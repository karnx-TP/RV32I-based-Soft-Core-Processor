module rv32i_core (clk,
    clkEn,
    dataBusInEn,
    rdEn,
    rstB,
    wrEn,
    RamMode,
    addr,
    dataBusIn,
    dataBusOut,
    inst_in,
    pc);
 input clk;
 input clkEn;
 input dataBusInEn;
 output rdEn;
 input rstB;
 output wrEn;
 output [3:0] RamMode;
 output [31:0] addr;
 input [31:0] dataBusIn;
 output [31:0] dataBusOut;
 input [31:0] inst_in;
 output [31:0] pc;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire \alu.b_type ;
 wire \alu.op_consShf ;
 wire \alu.r_type ;
 wire \brancher.funct3[0] ;
 wire \brancher.funct3[1] ;
 wire \brancher.funct3[2] ;
 wire \brancher.imm12_i_s[0] ;
 wire \brancher.imm12_i_s[10] ;
 wire \brancher.imm12_i_s[11] ;
 wire \brancher.imm12_i_s[1] ;
 wire \brancher.imm12_i_s[2] ;
 wire \brancher.imm12_i_s[3] ;
 wire \brancher.imm12_i_s[4] ;
 wire \brancher.imm12_i_s[5] ;
 wire \brancher.imm12_i_s[6] ;
 wire \brancher.imm12_i_s[7] ;
 wire \brancher.imm12_i_s[8] ;
 wire \brancher.imm12_i_s[9] ;
 wire \brancher.imm13_b[10] ;
 wire \brancher.imm13_b[11] ;
 wire \brancher.imm13_b[12] ;
 wire \brancher.imm13_b[1] ;
 wire \brancher.imm13_b[2] ;
 wire \brancher.imm13_b[3] ;
 wire \brancher.imm13_b[4] ;
 wire \brancher.imm13_b[5] ;
 wire \brancher.imm13_b[6] ;
 wire \brancher.imm13_b[7] ;
 wire \brancher.imm13_b[8] ;
 wire \brancher.imm13_b[9] ;
 wire \brancher.imm21_j[11] ;
 wire \brancher.imm21_j[15] ;
 wire \brancher.imm21_j[16] ;
 wire \brancher.imm21_j[17] ;
 wire \brancher.imm21_j[18] ;
 wire \brancher.imm21_j[19] ;
 wire \brancher.imm21_j[1] ;
 wire \brancher.imm21_j[2] ;
 wire \brancher.imm21_j[3] ;
 wire \brancher.imm21_j[4] ;
 wire \brancher.op_jal ;
 wire \brancher.op_jalr ;
 wire \brancher.pc_return[0] ;
 wire \brancher.pc_return[10] ;
 wire \brancher.pc_return[11] ;
 wire \brancher.pc_return[12] ;
 wire \brancher.pc_return[13] ;
 wire \brancher.pc_return[14] ;
 wire \brancher.pc_return[15] ;
 wire \brancher.pc_return[16] ;
 wire \brancher.pc_return[17] ;
 wire \brancher.pc_return[18] ;
 wire \brancher.pc_return[19] ;
 wire \brancher.pc_return[1] ;
 wire \brancher.pc_return[20] ;
 wire \brancher.pc_return[21] ;
 wire \brancher.pc_return[22] ;
 wire \brancher.pc_return[23] ;
 wire \brancher.pc_return[24] ;
 wire \brancher.pc_return[25] ;
 wire \brancher.pc_return[26] ;
 wire \brancher.pc_return[27] ;
 wire \brancher.pc_return[28] ;
 wire \brancher.pc_return[29] ;
 wire \brancher.pc_return[2] ;
 wire \brancher.pc_return[30] ;
 wire \brancher.pc_return[31] ;
 wire \brancher.pc_return[3] ;
 wire \brancher.pc_return[4] ;
 wire \brancher.pc_return[5] ;
 wire \brancher.pc_return[6] ;
 wire \brancher.pc_return[7] ;
 wire \brancher.pc_return[8] ;
 wire \brancher.pc_return[9] ;
 wire \brancher.rJumping ;
 wire \brancher.rPc_current_reg2[0] ;
 wire \brancher.rPc_current_reg2[10] ;
 wire \brancher.rPc_current_reg2[11] ;
 wire \brancher.rPc_current_reg2[12] ;
 wire \brancher.rPc_current_reg2[13] ;
 wire \brancher.rPc_current_reg2[14] ;
 wire \brancher.rPc_current_reg2[15] ;
 wire \brancher.rPc_current_reg2[16] ;
 wire \brancher.rPc_current_reg2[17] ;
 wire \brancher.rPc_current_reg2[18] ;
 wire \brancher.rPc_current_reg2[19] ;
 wire \brancher.rPc_current_reg2[1] ;
 wire \brancher.rPc_current_reg2[20] ;
 wire \brancher.rPc_current_reg2[21] ;
 wire \brancher.rPc_current_reg2[22] ;
 wire \brancher.rPc_current_reg2[23] ;
 wire \brancher.rPc_current_reg2[24] ;
 wire \brancher.rPc_current_reg2[25] ;
 wire \brancher.rPc_current_reg2[26] ;
 wire \brancher.rPc_current_reg2[27] ;
 wire \brancher.rPc_current_reg2[28] ;
 wire \brancher.rPc_current_reg2[29] ;
 wire \brancher.rPc_current_reg2[2] ;
 wire \brancher.rPc_current_reg2[30] ;
 wire \brancher.rPc_current_reg2[31] ;
 wire \brancher.rPc_current_reg2[3] ;
 wire \brancher.rPc_current_reg2[4] ;
 wire \brancher.rPc_current_reg2[5] ;
 wire \brancher.rPc_current_reg2[6] ;
 wire \brancher.rPc_current_reg2[7] ;
 wire \brancher.rPc_current_reg2[8] ;
 wire \brancher.rPc_current_reg2[9] ;
 wire \brancher.stall ;
 wire \dec.op_auipc ;
 wire \dec.op_intRegImm ;
 wire \dec.op_lui ;
 wire \dec.op_memLd ;
 wire \dec.op_memSt ;
 wire \dec.rInstrustion[0] ;
 wire \dec.rInstrustion[10] ;
 wire \dec.rInstrustion[11] ;
 wire \dec.rInstrustion[12] ;
 wire \dec.rInstrustion[13] ;
 wire \dec.rInstrustion[14] ;
 wire \dec.rInstrustion[15] ;
 wire \dec.rInstrustion[16] ;
 wire \dec.rInstrustion[17] ;
 wire \dec.rInstrustion[18] ;
 wire \dec.rInstrustion[19] ;
 wire \dec.rInstrustion[1] ;
 wire \dec.rInstrustion[20] ;
 wire \dec.rInstrustion[21] ;
 wire \dec.rInstrustion[22] ;
 wire \dec.rInstrustion[23] ;
 wire \dec.rInstrustion[24] ;
 wire \dec.rInstrustion[25] ;
 wire \dec.rInstrustion[26] ;
 wire \dec.rInstrustion[27] ;
 wire \dec.rInstrustion[28] ;
 wire \dec.rInstrustion[29] ;
 wire \dec.rInstrustion[2] ;
 wire \dec.rInstrustion[30] ;
 wire \dec.rInstrustion[31] ;
 wire \dec.rInstrustion[3] ;
 wire \dec.rInstrustion[4] ;
 wire \dec.rInstrustion[5] ;
 wire \dec.rInstrustion[6] ;
 wire \dec.rInstrustion[7] ;
 wire \dec.rInstrustion[8] ;
 wire \dec.rInstrustion[9] ;
 wire \dec.rStall ;
 wire rHazardStallRs1;
 wire rHazardStallRs2;
 wire rOp_memLd;
 wire rOp_memLd2;
 wire rRegWrEn;
 wire rRegWrEn2;
 wire \rReg_d2[0] ;
 wire \rReg_d2[1] ;
 wire \rReg_d2[2] ;
 wire \rReg_d2[3] ;
 wire \rReg_d2[4] ;
 wire \rReg_d[0] ;
 wire \rReg_d[1] ;
 wire \rReg_d[2] ;
 wire \rReg_d[3] ;
 wire \rReg_d[4] ;
 wire \rWrDataWB[0] ;
 wire \rWrDataWB[10] ;
 wire \rWrDataWB[11] ;
 wire \rWrDataWB[12] ;
 wire \rWrDataWB[13] ;
 wire \rWrDataWB[14] ;
 wire \rWrDataWB[15] ;
 wire \rWrDataWB[16] ;
 wire \rWrDataWB[17] ;
 wire \rWrDataWB[18] ;
 wire \rWrDataWB[19] ;
 wire \rWrDataWB[1] ;
 wire \rWrDataWB[20] ;
 wire \rWrDataWB[21] ;
 wire \rWrDataWB[22] ;
 wire \rWrDataWB[23] ;
 wire \rWrDataWB[24] ;
 wire \rWrDataWB[25] ;
 wire \rWrDataWB[26] ;
 wire \rWrDataWB[27] ;
 wire \rWrDataWB[28] ;
 wire \rWrDataWB[29] ;
 wire \rWrDataWB[2] ;
 wire \rWrDataWB[30] ;
 wire \rWrDataWB[31] ;
 wire \rWrDataWB[3] ;
 wire \rWrDataWB[4] ;
 wire \rWrDataWB[5] ;
 wire \rWrDataWB[6] ;
 wire \rWrDataWB[7] ;
 wire \rWrDataWB[8] ;
 wire \rWrDataWB[9] ;
 wire \rWrData[0] ;
 wire \rWrData[10] ;
 wire \rWrData[11] ;
 wire \rWrData[12] ;
 wire \rWrData[13] ;
 wire \rWrData[14] ;
 wire \rWrData[15] ;
 wire \rWrData[16] ;
 wire \rWrData[17] ;
 wire \rWrData[18] ;
 wire \rWrData[19] ;
 wire \rWrData[1] ;
 wire \rWrData[20] ;
 wire \rWrData[21] ;
 wire \rWrData[22] ;
 wire \rWrData[23] ;
 wire \rWrData[24] ;
 wire \rWrData[25] ;
 wire \rWrData[26] ;
 wire \rWrData[27] ;
 wire \rWrData[28] ;
 wire \rWrData[29] ;
 wire \rWrData[2] ;
 wire \rWrData[30] ;
 wire \rWrData[31] ;
 wire \rWrData[3] ;
 wire \rWrData[4] ;
 wire \rWrData[5] ;
 wire \rWrData[6] ;
 wire \rWrData[7] ;
 wire \rWrData[8] ;
 wire \rWrData[9] ;
 wire \reg_module.gprf[0] ;
 wire \reg_module.gprf[1000] ;
 wire \reg_module.gprf[1001] ;
 wire \reg_module.gprf[1002] ;
 wire \reg_module.gprf[1003] ;
 wire \reg_module.gprf[1004] ;
 wire \reg_module.gprf[1005] ;
 wire \reg_module.gprf[1006] ;
 wire \reg_module.gprf[1007] ;
 wire \reg_module.gprf[1008] ;
 wire \reg_module.gprf[1009] ;
 wire \reg_module.gprf[100] ;
 wire \reg_module.gprf[1010] ;
 wire \reg_module.gprf[1011] ;
 wire \reg_module.gprf[1012] ;
 wire \reg_module.gprf[1013] ;
 wire \reg_module.gprf[1014] ;
 wire \reg_module.gprf[1015] ;
 wire \reg_module.gprf[1016] ;
 wire \reg_module.gprf[1017] ;
 wire \reg_module.gprf[1018] ;
 wire \reg_module.gprf[1019] ;
 wire \reg_module.gprf[101] ;
 wire \reg_module.gprf[1020] ;
 wire \reg_module.gprf[1021] ;
 wire \reg_module.gprf[1022] ;
 wire \reg_module.gprf[1023] ;
 wire \reg_module.gprf[102] ;
 wire \reg_module.gprf[103] ;
 wire \reg_module.gprf[104] ;
 wire \reg_module.gprf[105] ;
 wire \reg_module.gprf[106] ;
 wire \reg_module.gprf[107] ;
 wire \reg_module.gprf[108] ;
 wire \reg_module.gprf[109] ;
 wire \reg_module.gprf[10] ;
 wire \reg_module.gprf[110] ;
 wire \reg_module.gprf[111] ;
 wire \reg_module.gprf[112] ;
 wire \reg_module.gprf[113] ;
 wire \reg_module.gprf[114] ;
 wire \reg_module.gprf[115] ;
 wire \reg_module.gprf[116] ;
 wire \reg_module.gprf[117] ;
 wire \reg_module.gprf[118] ;
 wire \reg_module.gprf[119] ;
 wire \reg_module.gprf[11] ;
 wire \reg_module.gprf[120] ;
 wire \reg_module.gprf[121] ;
 wire \reg_module.gprf[122] ;
 wire \reg_module.gprf[123] ;
 wire \reg_module.gprf[124] ;
 wire \reg_module.gprf[125] ;
 wire \reg_module.gprf[126] ;
 wire \reg_module.gprf[127] ;
 wire \reg_module.gprf[128] ;
 wire \reg_module.gprf[129] ;
 wire \reg_module.gprf[12] ;
 wire \reg_module.gprf[130] ;
 wire \reg_module.gprf[131] ;
 wire \reg_module.gprf[132] ;
 wire \reg_module.gprf[133] ;
 wire \reg_module.gprf[134] ;
 wire \reg_module.gprf[135] ;
 wire \reg_module.gprf[136] ;
 wire \reg_module.gprf[137] ;
 wire \reg_module.gprf[138] ;
 wire \reg_module.gprf[139] ;
 wire \reg_module.gprf[13] ;
 wire \reg_module.gprf[140] ;
 wire \reg_module.gprf[141] ;
 wire \reg_module.gprf[142] ;
 wire \reg_module.gprf[143] ;
 wire \reg_module.gprf[144] ;
 wire \reg_module.gprf[145] ;
 wire \reg_module.gprf[146] ;
 wire \reg_module.gprf[147] ;
 wire \reg_module.gprf[148] ;
 wire \reg_module.gprf[149] ;
 wire \reg_module.gprf[14] ;
 wire \reg_module.gprf[150] ;
 wire \reg_module.gprf[151] ;
 wire \reg_module.gprf[152] ;
 wire \reg_module.gprf[153] ;
 wire \reg_module.gprf[154] ;
 wire \reg_module.gprf[155] ;
 wire \reg_module.gprf[156] ;
 wire \reg_module.gprf[157] ;
 wire \reg_module.gprf[158] ;
 wire \reg_module.gprf[159] ;
 wire \reg_module.gprf[15] ;
 wire \reg_module.gprf[160] ;
 wire \reg_module.gprf[161] ;
 wire \reg_module.gprf[162] ;
 wire \reg_module.gprf[163] ;
 wire \reg_module.gprf[164] ;
 wire \reg_module.gprf[165] ;
 wire \reg_module.gprf[166] ;
 wire \reg_module.gprf[167] ;
 wire \reg_module.gprf[168] ;
 wire \reg_module.gprf[169] ;
 wire \reg_module.gprf[16] ;
 wire \reg_module.gprf[170] ;
 wire \reg_module.gprf[171] ;
 wire \reg_module.gprf[172] ;
 wire \reg_module.gprf[173] ;
 wire \reg_module.gprf[174] ;
 wire \reg_module.gprf[175] ;
 wire \reg_module.gprf[176] ;
 wire \reg_module.gprf[177] ;
 wire \reg_module.gprf[178] ;
 wire \reg_module.gprf[179] ;
 wire \reg_module.gprf[17] ;
 wire \reg_module.gprf[180] ;
 wire \reg_module.gprf[181] ;
 wire \reg_module.gprf[182] ;
 wire \reg_module.gprf[183] ;
 wire \reg_module.gprf[184] ;
 wire \reg_module.gprf[185] ;
 wire \reg_module.gprf[186] ;
 wire \reg_module.gprf[187] ;
 wire \reg_module.gprf[188] ;
 wire \reg_module.gprf[189] ;
 wire \reg_module.gprf[18] ;
 wire \reg_module.gprf[190] ;
 wire \reg_module.gprf[191] ;
 wire \reg_module.gprf[192] ;
 wire \reg_module.gprf[193] ;
 wire \reg_module.gprf[194] ;
 wire \reg_module.gprf[195] ;
 wire \reg_module.gprf[196] ;
 wire \reg_module.gprf[197] ;
 wire \reg_module.gprf[198] ;
 wire \reg_module.gprf[199] ;
 wire \reg_module.gprf[19] ;
 wire \reg_module.gprf[1] ;
 wire \reg_module.gprf[200] ;
 wire \reg_module.gprf[201] ;
 wire \reg_module.gprf[202] ;
 wire \reg_module.gprf[203] ;
 wire \reg_module.gprf[204] ;
 wire \reg_module.gprf[205] ;
 wire \reg_module.gprf[206] ;
 wire \reg_module.gprf[207] ;
 wire \reg_module.gprf[208] ;
 wire \reg_module.gprf[209] ;
 wire \reg_module.gprf[20] ;
 wire \reg_module.gprf[210] ;
 wire \reg_module.gprf[211] ;
 wire \reg_module.gprf[212] ;
 wire \reg_module.gprf[213] ;
 wire \reg_module.gprf[214] ;
 wire \reg_module.gprf[215] ;
 wire \reg_module.gprf[216] ;
 wire \reg_module.gprf[217] ;
 wire \reg_module.gprf[218] ;
 wire \reg_module.gprf[219] ;
 wire \reg_module.gprf[21] ;
 wire \reg_module.gprf[220] ;
 wire \reg_module.gprf[221] ;
 wire \reg_module.gprf[222] ;
 wire \reg_module.gprf[223] ;
 wire \reg_module.gprf[224] ;
 wire \reg_module.gprf[225] ;
 wire \reg_module.gprf[226] ;
 wire \reg_module.gprf[227] ;
 wire \reg_module.gprf[228] ;
 wire \reg_module.gprf[229] ;
 wire \reg_module.gprf[22] ;
 wire \reg_module.gprf[230] ;
 wire \reg_module.gprf[231] ;
 wire \reg_module.gprf[232] ;
 wire \reg_module.gprf[233] ;
 wire \reg_module.gprf[234] ;
 wire \reg_module.gprf[235] ;
 wire \reg_module.gprf[236] ;
 wire \reg_module.gprf[237] ;
 wire \reg_module.gprf[238] ;
 wire \reg_module.gprf[239] ;
 wire \reg_module.gprf[23] ;
 wire \reg_module.gprf[240] ;
 wire \reg_module.gprf[241] ;
 wire \reg_module.gprf[242] ;
 wire \reg_module.gprf[243] ;
 wire \reg_module.gprf[244] ;
 wire \reg_module.gprf[245] ;
 wire \reg_module.gprf[246] ;
 wire \reg_module.gprf[247] ;
 wire \reg_module.gprf[248] ;
 wire \reg_module.gprf[249] ;
 wire \reg_module.gprf[24] ;
 wire \reg_module.gprf[250] ;
 wire \reg_module.gprf[251] ;
 wire \reg_module.gprf[252] ;
 wire \reg_module.gprf[253] ;
 wire \reg_module.gprf[254] ;
 wire \reg_module.gprf[255] ;
 wire \reg_module.gprf[256] ;
 wire \reg_module.gprf[257] ;
 wire \reg_module.gprf[258] ;
 wire \reg_module.gprf[259] ;
 wire \reg_module.gprf[25] ;
 wire \reg_module.gprf[260] ;
 wire \reg_module.gprf[261] ;
 wire \reg_module.gprf[262] ;
 wire \reg_module.gprf[263] ;
 wire \reg_module.gprf[264] ;
 wire \reg_module.gprf[265] ;
 wire \reg_module.gprf[266] ;
 wire \reg_module.gprf[267] ;
 wire \reg_module.gprf[268] ;
 wire \reg_module.gprf[269] ;
 wire \reg_module.gprf[26] ;
 wire \reg_module.gprf[270] ;
 wire \reg_module.gprf[271] ;
 wire \reg_module.gprf[272] ;
 wire \reg_module.gprf[273] ;
 wire \reg_module.gprf[274] ;
 wire \reg_module.gprf[275] ;
 wire \reg_module.gprf[276] ;
 wire \reg_module.gprf[277] ;
 wire \reg_module.gprf[278] ;
 wire \reg_module.gprf[279] ;
 wire \reg_module.gprf[27] ;
 wire \reg_module.gprf[280] ;
 wire \reg_module.gprf[281] ;
 wire \reg_module.gprf[282] ;
 wire \reg_module.gprf[283] ;
 wire \reg_module.gprf[284] ;
 wire \reg_module.gprf[285] ;
 wire \reg_module.gprf[286] ;
 wire \reg_module.gprf[287] ;
 wire \reg_module.gprf[288] ;
 wire \reg_module.gprf[289] ;
 wire \reg_module.gprf[28] ;
 wire \reg_module.gprf[290] ;
 wire \reg_module.gprf[291] ;
 wire \reg_module.gprf[292] ;
 wire \reg_module.gprf[293] ;
 wire \reg_module.gprf[294] ;
 wire \reg_module.gprf[295] ;
 wire \reg_module.gprf[296] ;
 wire \reg_module.gprf[297] ;
 wire \reg_module.gprf[298] ;
 wire \reg_module.gprf[299] ;
 wire \reg_module.gprf[29] ;
 wire \reg_module.gprf[2] ;
 wire \reg_module.gprf[300] ;
 wire \reg_module.gprf[301] ;
 wire \reg_module.gprf[302] ;
 wire \reg_module.gprf[303] ;
 wire \reg_module.gprf[304] ;
 wire \reg_module.gprf[305] ;
 wire \reg_module.gprf[306] ;
 wire \reg_module.gprf[307] ;
 wire \reg_module.gprf[308] ;
 wire \reg_module.gprf[309] ;
 wire \reg_module.gprf[30] ;
 wire \reg_module.gprf[310] ;
 wire \reg_module.gprf[311] ;
 wire \reg_module.gprf[312] ;
 wire \reg_module.gprf[313] ;
 wire \reg_module.gprf[314] ;
 wire \reg_module.gprf[315] ;
 wire \reg_module.gprf[316] ;
 wire \reg_module.gprf[317] ;
 wire \reg_module.gprf[318] ;
 wire \reg_module.gprf[319] ;
 wire \reg_module.gprf[31] ;
 wire \reg_module.gprf[320] ;
 wire \reg_module.gprf[321] ;
 wire \reg_module.gprf[322] ;
 wire \reg_module.gprf[323] ;
 wire \reg_module.gprf[324] ;
 wire \reg_module.gprf[325] ;
 wire \reg_module.gprf[326] ;
 wire \reg_module.gprf[327] ;
 wire \reg_module.gprf[328] ;
 wire \reg_module.gprf[329] ;
 wire \reg_module.gprf[32] ;
 wire \reg_module.gprf[330] ;
 wire \reg_module.gprf[331] ;
 wire \reg_module.gprf[332] ;
 wire \reg_module.gprf[333] ;
 wire \reg_module.gprf[334] ;
 wire \reg_module.gprf[335] ;
 wire \reg_module.gprf[336] ;
 wire \reg_module.gprf[337] ;
 wire \reg_module.gprf[338] ;
 wire \reg_module.gprf[339] ;
 wire \reg_module.gprf[33] ;
 wire \reg_module.gprf[340] ;
 wire \reg_module.gprf[341] ;
 wire \reg_module.gprf[342] ;
 wire \reg_module.gprf[343] ;
 wire \reg_module.gprf[344] ;
 wire \reg_module.gprf[345] ;
 wire \reg_module.gprf[346] ;
 wire \reg_module.gprf[347] ;
 wire \reg_module.gprf[348] ;
 wire \reg_module.gprf[349] ;
 wire \reg_module.gprf[34] ;
 wire \reg_module.gprf[350] ;
 wire \reg_module.gprf[351] ;
 wire \reg_module.gprf[352] ;
 wire \reg_module.gprf[353] ;
 wire \reg_module.gprf[354] ;
 wire \reg_module.gprf[355] ;
 wire \reg_module.gprf[356] ;
 wire \reg_module.gprf[357] ;
 wire \reg_module.gprf[358] ;
 wire \reg_module.gprf[359] ;
 wire \reg_module.gprf[35] ;
 wire \reg_module.gprf[360] ;
 wire \reg_module.gprf[361] ;
 wire \reg_module.gprf[362] ;
 wire \reg_module.gprf[363] ;
 wire \reg_module.gprf[364] ;
 wire \reg_module.gprf[365] ;
 wire \reg_module.gprf[366] ;
 wire \reg_module.gprf[367] ;
 wire \reg_module.gprf[368] ;
 wire \reg_module.gprf[369] ;
 wire \reg_module.gprf[36] ;
 wire \reg_module.gprf[370] ;
 wire \reg_module.gprf[371] ;
 wire \reg_module.gprf[372] ;
 wire \reg_module.gprf[373] ;
 wire \reg_module.gprf[374] ;
 wire \reg_module.gprf[375] ;
 wire \reg_module.gprf[376] ;
 wire \reg_module.gprf[377] ;
 wire \reg_module.gprf[378] ;
 wire \reg_module.gprf[379] ;
 wire \reg_module.gprf[37] ;
 wire \reg_module.gprf[380] ;
 wire \reg_module.gprf[381] ;
 wire \reg_module.gprf[382] ;
 wire \reg_module.gprf[383] ;
 wire \reg_module.gprf[384] ;
 wire \reg_module.gprf[385] ;
 wire \reg_module.gprf[386] ;
 wire \reg_module.gprf[387] ;
 wire \reg_module.gprf[388] ;
 wire \reg_module.gprf[389] ;
 wire \reg_module.gprf[38] ;
 wire \reg_module.gprf[390] ;
 wire \reg_module.gprf[391] ;
 wire \reg_module.gprf[392] ;
 wire \reg_module.gprf[393] ;
 wire \reg_module.gprf[394] ;
 wire \reg_module.gprf[395] ;
 wire \reg_module.gprf[396] ;
 wire \reg_module.gprf[397] ;
 wire \reg_module.gprf[398] ;
 wire \reg_module.gprf[399] ;
 wire \reg_module.gprf[39] ;
 wire \reg_module.gprf[3] ;
 wire \reg_module.gprf[400] ;
 wire \reg_module.gprf[401] ;
 wire \reg_module.gprf[402] ;
 wire \reg_module.gprf[403] ;
 wire \reg_module.gprf[404] ;
 wire \reg_module.gprf[405] ;
 wire \reg_module.gprf[406] ;
 wire \reg_module.gprf[407] ;
 wire \reg_module.gprf[408] ;
 wire \reg_module.gprf[409] ;
 wire \reg_module.gprf[40] ;
 wire \reg_module.gprf[410] ;
 wire \reg_module.gprf[411] ;
 wire \reg_module.gprf[412] ;
 wire \reg_module.gprf[413] ;
 wire \reg_module.gprf[414] ;
 wire \reg_module.gprf[415] ;
 wire \reg_module.gprf[416] ;
 wire \reg_module.gprf[417] ;
 wire \reg_module.gprf[418] ;
 wire \reg_module.gprf[419] ;
 wire \reg_module.gprf[41] ;
 wire \reg_module.gprf[420] ;
 wire \reg_module.gprf[421] ;
 wire \reg_module.gprf[422] ;
 wire \reg_module.gprf[423] ;
 wire \reg_module.gprf[424] ;
 wire \reg_module.gprf[425] ;
 wire \reg_module.gprf[426] ;
 wire \reg_module.gprf[427] ;
 wire \reg_module.gprf[428] ;
 wire \reg_module.gprf[429] ;
 wire \reg_module.gprf[42] ;
 wire \reg_module.gprf[430] ;
 wire \reg_module.gprf[431] ;
 wire \reg_module.gprf[432] ;
 wire \reg_module.gprf[433] ;
 wire \reg_module.gprf[434] ;
 wire \reg_module.gprf[435] ;
 wire \reg_module.gprf[436] ;
 wire \reg_module.gprf[437] ;
 wire \reg_module.gprf[438] ;
 wire \reg_module.gprf[439] ;
 wire \reg_module.gprf[43] ;
 wire \reg_module.gprf[440] ;
 wire \reg_module.gprf[441] ;
 wire \reg_module.gprf[442] ;
 wire \reg_module.gprf[443] ;
 wire \reg_module.gprf[444] ;
 wire \reg_module.gprf[445] ;
 wire \reg_module.gprf[446] ;
 wire \reg_module.gprf[447] ;
 wire \reg_module.gprf[448] ;
 wire \reg_module.gprf[449] ;
 wire \reg_module.gprf[44] ;
 wire \reg_module.gprf[450] ;
 wire \reg_module.gprf[451] ;
 wire \reg_module.gprf[452] ;
 wire \reg_module.gprf[453] ;
 wire \reg_module.gprf[454] ;
 wire \reg_module.gprf[455] ;
 wire \reg_module.gprf[456] ;
 wire \reg_module.gprf[457] ;
 wire \reg_module.gprf[458] ;
 wire \reg_module.gprf[459] ;
 wire \reg_module.gprf[45] ;
 wire \reg_module.gprf[460] ;
 wire \reg_module.gprf[461] ;
 wire \reg_module.gprf[462] ;
 wire \reg_module.gprf[463] ;
 wire \reg_module.gprf[464] ;
 wire \reg_module.gprf[465] ;
 wire \reg_module.gprf[466] ;
 wire \reg_module.gprf[467] ;
 wire \reg_module.gprf[468] ;
 wire \reg_module.gprf[469] ;
 wire \reg_module.gprf[46] ;
 wire \reg_module.gprf[470] ;
 wire \reg_module.gprf[471] ;
 wire \reg_module.gprf[472] ;
 wire \reg_module.gprf[473] ;
 wire \reg_module.gprf[474] ;
 wire \reg_module.gprf[475] ;
 wire \reg_module.gprf[476] ;
 wire \reg_module.gprf[477] ;
 wire \reg_module.gprf[478] ;
 wire \reg_module.gprf[479] ;
 wire \reg_module.gprf[47] ;
 wire \reg_module.gprf[480] ;
 wire \reg_module.gprf[481] ;
 wire \reg_module.gprf[482] ;
 wire \reg_module.gprf[483] ;
 wire \reg_module.gprf[484] ;
 wire \reg_module.gprf[485] ;
 wire \reg_module.gprf[486] ;
 wire \reg_module.gprf[487] ;
 wire \reg_module.gprf[488] ;
 wire \reg_module.gprf[489] ;
 wire \reg_module.gprf[48] ;
 wire \reg_module.gprf[490] ;
 wire \reg_module.gprf[491] ;
 wire \reg_module.gprf[492] ;
 wire \reg_module.gprf[493] ;
 wire \reg_module.gprf[494] ;
 wire \reg_module.gprf[495] ;
 wire \reg_module.gprf[496] ;
 wire \reg_module.gprf[497] ;
 wire \reg_module.gprf[498] ;
 wire \reg_module.gprf[499] ;
 wire \reg_module.gprf[49] ;
 wire \reg_module.gprf[4] ;
 wire \reg_module.gprf[500] ;
 wire \reg_module.gprf[501] ;
 wire \reg_module.gprf[502] ;
 wire \reg_module.gprf[503] ;
 wire \reg_module.gprf[504] ;
 wire \reg_module.gprf[505] ;
 wire \reg_module.gprf[506] ;
 wire \reg_module.gprf[507] ;
 wire \reg_module.gprf[508] ;
 wire \reg_module.gprf[509] ;
 wire \reg_module.gprf[50] ;
 wire \reg_module.gprf[510] ;
 wire \reg_module.gprf[511] ;
 wire \reg_module.gprf[512] ;
 wire \reg_module.gprf[513] ;
 wire \reg_module.gprf[514] ;
 wire \reg_module.gprf[515] ;
 wire \reg_module.gprf[516] ;
 wire \reg_module.gprf[517] ;
 wire \reg_module.gprf[518] ;
 wire \reg_module.gprf[519] ;
 wire \reg_module.gprf[51] ;
 wire \reg_module.gprf[520] ;
 wire \reg_module.gprf[521] ;
 wire \reg_module.gprf[522] ;
 wire \reg_module.gprf[523] ;
 wire \reg_module.gprf[524] ;
 wire \reg_module.gprf[525] ;
 wire \reg_module.gprf[526] ;
 wire \reg_module.gprf[527] ;
 wire \reg_module.gprf[528] ;
 wire \reg_module.gprf[529] ;
 wire \reg_module.gprf[52] ;
 wire \reg_module.gprf[530] ;
 wire \reg_module.gprf[531] ;
 wire \reg_module.gprf[532] ;
 wire \reg_module.gprf[533] ;
 wire \reg_module.gprf[534] ;
 wire \reg_module.gprf[535] ;
 wire \reg_module.gprf[536] ;
 wire \reg_module.gprf[537] ;
 wire \reg_module.gprf[538] ;
 wire \reg_module.gprf[539] ;
 wire \reg_module.gprf[53] ;
 wire \reg_module.gprf[540] ;
 wire \reg_module.gprf[541] ;
 wire \reg_module.gprf[542] ;
 wire \reg_module.gprf[543] ;
 wire \reg_module.gprf[544] ;
 wire \reg_module.gprf[545] ;
 wire \reg_module.gprf[546] ;
 wire \reg_module.gprf[547] ;
 wire \reg_module.gprf[548] ;
 wire \reg_module.gprf[549] ;
 wire \reg_module.gprf[54] ;
 wire \reg_module.gprf[550] ;
 wire \reg_module.gprf[551] ;
 wire \reg_module.gprf[552] ;
 wire \reg_module.gprf[553] ;
 wire \reg_module.gprf[554] ;
 wire \reg_module.gprf[555] ;
 wire \reg_module.gprf[556] ;
 wire \reg_module.gprf[557] ;
 wire \reg_module.gprf[558] ;
 wire \reg_module.gprf[559] ;
 wire \reg_module.gprf[55] ;
 wire \reg_module.gprf[560] ;
 wire \reg_module.gprf[561] ;
 wire \reg_module.gprf[562] ;
 wire \reg_module.gprf[563] ;
 wire \reg_module.gprf[564] ;
 wire \reg_module.gprf[565] ;
 wire \reg_module.gprf[566] ;
 wire \reg_module.gprf[567] ;
 wire \reg_module.gprf[568] ;
 wire \reg_module.gprf[569] ;
 wire \reg_module.gprf[56] ;
 wire \reg_module.gprf[570] ;
 wire \reg_module.gprf[571] ;
 wire \reg_module.gprf[572] ;
 wire \reg_module.gprf[573] ;
 wire \reg_module.gprf[574] ;
 wire \reg_module.gprf[575] ;
 wire \reg_module.gprf[576] ;
 wire \reg_module.gprf[577] ;
 wire \reg_module.gprf[578] ;
 wire \reg_module.gprf[579] ;
 wire \reg_module.gprf[57] ;
 wire \reg_module.gprf[580] ;
 wire \reg_module.gprf[581] ;
 wire \reg_module.gprf[582] ;
 wire \reg_module.gprf[583] ;
 wire \reg_module.gprf[584] ;
 wire \reg_module.gprf[585] ;
 wire \reg_module.gprf[586] ;
 wire \reg_module.gprf[587] ;
 wire \reg_module.gprf[588] ;
 wire \reg_module.gprf[589] ;
 wire \reg_module.gprf[58] ;
 wire \reg_module.gprf[590] ;
 wire \reg_module.gprf[591] ;
 wire \reg_module.gprf[592] ;
 wire \reg_module.gprf[593] ;
 wire \reg_module.gprf[594] ;
 wire \reg_module.gprf[595] ;
 wire \reg_module.gprf[596] ;
 wire \reg_module.gprf[597] ;
 wire \reg_module.gprf[598] ;
 wire \reg_module.gprf[599] ;
 wire \reg_module.gprf[59] ;
 wire \reg_module.gprf[5] ;
 wire \reg_module.gprf[600] ;
 wire \reg_module.gprf[601] ;
 wire \reg_module.gprf[602] ;
 wire \reg_module.gprf[603] ;
 wire \reg_module.gprf[604] ;
 wire \reg_module.gprf[605] ;
 wire \reg_module.gprf[606] ;
 wire \reg_module.gprf[607] ;
 wire \reg_module.gprf[608] ;
 wire \reg_module.gprf[609] ;
 wire \reg_module.gprf[60] ;
 wire \reg_module.gprf[610] ;
 wire \reg_module.gprf[611] ;
 wire \reg_module.gprf[612] ;
 wire \reg_module.gprf[613] ;
 wire \reg_module.gprf[614] ;
 wire \reg_module.gprf[615] ;
 wire \reg_module.gprf[616] ;
 wire \reg_module.gprf[617] ;
 wire \reg_module.gprf[618] ;
 wire \reg_module.gprf[619] ;
 wire \reg_module.gprf[61] ;
 wire \reg_module.gprf[620] ;
 wire \reg_module.gprf[621] ;
 wire \reg_module.gprf[622] ;
 wire \reg_module.gprf[623] ;
 wire \reg_module.gprf[624] ;
 wire \reg_module.gprf[625] ;
 wire \reg_module.gprf[626] ;
 wire \reg_module.gprf[627] ;
 wire \reg_module.gprf[628] ;
 wire \reg_module.gprf[629] ;
 wire \reg_module.gprf[62] ;
 wire \reg_module.gprf[630] ;
 wire \reg_module.gprf[631] ;
 wire \reg_module.gprf[632] ;
 wire \reg_module.gprf[633] ;
 wire \reg_module.gprf[634] ;
 wire \reg_module.gprf[635] ;
 wire \reg_module.gprf[636] ;
 wire \reg_module.gprf[637] ;
 wire \reg_module.gprf[638] ;
 wire \reg_module.gprf[639] ;
 wire \reg_module.gprf[63] ;
 wire \reg_module.gprf[640] ;
 wire \reg_module.gprf[641] ;
 wire \reg_module.gprf[642] ;
 wire \reg_module.gprf[643] ;
 wire \reg_module.gprf[644] ;
 wire \reg_module.gprf[645] ;
 wire \reg_module.gprf[646] ;
 wire \reg_module.gprf[647] ;
 wire \reg_module.gprf[648] ;
 wire \reg_module.gprf[649] ;
 wire \reg_module.gprf[64] ;
 wire \reg_module.gprf[650] ;
 wire \reg_module.gprf[651] ;
 wire \reg_module.gprf[652] ;
 wire \reg_module.gprf[653] ;
 wire \reg_module.gprf[654] ;
 wire \reg_module.gprf[655] ;
 wire \reg_module.gprf[656] ;
 wire \reg_module.gprf[657] ;
 wire \reg_module.gprf[658] ;
 wire \reg_module.gprf[659] ;
 wire \reg_module.gprf[65] ;
 wire \reg_module.gprf[660] ;
 wire \reg_module.gprf[661] ;
 wire \reg_module.gprf[662] ;
 wire \reg_module.gprf[663] ;
 wire \reg_module.gprf[664] ;
 wire \reg_module.gprf[665] ;
 wire \reg_module.gprf[666] ;
 wire \reg_module.gprf[667] ;
 wire \reg_module.gprf[668] ;
 wire \reg_module.gprf[669] ;
 wire \reg_module.gprf[66] ;
 wire \reg_module.gprf[670] ;
 wire \reg_module.gprf[671] ;
 wire \reg_module.gprf[672] ;
 wire \reg_module.gprf[673] ;
 wire \reg_module.gprf[674] ;
 wire \reg_module.gprf[675] ;
 wire \reg_module.gprf[676] ;
 wire \reg_module.gprf[677] ;
 wire \reg_module.gprf[678] ;
 wire \reg_module.gprf[679] ;
 wire \reg_module.gprf[67] ;
 wire \reg_module.gprf[680] ;
 wire \reg_module.gprf[681] ;
 wire \reg_module.gprf[682] ;
 wire \reg_module.gprf[683] ;
 wire \reg_module.gprf[684] ;
 wire \reg_module.gprf[685] ;
 wire \reg_module.gprf[686] ;
 wire \reg_module.gprf[687] ;
 wire \reg_module.gprf[688] ;
 wire \reg_module.gprf[689] ;
 wire \reg_module.gprf[68] ;
 wire \reg_module.gprf[690] ;
 wire \reg_module.gprf[691] ;
 wire \reg_module.gprf[692] ;
 wire \reg_module.gprf[693] ;
 wire \reg_module.gprf[694] ;
 wire \reg_module.gprf[695] ;
 wire \reg_module.gprf[696] ;
 wire \reg_module.gprf[697] ;
 wire \reg_module.gprf[698] ;
 wire \reg_module.gprf[699] ;
 wire \reg_module.gprf[69] ;
 wire \reg_module.gprf[6] ;
 wire \reg_module.gprf[700] ;
 wire \reg_module.gprf[701] ;
 wire \reg_module.gprf[702] ;
 wire \reg_module.gprf[703] ;
 wire \reg_module.gprf[704] ;
 wire \reg_module.gprf[705] ;
 wire \reg_module.gprf[706] ;
 wire \reg_module.gprf[707] ;
 wire \reg_module.gprf[708] ;
 wire \reg_module.gprf[709] ;
 wire \reg_module.gprf[70] ;
 wire \reg_module.gprf[710] ;
 wire \reg_module.gprf[711] ;
 wire \reg_module.gprf[712] ;
 wire \reg_module.gprf[713] ;
 wire \reg_module.gprf[714] ;
 wire \reg_module.gprf[715] ;
 wire \reg_module.gprf[716] ;
 wire \reg_module.gprf[717] ;
 wire \reg_module.gprf[718] ;
 wire \reg_module.gprf[719] ;
 wire \reg_module.gprf[71] ;
 wire \reg_module.gprf[720] ;
 wire \reg_module.gprf[721] ;
 wire \reg_module.gprf[722] ;
 wire \reg_module.gprf[723] ;
 wire \reg_module.gprf[724] ;
 wire \reg_module.gprf[725] ;
 wire \reg_module.gprf[726] ;
 wire \reg_module.gprf[727] ;
 wire \reg_module.gprf[728] ;
 wire \reg_module.gprf[729] ;
 wire \reg_module.gprf[72] ;
 wire \reg_module.gprf[730] ;
 wire \reg_module.gprf[731] ;
 wire \reg_module.gprf[732] ;
 wire \reg_module.gprf[733] ;
 wire \reg_module.gprf[734] ;
 wire \reg_module.gprf[735] ;
 wire \reg_module.gprf[736] ;
 wire \reg_module.gprf[737] ;
 wire \reg_module.gprf[738] ;
 wire \reg_module.gprf[739] ;
 wire \reg_module.gprf[73] ;
 wire \reg_module.gprf[740] ;
 wire \reg_module.gprf[741] ;
 wire \reg_module.gprf[742] ;
 wire \reg_module.gprf[743] ;
 wire \reg_module.gprf[744] ;
 wire \reg_module.gprf[745] ;
 wire \reg_module.gprf[746] ;
 wire \reg_module.gprf[747] ;
 wire \reg_module.gprf[748] ;
 wire \reg_module.gprf[749] ;
 wire \reg_module.gprf[74] ;
 wire \reg_module.gprf[750] ;
 wire \reg_module.gprf[751] ;
 wire \reg_module.gprf[752] ;
 wire \reg_module.gprf[753] ;
 wire \reg_module.gprf[754] ;
 wire \reg_module.gprf[755] ;
 wire \reg_module.gprf[756] ;
 wire \reg_module.gprf[757] ;
 wire \reg_module.gprf[758] ;
 wire \reg_module.gprf[759] ;
 wire \reg_module.gprf[75] ;
 wire \reg_module.gprf[760] ;
 wire \reg_module.gprf[761] ;
 wire \reg_module.gprf[762] ;
 wire \reg_module.gprf[763] ;
 wire \reg_module.gprf[764] ;
 wire \reg_module.gprf[765] ;
 wire \reg_module.gprf[766] ;
 wire \reg_module.gprf[767] ;
 wire \reg_module.gprf[768] ;
 wire \reg_module.gprf[769] ;
 wire \reg_module.gprf[76] ;
 wire \reg_module.gprf[770] ;
 wire \reg_module.gprf[771] ;
 wire \reg_module.gprf[772] ;
 wire \reg_module.gprf[773] ;
 wire \reg_module.gprf[774] ;
 wire \reg_module.gprf[775] ;
 wire \reg_module.gprf[776] ;
 wire \reg_module.gprf[777] ;
 wire \reg_module.gprf[778] ;
 wire \reg_module.gprf[779] ;
 wire \reg_module.gprf[77] ;
 wire \reg_module.gprf[780] ;
 wire \reg_module.gprf[781] ;
 wire \reg_module.gprf[782] ;
 wire \reg_module.gprf[783] ;
 wire \reg_module.gprf[784] ;
 wire \reg_module.gprf[785] ;
 wire \reg_module.gprf[786] ;
 wire \reg_module.gprf[787] ;
 wire \reg_module.gprf[788] ;
 wire \reg_module.gprf[789] ;
 wire \reg_module.gprf[78] ;
 wire \reg_module.gprf[790] ;
 wire \reg_module.gprf[791] ;
 wire \reg_module.gprf[792] ;
 wire \reg_module.gprf[793] ;
 wire \reg_module.gprf[794] ;
 wire \reg_module.gprf[795] ;
 wire \reg_module.gprf[796] ;
 wire \reg_module.gprf[797] ;
 wire \reg_module.gprf[798] ;
 wire \reg_module.gprf[799] ;
 wire \reg_module.gprf[79] ;
 wire \reg_module.gprf[7] ;
 wire \reg_module.gprf[800] ;
 wire \reg_module.gprf[801] ;
 wire \reg_module.gprf[802] ;
 wire \reg_module.gprf[803] ;
 wire \reg_module.gprf[804] ;
 wire \reg_module.gprf[805] ;
 wire \reg_module.gprf[806] ;
 wire \reg_module.gprf[807] ;
 wire \reg_module.gprf[808] ;
 wire \reg_module.gprf[809] ;
 wire \reg_module.gprf[80] ;
 wire \reg_module.gprf[810] ;
 wire \reg_module.gprf[811] ;
 wire \reg_module.gprf[812] ;
 wire \reg_module.gprf[813] ;
 wire \reg_module.gprf[814] ;
 wire \reg_module.gprf[815] ;
 wire \reg_module.gprf[816] ;
 wire \reg_module.gprf[817] ;
 wire \reg_module.gprf[818] ;
 wire \reg_module.gprf[819] ;
 wire \reg_module.gprf[81] ;
 wire \reg_module.gprf[820] ;
 wire \reg_module.gprf[821] ;
 wire \reg_module.gprf[822] ;
 wire \reg_module.gprf[823] ;
 wire \reg_module.gprf[824] ;
 wire \reg_module.gprf[825] ;
 wire \reg_module.gprf[826] ;
 wire \reg_module.gprf[827] ;
 wire \reg_module.gprf[828] ;
 wire \reg_module.gprf[829] ;
 wire \reg_module.gprf[82] ;
 wire \reg_module.gprf[830] ;
 wire \reg_module.gprf[831] ;
 wire \reg_module.gprf[832] ;
 wire \reg_module.gprf[833] ;
 wire \reg_module.gprf[834] ;
 wire \reg_module.gprf[835] ;
 wire \reg_module.gprf[836] ;
 wire \reg_module.gprf[837] ;
 wire \reg_module.gprf[838] ;
 wire \reg_module.gprf[839] ;
 wire \reg_module.gprf[83] ;
 wire \reg_module.gprf[840] ;
 wire \reg_module.gprf[841] ;
 wire \reg_module.gprf[842] ;
 wire \reg_module.gprf[843] ;
 wire \reg_module.gprf[844] ;
 wire \reg_module.gprf[845] ;
 wire \reg_module.gprf[846] ;
 wire \reg_module.gprf[847] ;
 wire \reg_module.gprf[848] ;
 wire \reg_module.gprf[849] ;
 wire \reg_module.gprf[84] ;
 wire \reg_module.gprf[850] ;
 wire \reg_module.gprf[851] ;
 wire \reg_module.gprf[852] ;
 wire \reg_module.gprf[853] ;
 wire \reg_module.gprf[854] ;
 wire \reg_module.gprf[855] ;
 wire \reg_module.gprf[856] ;
 wire \reg_module.gprf[857] ;
 wire \reg_module.gprf[858] ;
 wire \reg_module.gprf[859] ;
 wire \reg_module.gprf[85] ;
 wire \reg_module.gprf[860] ;
 wire \reg_module.gprf[861] ;
 wire \reg_module.gprf[862] ;
 wire \reg_module.gprf[863] ;
 wire \reg_module.gprf[864] ;
 wire \reg_module.gprf[865] ;
 wire \reg_module.gprf[866] ;
 wire \reg_module.gprf[867] ;
 wire \reg_module.gprf[868] ;
 wire \reg_module.gprf[869] ;
 wire \reg_module.gprf[86] ;
 wire \reg_module.gprf[870] ;
 wire \reg_module.gprf[871] ;
 wire \reg_module.gprf[872] ;
 wire \reg_module.gprf[873] ;
 wire \reg_module.gprf[874] ;
 wire \reg_module.gprf[875] ;
 wire \reg_module.gprf[876] ;
 wire \reg_module.gprf[877] ;
 wire \reg_module.gprf[878] ;
 wire \reg_module.gprf[879] ;
 wire \reg_module.gprf[87] ;
 wire \reg_module.gprf[880] ;
 wire \reg_module.gprf[881] ;
 wire \reg_module.gprf[882] ;
 wire \reg_module.gprf[883] ;
 wire \reg_module.gprf[884] ;
 wire \reg_module.gprf[885] ;
 wire \reg_module.gprf[886] ;
 wire \reg_module.gprf[887] ;
 wire \reg_module.gprf[888] ;
 wire \reg_module.gprf[889] ;
 wire \reg_module.gprf[88] ;
 wire \reg_module.gprf[890] ;
 wire \reg_module.gprf[891] ;
 wire \reg_module.gprf[892] ;
 wire \reg_module.gprf[893] ;
 wire \reg_module.gprf[894] ;
 wire \reg_module.gprf[895] ;
 wire \reg_module.gprf[896] ;
 wire \reg_module.gprf[897] ;
 wire \reg_module.gprf[898] ;
 wire \reg_module.gprf[899] ;
 wire \reg_module.gprf[89] ;
 wire \reg_module.gprf[8] ;
 wire \reg_module.gprf[900] ;
 wire \reg_module.gprf[901] ;
 wire \reg_module.gprf[902] ;
 wire \reg_module.gprf[903] ;
 wire \reg_module.gprf[904] ;
 wire \reg_module.gprf[905] ;
 wire \reg_module.gprf[906] ;
 wire \reg_module.gprf[907] ;
 wire \reg_module.gprf[908] ;
 wire \reg_module.gprf[909] ;
 wire \reg_module.gprf[90] ;
 wire \reg_module.gprf[910] ;
 wire \reg_module.gprf[911] ;
 wire \reg_module.gprf[912] ;
 wire \reg_module.gprf[913] ;
 wire \reg_module.gprf[914] ;
 wire \reg_module.gprf[915] ;
 wire \reg_module.gprf[916] ;
 wire \reg_module.gprf[917] ;
 wire \reg_module.gprf[918] ;
 wire \reg_module.gprf[919] ;
 wire \reg_module.gprf[91] ;
 wire \reg_module.gprf[920] ;
 wire \reg_module.gprf[921] ;
 wire \reg_module.gprf[922] ;
 wire \reg_module.gprf[923] ;
 wire \reg_module.gprf[924] ;
 wire \reg_module.gprf[925] ;
 wire \reg_module.gprf[926] ;
 wire \reg_module.gprf[927] ;
 wire \reg_module.gprf[928] ;
 wire \reg_module.gprf[929] ;
 wire \reg_module.gprf[92] ;
 wire \reg_module.gprf[930] ;
 wire \reg_module.gprf[931] ;
 wire \reg_module.gprf[932] ;
 wire \reg_module.gprf[933] ;
 wire \reg_module.gprf[934] ;
 wire \reg_module.gprf[935] ;
 wire \reg_module.gprf[936] ;
 wire \reg_module.gprf[937] ;
 wire \reg_module.gprf[938] ;
 wire \reg_module.gprf[939] ;
 wire \reg_module.gprf[93] ;
 wire \reg_module.gprf[940] ;
 wire \reg_module.gprf[941] ;
 wire \reg_module.gprf[942] ;
 wire \reg_module.gprf[943] ;
 wire \reg_module.gprf[944] ;
 wire \reg_module.gprf[945] ;
 wire \reg_module.gprf[946] ;
 wire \reg_module.gprf[947] ;
 wire \reg_module.gprf[948] ;
 wire \reg_module.gprf[949] ;
 wire \reg_module.gprf[94] ;
 wire \reg_module.gprf[950] ;
 wire \reg_module.gprf[951] ;
 wire \reg_module.gprf[952] ;
 wire \reg_module.gprf[953] ;
 wire \reg_module.gprf[954] ;
 wire \reg_module.gprf[955] ;
 wire \reg_module.gprf[956] ;
 wire \reg_module.gprf[957] ;
 wire \reg_module.gprf[958] ;
 wire \reg_module.gprf[959] ;
 wire \reg_module.gprf[95] ;
 wire \reg_module.gprf[960] ;
 wire \reg_module.gprf[961] ;
 wire \reg_module.gprf[962] ;
 wire \reg_module.gprf[963] ;
 wire \reg_module.gprf[964] ;
 wire \reg_module.gprf[965] ;
 wire \reg_module.gprf[966] ;
 wire \reg_module.gprf[967] ;
 wire \reg_module.gprf[968] ;
 wire \reg_module.gprf[969] ;
 wire \reg_module.gprf[96] ;
 wire \reg_module.gprf[970] ;
 wire \reg_module.gprf[971] ;
 wire \reg_module.gprf[972] ;
 wire \reg_module.gprf[973] ;
 wire \reg_module.gprf[974] ;
 wire \reg_module.gprf[975] ;
 wire \reg_module.gprf[976] ;
 wire \reg_module.gprf[977] ;
 wire \reg_module.gprf[978] ;
 wire \reg_module.gprf[979] ;
 wire \reg_module.gprf[97] ;
 wire \reg_module.gprf[980] ;
 wire \reg_module.gprf[981] ;
 wire \reg_module.gprf[982] ;
 wire \reg_module.gprf[983] ;
 wire \reg_module.gprf[984] ;
 wire \reg_module.gprf[985] ;
 wire \reg_module.gprf[986] ;
 wire \reg_module.gprf[987] ;
 wire \reg_module.gprf[988] ;
 wire \reg_module.gprf[989] ;
 wire \reg_module.gprf[98] ;
 wire \reg_module.gprf[990] ;
 wire \reg_module.gprf[991] ;
 wire \reg_module.gprf[992] ;
 wire \reg_module.gprf[993] ;
 wire \reg_module.gprf[994] ;
 wire \reg_module.gprf[995] ;
 wire \reg_module.gprf[996] ;
 wire \reg_module.gprf[997] ;
 wire \reg_module.gprf[998] ;
 wire \reg_module.gprf[999] ;
 wire \reg_module.gprf[99] ;
 wire \reg_module.gprf[9] ;
 wire wRamByteEn;
 wire wRamHalfEn;
 wire wRamWordEn;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;

 sky130_fd_sc_hd__inv_2 _06118_ (.A(net156),
    .Y(_01203_));
 sky130_fd_sc_hd__inv_2 _06119_ (.A(net155),
    .Y(_01204_));
 sky130_fd_sc_hd__inv_2 _06120_ (.A(net154),
    .Y(_01205_));
 sky130_fd_sc_hd__inv_2 _06121_ (.A(net145),
    .Y(_01206_));
 sky130_fd_sc_hd__inv_2 _06122_ (.A(net953),
    .Y(_01207_));
 sky130_fd_sc_hd__clkinv_4 _06123_ (.A(net957),
    .Y(_01208_));
 sky130_fd_sc_hd__inv_2 _06124_ (.A(\alu.b_type ),
    .Y(_01209_));
 sky130_fd_sc_hd__inv_2 _06125_ (.A(net992),
    .Y(_01210_));
 sky130_fd_sc_hd__inv_2 _06126_ (.A(net984),
    .Y(_01211_));
 sky130_fd_sc_hd__inv_2 _06127_ (.A(net1066),
    .Y(_01212_));
 sky130_fd_sc_hd__inv_2 _06128_ (.A(\rReg_d2[0] ),
    .Y(_01213_));
 sky130_fd_sc_hd__inv_2 _06129_ (.A(net968),
    .Y(_01214_));
 sky130_fd_sc_hd__inv_2 _06130_ (.A(\rWrDataWB[31] ),
    .Y(_01215_));
 sky130_fd_sc_hd__inv_2 _06131_ (.A(\rReg_d[2] ),
    .Y(_01216_));
 sky130_fd_sc_hd__inv_2 _06132_ (.A(net845),
    .Y(_01217_));
 sky130_fd_sc_hd__inv_2 _06133_ (.A(net943),
    .Y(_01218_));
 sky130_fd_sc_hd__inv_2 _06134_ (.A(net944),
    .Y(_01219_));
 sky130_fd_sc_hd__inv_2 _06135_ (.A(net857),
    .Y(_01220_));
 sky130_fd_sc_hd__inv_2 _06136_ (.A(net848),
    .Y(_01221_));
 sky130_fd_sc_hd__inv_2 _06137_ (.A(net938),
    .Y(_01222_));
 sky130_fd_sc_hd__inv_2 _06138_ (.A(\brancher.imm12_i_s[10] ),
    .Y(_01223_));
 sky130_fd_sc_hd__inv_2 _06139_ (.A(\brancher.imm12_i_s[9] ),
    .Y(_01224_));
 sky130_fd_sc_hd__inv_2 _06140_ (.A(\brancher.imm12_i_s[7] ),
    .Y(_01225_));
 sky130_fd_sc_hd__inv_2 _06141_ (.A(\brancher.imm12_i_s[6] ),
    .Y(_01226_));
 sky130_fd_sc_hd__nor2_1 _06142_ (.A(net813),
    .B(net847),
    .Y(wRamWordEn));
 sky130_fd_sc_hd__nor2_1 _06143_ (.A(net846),
    .B(net847),
    .Y(wRamByteEn));
 sky130_fd_sc_hd__nand2_2 _06144_ (.A(net813),
    .B(net847),
    .Y(_01227_));
 sky130_fd_sc_hd__inv_2 _06145_ (.A(_01227_),
    .Y(wRamHalfEn));
 sky130_fd_sc_hd__xnor2_1 _06146_ (.A(net1046),
    .B(\rReg_d[0] ),
    .Y(_01228_));
 sky130_fd_sc_hd__or4_1 _06147_ (.A(\rReg_d[0] ),
    .B(\rReg_d[1] ),
    .C(\rReg_d[3] ),
    .D(\rReg_d[4] ),
    .X(_01229_));
 sky130_fd_sc_hd__nand2b_1 _06148_ (.A_N(net986),
    .B(\rReg_d[3] ),
    .Y(_01230_));
 sky130_fd_sc_hd__nand2b_1 _06149_ (.A_N(\rReg_d[3] ),
    .B(net986),
    .Y(_01231_));
 sky130_fd_sc_hd__xnor2_1 _06150_ (.A(net1067),
    .B(\rReg_d[4] ),
    .Y(_01232_));
 sky130_fd_sc_hd__xnor2_1 _06151_ (.A(net1012),
    .B(\rReg_d[1] ),
    .Y(_01233_));
 sky130_fd_sc_hd__o211a_1 _06152_ (.A1(net994),
    .A2(_01216_),
    .B1(_01230_),
    .C1(_01231_),
    .X(_01234_));
 sky130_fd_sc_hd__o211a_1 _06153_ (.A1(net827),
    .A2(\rReg_d[2] ),
    .B1(rRegWrEn),
    .C1(_01228_),
    .X(_01235_));
 sky130_fd_sc_hd__o211a_1 _06154_ (.A1(\rReg_d[2] ),
    .A2(_01229_),
    .B1(_01232_),
    .C1(_01233_),
    .X(_01236_));
 sky130_fd_sc_hd__and3_2 _06155_ (.A(_01234_),
    .B(_01235_),
    .C(_01236_),
    .X(_01237_));
 sky130_fd_sc_hd__nand3_4 _06156_ (.A(_01234_),
    .B(_01235_),
    .C(_01236_),
    .Y(_01238_));
 sky130_fd_sc_hd__or4bb_1 _06157_ (.A(rHazardStallRs1),
    .B(rHazardStallRs2),
    .C_N(rOp_memLd),
    .D_N(net1),
    .X(_01239_));
 sky130_fd_sc_hd__nor2_1 _06158_ (.A(net617),
    .B(_01239_),
    .Y(_00000_));
 sky130_fd_sc_hd__xnor2_1 _06159_ (.A(\rReg_d[0] ),
    .B(net917),
    .Y(_01240_));
 sky130_fd_sc_hd__xnor2_1 _06160_ (.A(\rReg_d[4] ),
    .B(net939),
    .Y(_01241_));
 sky130_fd_sc_hd__o211a_1 _06161_ (.A1(\rReg_d[2] ),
    .A2(_01229_),
    .B1(_01240_),
    .C1(_01241_),
    .X(_01242_));
 sky130_fd_sc_hd__nor2_1 _06162_ (.A(\rReg_d[1] ),
    .B(net880),
    .Y(_01243_));
 sky130_fd_sc_hd__and2_1 _06163_ (.A(\rReg_d[1] ),
    .B(net880),
    .X(_01244_));
 sky130_fd_sc_hd__o221a_1 _06164_ (.A1(\rReg_d[2] ),
    .A2(net802),
    .B1(_01243_),
    .B2(_01244_),
    .C1(rRegWrEn),
    .X(_01245_));
 sky130_fd_sc_hd__nand2b_1 _06165_ (.A_N(\rReg_d[3] ),
    .B(net851),
    .Y(_01246_));
 sky130_fd_sc_hd__nand2b_1 _06166_ (.A_N(net851),
    .B(\rReg_d[3] ),
    .Y(_01247_));
 sky130_fd_sc_hd__o211a_1 _06167_ (.A1(_01216_),
    .A2(net860),
    .B1(_01246_),
    .C1(_01247_),
    .X(_01248_));
 sky130_fd_sc_hd__and3_2 _06168_ (.A(_01242_),
    .B(_01245_),
    .C(_01248_),
    .X(_01249_));
 sky130_fd_sc_hd__nand3_4 _06169_ (.A(_01242_),
    .B(_01245_),
    .C(_01248_),
    .Y(_01250_));
 sky130_fd_sc_hd__nor2_1 _06170_ (.A(_01239_),
    .B(net603),
    .Y(_00001_));
 sky130_fd_sc_hd__nor2_1 _06171_ (.A(_00000_),
    .B(_00001_),
    .Y(_01251_));
 sky130_fd_sc_hd__inv_2 _06172_ (.A(net266),
    .Y(\brancher.stall ));
 sky130_fd_sc_hd__or2_1 _06173_ (.A(\rWrData[0] ),
    .B(net617),
    .X(_01252_));
 sky130_fd_sc_hd__nor3_1 _06174_ (.A(\rReg_d2[0] ),
    .B(net970),
    .C(net968),
    .Y(_01253_));
 sky130_fd_sc_hd__or4_2 _06175_ (.A(\rReg_d2[0] ),
    .B(net969),
    .C(net968),
    .D(net966),
    .X(_01254_));
 sky130_fd_sc_hd__a21o_1 _06176_ (.A1(net815),
    .A2(_01254_),
    .B1(\rReg_d2[4] ),
    .X(_01255_));
 sky130_fd_sc_hd__and2b_1 _06177_ (.A_N(net1012),
    .B(net969),
    .X(_01256_));
 sky130_fd_sc_hd__and2b_1 _06178_ (.A_N(net1067),
    .B(\rReg_d2[4] ),
    .X(_01257_));
 sky130_fd_sc_hd__and2b_1 _06179_ (.A_N(net969),
    .B(net1012),
    .X(_01258_));
 sky130_fd_sc_hd__a2111oi_1 _06180_ (.A1(net1046),
    .A2(_01213_),
    .B1(_01256_),
    .C1(_01257_),
    .D1(_01258_),
    .Y(_01259_));
 sky130_fd_sc_hd__xnor2_1 _06181_ (.A(net987),
    .B(net966),
    .Y(_01260_));
 sky130_fd_sc_hd__xnor2_1 _06182_ (.A(net994),
    .B(net968),
    .Y(_01261_));
 sky130_fd_sc_hd__o2111a_1 _06183_ (.A1(net1046),
    .A2(_01213_),
    .B1(rRegWrEn2),
    .C1(_01260_),
    .D1(_01261_),
    .X(_01262_));
 sky130_fd_sc_hd__a31oi_1 _06184_ (.A1(_01255_),
    .A2(_01259_),
    .A3(_01262_),
    .B1(rHazardStallRs1),
    .Y(_01263_));
 sky130_fd_sc_hd__a31o_2 _06185_ (.A1(_01255_),
    .A2(net744),
    .A3(_01262_),
    .B1(rHazardStallRs1),
    .X(_01264_));
 sky130_fd_sc_hd__mux4_1 _06186_ (.A0(\reg_module.gprf[352] ),
    .A1(\reg_module.gprf[320] ),
    .A2(\reg_module.gprf[288] ),
    .A3(\reg_module.gprf[256] ),
    .S0(net1044),
    .S1(net1010),
    .X(_01265_));
 sky130_fd_sc_hd__mux4_1 _06187_ (.A0(\reg_module.gprf[480] ),
    .A1(\reg_module.gprf[448] ),
    .A2(\reg_module.gprf[416] ),
    .A3(\reg_module.gprf[384] ),
    .S0(net1044),
    .S1(net1010),
    .X(_01266_));
 sky130_fd_sc_hd__mux4_1 _06188_ (.A0(\reg_module.gprf[96] ),
    .A1(\reg_module.gprf[64] ),
    .A2(\reg_module.gprf[32] ),
    .A3(\reg_module.gprf[0] ),
    .S0(net1035),
    .S1(net1001),
    .X(_01267_));
 sky130_fd_sc_hd__mux4_1 _06189_ (.A0(\reg_module.gprf[224] ),
    .A1(\reg_module.gprf[192] ),
    .A2(\reg_module.gprf[160] ),
    .A3(\reg_module.gprf[128] ),
    .S0(net1036),
    .S1(net1002),
    .X(_01268_));
 sky130_fd_sc_hd__mux4_1 _06190_ (.A0(_01265_),
    .A1(_01266_),
    .A2(_01267_),
    .A3(_01268_),
    .S0(net823),
    .S1(net985),
    .X(_01269_));
 sky130_fd_sc_hd__nand2_1 _06191_ (.A(net1066),
    .B(_01269_),
    .Y(_01270_));
 sky130_fd_sc_hd__mux4_1 _06192_ (.A0(\reg_module.gprf[864] ),
    .A1(\reg_module.gprf[832] ),
    .A2(\reg_module.gprf[800] ),
    .A3(\reg_module.gprf[768] ),
    .S0(net1044),
    .S1(net1010),
    .X(_01271_));
 sky130_fd_sc_hd__mux4_1 _06193_ (.A0(\reg_module.gprf[992] ),
    .A1(\reg_module.gprf[960] ),
    .A2(\reg_module.gprf[928] ),
    .A3(\reg_module.gprf[896] ),
    .S0(net1044),
    .S1(net1010),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _06194_ (.A0(_01271_),
    .A1(_01272_),
    .S(net827),
    .X(_01273_));
 sky130_fd_sc_hd__nor2_1 _06195_ (.A(net986),
    .B(_01273_),
    .Y(_01274_));
 sky130_fd_sc_hd__mux4_1 _06196_ (.A0(\reg_module.gprf[736] ),
    .A1(\reg_module.gprf[704] ),
    .A2(\reg_module.gprf[672] ),
    .A3(\reg_module.gprf[640] ),
    .S0(net1035),
    .S1(net1001),
    .X(_01275_));
 sky130_fd_sc_hd__mux4_1 _06197_ (.A0(\reg_module.gprf[608] ),
    .A1(\reg_module.gprf[576] ),
    .A2(\reg_module.gprf[544] ),
    .A3(\reg_module.gprf[512] ),
    .S0(net1041),
    .S1(net1007),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _06198_ (.A0(_01275_),
    .A1(_01276_),
    .S(net992),
    .X(_01277_));
 sky130_fd_sc_hd__o21ai_1 _06199_ (.A1(net820),
    .A2(_01277_),
    .B1(net815),
    .Y(_01278_));
 sky130_fd_sc_hd__o21ai_2 _06200_ (.A1(_01274_),
    .A2(_01278_),
    .B1(_01270_),
    .Y(_01279_));
 sky130_fd_sc_hd__o211a_1 _06201_ (.A1(_01274_),
    .A2(_01278_),
    .B1(net595),
    .C1(_01270_),
    .X(_01280_));
 sky130_fd_sc_hd__nor2_1 _06202_ (.A(\rWrDataWB[0] ),
    .B(net595),
    .Y(_01281_));
 sky130_fd_sc_hd__o21ai_1 _06203_ (.A1(_01280_),
    .A2(_01281_),
    .B1(net617),
    .Y(_01282_));
 sky130_fd_sc_hd__and3_1 _06204_ (.A(\brancher.imm12_i_s[0] ),
    .B(_01252_),
    .C(_01282_),
    .X(_01283_));
 sky130_fd_sc_hd__nor2_4 _06205_ (.A(\dec.op_memSt ),
    .B(\dec.op_memLd ),
    .Y(_01284_));
 sky130_fd_sc_hd__or2_1 _06206_ (.A(\dec.op_memSt ),
    .B(\dec.op_memLd ),
    .X(_01285_));
 sky130_fd_sc_hd__a21o_1 _06207_ (.A1(_01252_),
    .A2(_01282_),
    .B1(\brancher.imm12_i_s[0] ),
    .X(_01286_));
 sky130_fd_sc_hd__and3b_1 _06208_ (.A_N(_01283_),
    .B(net772),
    .C(_01286_),
    .X(net71));
 sky130_fd_sc_hd__and2_1 _06209_ (.A(\rWrData[1] ),
    .B(net623),
    .X(_01287_));
 sky130_fd_sc_hd__mux4_1 _06210_ (.A0(\reg_module.gprf[353] ),
    .A1(\reg_module.gprf[321] ),
    .A2(\reg_module.gprf[289] ),
    .A3(\reg_module.gprf[257] ),
    .S0(net1045),
    .S1(net1011),
    .X(_01288_));
 sky130_fd_sc_hd__mux4_1 _06211_ (.A0(\reg_module.gprf[481] ),
    .A1(\reg_module.gprf[449] ),
    .A2(\reg_module.gprf[417] ),
    .A3(\reg_module.gprf[385] ),
    .S0(net1046),
    .S1(net1012),
    .X(_01289_));
 sky130_fd_sc_hd__mux4_1 _06212_ (.A0(\reg_module.gprf[97] ),
    .A1(\reg_module.gprf[65] ),
    .A2(\reg_module.gprf[33] ),
    .A3(\reg_module.gprf[1] ),
    .S0(net1045),
    .S1(net1011),
    .X(_01290_));
 sky130_fd_sc_hd__mux4_1 _06213_ (.A0(\reg_module.gprf[225] ),
    .A1(\reg_module.gprf[193] ),
    .A2(\reg_module.gprf[161] ),
    .A3(\reg_module.gprf[129] ),
    .S0(net1046),
    .S1(net1011),
    .X(_01291_));
 sky130_fd_sc_hd__mux4_1 _06214_ (.A0(_01288_),
    .A1(_01289_),
    .A2(_01290_),
    .A3(_01291_),
    .S0(net827),
    .S1(net986),
    .X(_01292_));
 sky130_fd_sc_hd__nor2_1 _06215_ (.A(net815),
    .B(_01292_),
    .Y(_01293_));
 sky130_fd_sc_hd__mux4_1 _06216_ (.A0(\reg_module.gprf[609] ),
    .A1(\reg_module.gprf[577] ),
    .A2(\reg_module.gprf[545] ),
    .A3(\reg_module.gprf[513] ),
    .S0(net1047),
    .S1(net1013),
    .X(_01294_));
 sky130_fd_sc_hd__mux4_1 _06217_ (.A0(\reg_module.gprf[737] ),
    .A1(\reg_module.gprf[705] ),
    .A2(\reg_module.gprf[673] ),
    .A3(\reg_module.gprf[641] ),
    .S0(net1047),
    .S1(net1013),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _06218_ (.A0(_01294_),
    .A1(_01295_),
    .S(net827),
    .X(_01296_));
 sky130_fd_sc_hd__nand2_1 _06219_ (.A(net986),
    .B(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hd__mux4_1 _06220_ (.A0(\reg_module.gprf[865] ),
    .A1(\reg_module.gprf[833] ),
    .A2(\reg_module.gprf[801] ),
    .A3(\reg_module.gprf[769] ),
    .S0(net1045),
    .S1(net1011),
    .X(_01298_));
 sky130_fd_sc_hd__mux4_1 _06221_ (.A0(\reg_module.gprf[993] ),
    .A1(\reg_module.gprf[961] ),
    .A2(\reg_module.gprf[929] ),
    .A3(\reg_module.gprf[897] ),
    .S0(net1046),
    .S1(net1012),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _06222_ (.A0(_01298_),
    .A1(_01299_),
    .S(net827),
    .X(_01300_));
 sky130_fd_sc_hd__a21oi_1 _06223_ (.A1(net820),
    .A2(_01300_),
    .B1(net1067),
    .Y(_01301_));
 sky130_fd_sc_hd__a21oi_1 _06224_ (.A1(_01297_),
    .A2(_01301_),
    .B1(_01293_),
    .Y(_01302_));
 sky130_fd_sc_hd__a211o_1 _06225_ (.A1(_01297_),
    .A2(_01301_),
    .B1(net589),
    .C1(_01293_),
    .X(_01303_));
 sky130_fd_sc_hd__nand2_1 _06226_ (.A(\rWrDataWB[1] ),
    .B(net589),
    .Y(_01304_));
 sky130_fd_sc_hd__a21oi_1 _06227_ (.A1(_01303_),
    .A2(_01304_),
    .B1(net623),
    .Y(_01305_));
 sky130_fd_sc_hd__o21a_1 _06228_ (.A1(_01287_),
    .A2(_01305_),
    .B1(\brancher.imm12_i_s[1] ),
    .X(_01306_));
 sky130_fd_sc_hd__or3_1 _06229_ (.A(\brancher.imm12_i_s[1] ),
    .B(_01287_),
    .C(_01305_),
    .X(_01307_));
 sky130_fd_sc_hd__and2b_1 _06230_ (.A_N(_01306_),
    .B(_01307_),
    .X(_01308_));
 sky130_fd_sc_hd__o21ai_1 _06231_ (.A1(_01283_),
    .A2(_01308_),
    .B1(net772),
    .Y(_01309_));
 sky130_fd_sc_hd__a21oi_2 _06232_ (.A1(_01283_),
    .A2(_01308_),
    .B1(_01309_),
    .Y(net82));
 sky130_fd_sc_hd__or2_1 _06233_ (.A(\rWrData[2] ),
    .B(net618),
    .X(_01310_));
 sky130_fd_sc_hd__mux4_1 _06234_ (.A0(\reg_module.gprf[354] ),
    .A1(\reg_module.gprf[322] ),
    .A2(\reg_module.gprf[290] ),
    .A3(\reg_module.gprf[258] ),
    .S0(net1041),
    .S1(net1007),
    .X(_01311_));
 sky130_fd_sc_hd__mux4_1 _06235_ (.A0(\reg_module.gprf[482] ),
    .A1(\reg_module.gprf[450] ),
    .A2(\reg_module.gprf[418] ),
    .A3(\reg_module.gprf[386] ),
    .S0(net1041),
    .S1(net1007),
    .X(_01312_));
 sky130_fd_sc_hd__mux2_1 _06236_ (.A0(_01311_),
    .A1(_01312_),
    .S(net826),
    .X(_01313_));
 sky130_fd_sc_hd__mux4_1 _06237_ (.A0(\reg_module.gprf[98] ),
    .A1(\reg_module.gprf[66] ),
    .A2(\reg_module.gprf[34] ),
    .A3(\reg_module.gprf[2] ),
    .S0(net1041),
    .S1(net1007),
    .X(_01314_));
 sky130_fd_sc_hd__mux4_1 _06238_ (.A0(\reg_module.gprf[226] ),
    .A1(\reg_module.gprf[194] ),
    .A2(\reg_module.gprf[162] ),
    .A3(\reg_module.gprf[130] ),
    .S0(net1041),
    .S1(net1007),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _06239_ (.A0(_01314_),
    .A1(_01315_),
    .S(net826),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _06240_ (.A0(_01313_),
    .A1(_01316_),
    .S(net987),
    .X(_01317_));
 sky130_fd_sc_hd__mux4_1 _06241_ (.A0(\reg_module.gprf[610] ),
    .A1(\reg_module.gprf[578] ),
    .A2(\reg_module.gprf[546] ),
    .A3(\reg_module.gprf[514] ),
    .S0(net1035),
    .S1(net1001),
    .X(_01318_));
 sky130_fd_sc_hd__or2_1 _06242_ (.A(net824),
    .B(_01318_),
    .X(_01319_));
 sky130_fd_sc_hd__mux4_1 _06243_ (.A0(\reg_module.gprf[738] ),
    .A1(\reg_module.gprf[706] ),
    .A2(\reg_module.gprf[674] ),
    .A3(\reg_module.gprf[642] ),
    .S0(net1035),
    .S1(net1001),
    .X(_01320_));
 sky130_fd_sc_hd__o21a_1 _06244_ (.A1(net992),
    .A2(_01320_),
    .B1(net984),
    .X(_01321_));
 sky130_fd_sc_hd__mux4_1 _06245_ (.A0(\reg_module.gprf[866] ),
    .A1(\reg_module.gprf[834] ),
    .A2(\reg_module.gprf[802] ),
    .A3(\reg_module.gprf[770] ),
    .S0(net1041),
    .S1(net1007),
    .X(_01322_));
 sky130_fd_sc_hd__mux4_1 _06246_ (.A0(\reg_module.gprf[994] ),
    .A1(\reg_module.gprf[962] ),
    .A2(\reg_module.gprf[930] ),
    .A3(\reg_module.gprf[898] ),
    .S0(net1041),
    .S1(net1007),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _06247_ (.A0(_01322_),
    .A1(_01323_),
    .S(net824),
    .X(_01324_));
 sky130_fd_sc_hd__a221o_1 _06248_ (.A1(_01319_),
    .A2(_01321_),
    .B1(_01324_),
    .B2(net818),
    .C1(net1066),
    .X(_01325_));
 sky130_fd_sc_hd__o21a_2 _06249_ (.A1(net815),
    .A2(_01317_),
    .B1(_01325_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _06250_ (.A0(\rWrDataWB[2] ),
    .A1(_01326_),
    .S(net597),
    .X(_01327_));
 sky130_fd_sc_hd__o21a_1 _06251_ (.A1(net623),
    .A2(_01327_),
    .B1(_01310_),
    .X(_01328_));
 sky130_fd_sc_hd__nand2_1 _06252_ (.A(\brancher.imm12_i_s[2] ),
    .B(_01328_),
    .Y(_01329_));
 sky130_fd_sc_hd__xnor2_1 _06253_ (.A(\brancher.imm12_i_s[2] ),
    .B(_01328_),
    .Y(_01330_));
 sky130_fd_sc_hd__a21oi_1 _06254_ (.A1(_01283_),
    .A2(_01307_),
    .B1(_01306_),
    .Y(_01331_));
 sky130_fd_sc_hd__xnor2_1 _06255_ (.A(_01330_),
    .B(_01331_),
    .Y(_01332_));
 sky130_fd_sc_hd__nor2_1 _06256_ (.A(net773),
    .B(_01332_),
    .Y(net93));
 sky130_fd_sc_hd__mux4_1 _06257_ (.A0(\reg_module.gprf[355] ),
    .A1(\reg_module.gprf[323] ),
    .A2(\reg_module.gprf[291] ),
    .A3(\reg_module.gprf[259] ),
    .S0(net1035),
    .S1(net1001),
    .X(_01333_));
 sky130_fd_sc_hd__mux4_1 _06258_ (.A0(\reg_module.gprf[483] ),
    .A1(\reg_module.gprf[451] ),
    .A2(\reg_module.gprf[419] ),
    .A3(\reg_module.gprf[387] ),
    .S0(net1035),
    .S1(net1001),
    .X(_01334_));
 sky130_fd_sc_hd__mux4_1 _06259_ (.A0(\reg_module.gprf[99] ),
    .A1(\reg_module.gprf[67] ),
    .A2(\reg_module.gprf[35] ),
    .A3(\reg_module.gprf[3] ),
    .S0(net1032),
    .S1(net998),
    .X(_01335_));
 sky130_fd_sc_hd__mux4_1 _06260_ (.A0(\reg_module.gprf[227] ),
    .A1(\reg_module.gprf[195] ),
    .A2(\reg_module.gprf[163] ),
    .A3(\reg_module.gprf[131] ),
    .S0(net1036),
    .S1(net1002),
    .X(_01336_));
 sky130_fd_sc_hd__mux4_1 _06261_ (.A0(_01333_),
    .A1(_01334_),
    .A2(_01335_),
    .A3(_01336_),
    .S0(net823),
    .S1(net984),
    .X(_01337_));
 sky130_fd_sc_hd__mux4_1 _06262_ (.A0(\reg_module.gprf[867] ),
    .A1(\reg_module.gprf[835] ),
    .A2(\reg_module.gprf[803] ),
    .A3(\reg_module.gprf[771] ),
    .S0(net1035),
    .S1(net1001),
    .X(_01338_));
 sky130_fd_sc_hd__or2_1 _06263_ (.A(net824),
    .B(_01338_),
    .X(_01339_));
 sky130_fd_sc_hd__mux4_1 _06264_ (.A0(\reg_module.gprf[995] ),
    .A1(\reg_module.gprf[963] ),
    .A2(\reg_module.gprf[931] ),
    .A3(\reg_module.gprf[899] ),
    .S0(net1035),
    .S1(net1001),
    .X(_01340_));
 sky130_fd_sc_hd__o21a_1 _06265_ (.A1(net993),
    .A2(_01340_),
    .B1(net818),
    .X(_01341_));
 sky130_fd_sc_hd__mux4_1 _06266_ (.A0(\reg_module.gprf[739] ),
    .A1(\reg_module.gprf[707] ),
    .A2(\reg_module.gprf[675] ),
    .A3(\reg_module.gprf[643] ),
    .S0(net1035),
    .S1(net1001),
    .X(_01342_));
 sky130_fd_sc_hd__mux4_1 _06267_ (.A0(\reg_module.gprf[611] ),
    .A1(\reg_module.gprf[579] ),
    .A2(\reg_module.gprf[547] ),
    .A3(\reg_module.gprf[515] ),
    .S0(net1035),
    .S1(net1001),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _06268_ (.A0(_01342_),
    .A1(_01343_),
    .S(net993),
    .X(_01344_));
 sky130_fd_sc_hd__a221o_1 _06269_ (.A1(_01339_),
    .A2(_01341_),
    .B1(_01344_),
    .B2(net984),
    .C1(net1066),
    .X(_01345_));
 sky130_fd_sc_hd__o21a_2 _06270_ (.A1(net814),
    .A2(_01337_),
    .B1(_01345_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _06271_ (.A0(\rWrDataWB[3] ),
    .A1(_01346_),
    .S(net595),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _06272_ (.A0(\rWrData[3] ),
    .A1(_01347_),
    .S(net617),
    .X(_01348_));
 sky130_fd_sc_hd__nand2_1 _06273_ (.A(\brancher.imm12_i_s[3] ),
    .B(_01348_),
    .Y(_01349_));
 sky130_fd_sc_hd__or2_1 _06274_ (.A(\brancher.imm12_i_s[3] ),
    .B(_01348_),
    .X(_01350_));
 sky130_fd_sc_hd__nand2_1 _06275_ (.A(_01349_),
    .B(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__o21a_1 _06276_ (.A1(_01330_),
    .A2(_01331_),
    .B1(_01329_),
    .X(_01352_));
 sky130_fd_sc_hd__o21ai_1 _06277_ (.A1(_01351_),
    .A2(_01352_),
    .B1(net772),
    .Y(_01353_));
 sky130_fd_sc_hd__a21oi_1 _06278_ (.A1(_01351_),
    .A2(_01352_),
    .B1(_01353_),
    .Y(net96));
 sky130_fd_sc_hd__mux4_1 _06279_ (.A0(\reg_module.gprf[356] ),
    .A1(\reg_module.gprf[324] ),
    .A2(\reg_module.gprf[292] ),
    .A3(\reg_module.gprf[260] ),
    .S0(net1045),
    .S1(net1011),
    .X(_01354_));
 sky130_fd_sc_hd__mux4_1 _06280_ (.A0(\reg_module.gprf[484] ),
    .A1(\reg_module.gprf[452] ),
    .A2(\reg_module.gprf[420] ),
    .A3(\reg_module.gprf[388] ),
    .S0(net1045),
    .S1(net1012),
    .X(_01355_));
 sky130_fd_sc_hd__mux4_1 _06281_ (.A0(\reg_module.gprf[100] ),
    .A1(\reg_module.gprf[68] ),
    .A2(\reg_module.gprf[36] ),
    .A3(\reg_module.gprf[4] ),
    .S0(net1045),
    .S1(net1011),
    .X(_01356_));
 sky130_fd_sc_hd__mux4_1 _06282_ (.A0(\reg_module.gprf[228] ),
    .A1(\reg_module.gprf[196] ),
    .A2(\reg_module.gprf[164] ),
    .A3(\reg_module.gprf[132] ),
    .S0(net1045),
    .S1(net1011),
    .X(_01357_));
 sky130_fd_sc_hd__mux4_1 _06283_ (.A0(_01354_),
    .A1(_01355_),
    .A2(_01356_),
    .A3(_01357_),
    .S0(net828),
    .S1(net986),
    .X(_01358_));
 sky130_fd_sc_hd__mux4_1 _06284_ (.A0(\reg_module.gprf[868] ),
    .A1(\reg_module.gprf[836] ),
    .A2(\reg_module.gprf[804] ),
    .A3(\reg_module.gprf[772] ),
    .S0(net1046),
    .S1(net1012),
    .X(_01359_));
 sky130_fd_sc_hd__or2_1 _06285_ (.A(net827),
    .B(_01359_),
    .X(_01360_));
 sky130_fd_sc_hd__mux4_1 _06286_ (.A0(\reg_module.gprf[996] ),
    .A1(\reg_module.gprf[964] ),
    .A2(\reg_module.gprf[932] ),
    .A3(\reg_module.gprf[900] ),
    .S0(net1046),
    .S1(net1012),
    .X(_01361_));
 sky130_fd_sc_hd__o211a_1 _06287_ (.A1(net994),
    .A2(_01361_),
    .B1(_01360_),
    .C1(net820),
    .X(_01362_));
 sky130_fd_sc_hd__mux4_1 _06288_ (.A0(\reg_module.gprf[740] ),
    .A1(\reg_module.gprf[708] ),
    .A2(\reg_module.gprf[676] ),
    .A3(\reg_module.gprf[644] ),
    .S0(net1045),
    .S1(net1011),
    .X(_01363_));
 sky130_fd_sc_hd__mux4_1 _06289_ (.A0(\reg_module.gprf[612] ),
    .A1(\reg_module.gprf[580] ),
    .A2(\reg_module.gprf[548] ),
    .A3(\reg_module.gprf[516] ),
    .S0(net1045),
    .S1(net1011),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _06290_ (.A0(_01363_),
    .A1(_01364_),
    .S(net994),
    .X(_01365_));
 sky130_fd_sc_hd__a21o_1 _06291_ (.A1(net986),
    .A2(_01365_),
    .B1(net1067),
    .X(_01366_));
 sky130_fd_sc_hd__o22a_1 _06292_ (.A1(net815),
    .A2(_01358_),
    .B1(_01362_),
    .B2(_01366_),
    .X(_01367_));
 sky130_fd_sc_hd__o221a_1 _06293_ (.A1(net815),
    .A2(_01358_),
    .B1(_01362_),
    .B2(_01366_),
    .C1(net595),
    .X(_01368_));
 sky130_fd_sc_hd__a21o_1 _06294_ (.A1(\rWrDataWB[4] ),
    .A2(net589),
    .B1(net624),
    .X(_01369_));
 sky130_fd_sc_hd__o22a_1 _06295_ (.A1(\rWrData[4] ),
    .A2(net617),
    .B1(_01368_),
    .B2(_01369_),
    .X(_01370_));
 sky130_fd_sc_hd__nand2_1 _06296_ (.A(\brancher.imm12_i_s[4] ),
    .B(_01370_),
    .Y(_01371_));
 sky130_fd_sc_hd__or2_1 _06297_ (.A(\brancher.imm12_i_s[4] ),
    .B(_01370_),
    .X(_01372_));
 sky130_fd_sc_hd__nand2_1 _06298_ (.A(_01371_),
    .B(_01372_),
    .Y(_01373_));
 sky130_fd_sc_hd__o21a_1 _06299_ (.A1(_01351_),
    .A2(_01352_),
    .B1(_01349_),
    .X(_01374_));
 sky130_fd_sc_hd__o21ai_1 _06300_ (.A1(_01373_),
    .A2(_01374_),
    .B1(net772),
    .Y(_01375_));
 sky130_fd_sc_hd__a21oi_1 _06301_ (.A1(_01373_),
    .A2(_01374_),
    .B1(_01375_),
    .Y(net97));
 sky130_fd_sc_hd__mux4_1 _06302_ (.A0(\reg_module.gprf[357] ),
    .A1(\reg_module.gprf[325] ),
    .A2(\reg_module.gprf[293] ),
    .A3(\reg_module.gprf[261] ),
    .S0(net1043),
    .S1(net1009),
    .X(_01376_));
 sky130_fd_sc_hd__mux4_1 _06303_ (.A0(\reg_module.gprf[485] ),
    .A1(\reg_module.gprf[453] ),
    .A2(\reg_module.gprf[421] ),
    .A3(\reg_module.gprf[389] ),
    .S0(net1043),
    .S1(net1009),
    .X(_01377_));
 sky130_fd_sc_hd__mux4_1 _06304_ (.A0(\reg_module.gprf[101] ),
    .A1(\reg_module.gprf[69] ),
    .A2(\reg_module.gprf[37] ),
    .A3(\reg_module.gprf[5] ),
    .S0(net1043),
    .S1(net1009),
    .X(_01378_));
 sky130_fd_sc_hd__mux4_1 _06305_ (.A0(\reg_module.gprf[229] ),
    .A1(\reg_module.gprf[197] ),
    .A2(\reg_module.gprf[165] ),
    .A3(\reg_module.gprf[133] ),
    .S0(net1043),
    .S1(net1009),
    .X(_01379_));
 sky130_fd_sc_hd__mux4_1 _06306_ (.A0(_01376_),
    .A1(_01377_),
    .A2(_01378_),
    .A3(_01379_),
    .S0(net827),
    .S1(net986),
    .X(_01380_));
 sky130_fd_sc_hd__mux4_1 _06307_ (.A0(\reg_module.gprf[869] ),
    .A1(\reg_module.gprf[837] ),
    .A2(\reg_module.gprf[805] ),
    .A3(\reg_module.gprf[773] ),
    .S0(net1043),
    .S1(net1009),
    .X(_01381_));
 sky130_fd_sc_hd__mux4_1 _06308_ (.A0(\reg_module.gprf[997] ),
    .A1(\reg_module.gprf[965] ),
    .A2(\reg_module.gprf[933] ),
    .A3(\reg_module.gprf[901] ),
    .S0(net1043),
    .S1(net1009),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _06309_ (.A0(_01381_),
    .A1(_01382_),
    .S(net827),
    .X(_01383_));
 sky130_fd_sc_hd__mux4_1 _06310_ (.A0(\reg_module.gprf[741] ),
    .A1(\reg_module.gprf[709] ),
    .A2(\reg_module.gprf[677] ),
    .A3(\reg_module.gprf[645] ),
    .S0(net1034),
    .S1(net1000),
    .X(_01384_));
 sky130_fd_sc_hd__mux4_1 _06311_ (.A0(\reg_module.gprf[613] ),
    .A1(\reg_module.gprf[581] ),
    .A2(\reg_module.gprf[549] ),
    .A3(\reg_module.gprf[517] ),
    .S0(net1043),
    .S1(net1009),
    .X(_01385_));
 sky130_fd_sc_hd__or2_1 _06312_ (.A(net824),
    .B(_01385_),
    .X(_01386_));
 sky130_fd_sc_hd__o211a_1 _06313_ (.A1(net992),
    .A2(_01384_),
    .B1(_01386_),
    .C1(net985),
    .X(_01387_));
 sky130_fd_sc_hd__a21o_1 _06314_ (.A1(net820),
    .A2(_01383_),
    .B1(net1067),
    .X(_01388_));
 sky130_fd_sc_hd__o22a_1 _06315_ (.A1(net815),
    .A2(_01380_),
    .B1(_01387_),
    .B2(_01388_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _06316_ (.A0(\rWrDataWB[5] ),
    .A1(_01389_),
    .S(net595),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _06317_ (.A0(\rWrData[5] ),
    .A1(_01390_),
    .S(net616),
    .X(_01391_));
 sky130_fd_sc_hd__nand2_1 _06318_ (.A(\brancher.imm12_i_s[5] ),
    .B(_01391_),
    .Y(_01392_));
 sky130_fd_sc_hd__or2_1 _06319_ (.A(\brancher.imm12_i_s[5] ),
    .B(_01391_),
    .X(_01393_));
 sky130_fd_sc_hd__nand2_1 _06320_ (.A(_01392_),
    .B(_01393_),
    .Y(_01394_));
 sky130_fd_sc_hd__o21a_1 _06321_ (.A1(_01373_),
    .A2(_01374_),
    .B1(_01371_),
    .X(_01395_));
 sky130_fd_sc_hd__o21ai_1 _06322_ (.A1(_01394_),
    .A2(_01395_),
    .B1(net772),
    .Y(_01396_));
 sky130_fd_sc_hd__a21oi_1 _06323_ (.A1(_01394_),
    .A2(_01395_),
    .B1(_01396_),
    .Y(net98));
 sky130_fd_sc_hd__mux4_1 _06324_ (.A0(\reg_module.gprf[230] ),
    .A1(\reg_module.gprf[198] ),
    .A2(\reg_module.gprf[166] ),
    .A3(\reg_module.gprf[134] ),
    .S0(net1033),
    .S1(net999),
    .X(_01397_));
 sky130_fd_sc_hd__mux4_1 _06325_ (.A0(\reg_module.gprf[102] ),
    .A1(\reg_module.gprf[70] ),
    .A2(\reg_module.gprf[38] ),
    .A3(\reg_module.gprf[6] ),
    .S0(net1033),
    .S1(net999),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _06326_ (.A0(_01397_),
    .A1(_01398_),
    .S(net992),
    .X(_01399_));
 sky130_fd_sc_hd__mux4_1 _06327_ (.A0(\reg_module.gprf[358] ),
    .A1(\reg_module.gprf[326] ),
    .A2(\reg_module.gprf[294] ),
    .A3(\reg_module.gprf[262] ),
    .S0(net1033),
    .S1(net999),
    .X(_01400_));
 sky130_fd_sc_hd__mux4_1 _06328_ (.A0(\reg_module.gprf[486] ),
    .A1(\reg_module.gprf[454] ),
    .A2(\reg_module.gprf[422] ),
    .A3(\reg_module.gprf[390] ),
    .S0(net1033),
    .S1(net999),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _06329_ (.A0(_01400_),
    .A1(_01401_),
    .S(net823),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _06330_ (.A0(_01399_),
    .A1(_01402_),
    .S(net818),
    .X(_01403_));
 sky130_fd_sc_hd__mux4_1 _06331_ (.A0(\reg_module.gprf[870] ),
    .A1(\reg_module.gprf[838] ),
    .A2(\reg_module.gprf[806] ),
    .A3(\reg_module.gprf[774] ),
    .S0(net1034),
    .S1(net1000),
    .X(_01404_));
 sky130_fd_sc_hd__mux4_1 _06332_ (.A0(\reg_module.gprf[998] ),
    .A1(\reg_module.gprf[966] ),
    .A2(\reg_module.gprf[934] ),
    .A3(\reg_module.gprf[902] ),
    .S0(net1034),
    .S1(net1000),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _06333_ (.A0(_01404_),
    .A1(_01405_),
    .S(net824),
    .X(_01406_));
 sky130_fd_sc_hd__mux4_1 _06334_ (.A0(\reg_module.gprf[742] ),
    .A1(\reg_module.gprf[710] ),
    .A2(\reg_module.gprf[678] ),
    .A3(\reg_module.gprf[646] ),
    .S0(net1033),
    .S1(net999),
    .X(_01407_));
 sky130_fd_sc_hd__mux4_1 _06335_ (.A0(\reg_module.gprf[614] ),
    .A1(\reg_module.gprf[582] ),
    .A2(\reg_module.gprf[550] ),
    .A3(\reg_module.gprf[518] ),
    .S0(net1033),
    .S1(net999),
    .X(_01408_));
 sky130_fd_sc_hd__mux2_1 _06336_ (.A0(_01407_),
    .A1(_01408_),
    .S(net992),
    .X(_01409_));
 sky130_fd_sc_hd__nand2_1 _06337_ (.A(net984),
    .B(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hd__a21oi_1 _06338_ (.A1(net818),
    .A2(_01406_),
    .B1(net1066),
    .Y(_01411_));
 sky130_fd_sc_hd__a2bb2o_2 _06339_ (.A1_N(net814),
    .A2_N(_01403_),
    .B1(_01410_),
    .B2(_01411_),
    .X(_01412_));
 sky130_fd_sc_hd__nor2_1 _06340_ (.A(net587),
    .B(_01412_),
    .Y(_01413_));
 sky130_fd_sc_hd__a21o_1 _06341_ (.A1(\rWrDataWB[6] ),
    .A2(net587),
    .B1(net622),
    .X(_01414_));
 sky130_fd_sc_hd__o22a_1 _06342_ (.A1(\rWrData[6] ),
    .A2(net616),
    .B1(_01413_),
    .B2(_01414_),
    .X(_01415_));
 sky130_fd_sc_hd__nand2_1 _06343_ (.A(\brancher.imm12_i_s[6] ),
    .B(_01415_),
    .Y(_01416_));
 sky130_fd_sc_hd__or2_1 _06344_ (.A(\brancher.imm12_i_s[6] ),
    .B(_01415_),
    .X(_01417_));
 sky130_fd_sc_hd__nand2_1 _06345_ (.A(_01416_),
    .B(_01417_),
    .Y(_01418_));
 sky130_fd_sc_hd__o21a_1 _06346_ (.A1(_01394_),
    .A2(_01395_),
    .B1(_01392_),
    .X(_01419_));
 sky130_fd_sc_hd__a21o_1 _06347_ (.A1(_01418_),
    .A2(_01419_),
    .B1(net773),
    .X(_01420_));
 sky130_fd_sc_hd__o21ba_1 _06348_ (.A1(_01418_),
    .A2(_01419_),
    .B1_N(_01420_),
    .X(net99));
 sky130_fd_sc_hd__mux4_1 _06349_ (.A0(\reg_module.gprf[359] ),
    .A1(\reg_module.gprf[327] ),
    .A2(\reg_module.gprf[295] ),
    .A3(\reg_module.gprf[263] ),
    .S0(net1034),
    .S1(net1002),
    .X(_01421_));
 sky130_fd_sc_hd__mux4_1 _06350_ (.A0(\reg_module.gprf[487] ),
    .A1(\reg_module.gprf[455] ),
    .A2(\reg_module.gprf[423] ),
    .A3(\reg_module.gprf[391] ),
    .S0(net1034),
    .S1(net1000),
    .X(_01422_));
 sky130_fd_sc_hd__or2_1 _06351_ (.A(net992),
    .B(_01422_),
    .X(_01423_));
 sky130_fd_sc_hd__o21a_1 _06352_ (.A1(net824),
    .A2(_01421_),
    .B1(net818),
    .X(_01424_));
 sky130_fd_sc_hd__mux4_1 _06353_ (.A0(\reg_module.gprf[103] ),
    .A1(\reg_module.gprf[71] ),
    .A2(\reg_module.gprf[39] ),
    .A3(\reg_module.gprf[7] ),
    .S0(net1034),
    .S1(net1000),
    .X(_01425_));
 sky130_fd_sc_hd__mux4_1 _06354_ (.A0(\reg_module.gprf[231] ),
    .A1(\reg_module.gprf[199] ),
    .A2(\reg_module.gprf[167] ),
    .A3(\reg_module.gprf[135] ),
    .S0(net1034),
    .S1(net1000),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _06355_ (.A0(_01425_),
    .A1(_01426_),
    .S(net824),
    .X(_01427_));
 sky130_fd_sc_hd__a221o_1 _06356_ (.A1(_01423_),
    .A2(_01424_),
    .B1(_01427_),
    .B2(net984),
    .C1(net814),
    .X(_01428_));
 sky130_fd_sc_hd__mux4_1 _06357_ (.A0(\reg_module.gprf[615] ),
    .A1(\reg_module.gprf[583] ),
    .A2(\reg_module.gprf[551] ),
    .A3(\reg_module.gprf[519] ),
    .S0(net1034),
    .S1(net1000),
    .X(_01429_));
 sky130_fd_sc_hd__or2_1 _06358_ (.A(net824),
    .B(_01429_),
    .X(_01430_));
 sky130_fd_sc_hd__mux4_1 _06359_ (.A0(\reg_module.gprf[743] ),
    .A1(\reg_module.gprf[711] ),
    .A2(\reg_module.gprf[679] ),
    .A3(\reg_module.gprf[647] ),
    .S0(net1036),
    .S1(net1000),
    .X(_01431_));
 sky130_fd_sc_hd__o21a_1 _06360_ (.A1(net993),
    .A2(_01431_),
    .B1(net984),
    .X(_01432_));
 sky130_fd_sc_hd__mux4_1 _06361_ (.A0(\reg_module.gprf[871] ),
    .A1(\reg_module.gprf[839] ),
    .A2(\reg_module.gprf[807] ),
    .A3(\reg_module.gprf[775] ),
    .S0(net1034),
    .S1(net1000),
    .X(_01433_));
 sky130_fd_sc_hd__mux4_1 _06362_ (.A0(\reg_module.gprf[999] ),
    .A1(\reg_module.gprf[967] ),
    .A2(\reg_module.gprf[935] ),
    .A3(\reg_module.gprf[903] ),
    .S0(net1034),
    .S1(net1000),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _06363_ (.A0(_01433_),
    .A1(_01434_),
    .S(net824),
    .X(_01435_));
 sky130_fd_sc_hd__a221o_1 _06364_ (.A1(_01430_),
    .A2(_01432_),
    .B1(_01435_),
    .B2(net818),
    .C1(net1066),
    .X(_01436_));
 sky130_fd_sc_hd__nand2_1 _06365_ (.A(_01428_),
    .B(_01436_),
    .Y(_01437_));
 sky130_fd_sc_hd__and3_1 _06366_ (.A(net595),
    .B(_01428_),
    .C(_01436_),
    .X(_01438_));
 sky130_fd_sc_hd__a21o_1 _06367_ (.A1(\rWrDataWB[7] ),
    .A2(net587),
    .B1(net622),
    .X(_01439_));
 sky130_fd_sc_hd__o22a_1 _06368_ (.A1(\rWrData[7] ),
    .A2(net616),
    .B1(_01438_),
    .B2(_01439_),
    .X(_01440_));
 sky130_fd_sc_hd__and2_1 _06369_ (.A(\brancher.imm12_i_s[7] ),
    .B(_01440_),
    .X(_01441_));
 sky130_fd_sc_hd__nor2_1 _06370_ (.A(\brancher.imm12_i_s[7] ),
    .B(_01440_),
    .Y(_01442_));
 sky130_fd_sc_hd__or2_1 _06371_ (.A(_01441_),
    .B(_01442_),
    .X(_01443_));
 sky130_fd_sc_hd__o21a_1 _06372_ (.A1(_01418_),
    .A2(_01419_),
    .B1(_01416_),
    .X(_01444_));
 sky130_fd_sc_hd__a21o_1 _06373_ (.A1(_01443_),
    .A2(_01444_),
    .B1(net773),
    .X(_01445_));
 sky130_fd_sc_hd__o21ba_1 _06374_ (.A1(_01443_),
    .A2(_01444_),
    .B1_N(_01445_),
    .X(net100));
 sky130_fd_sc_hd__or2_2 _06375_ (.A(\rWrData[8] ),
    .B(net617),
    .X(_01446_));
 sky130_fd_sc_hd__mux4_1 _06376_ (.A0(\reg_module.gprf[360] ),
    .A1(\reg_module.gprf[328] ),
    .A2(\reg_module.gprf[296] ),
    .A3(\reg_module.gprf[264] ),
    .S0(net1043),
    .S1(net1010),
    .X(_01447_));
 sky130_fd_sc_hd__mux4_1 _06377_ (.A0(\reg_module.gprf[488] ),
    .A1(\reg_module.gprf[456] ),
    .A2(\reg_module.gprf[424] ),
    .A3(\reg_module.gprf[392] ),
    .S0(net1044),
    .S1(net1009),
    .X(_01448_));
 sky130_fd_sc_hd__mux4_1 _06378_ (.A0(\reg_module.gprf[104] ),
    .A1(\reg_module.gprf[72] ),
    .A2(\reg_module.gprf[40] ),
    .A3(\reg_module.gprf[8] ),
    .S0(net1044),
    .S1(net1009),
    .X(_01449_));
 sky130_fd_sc_hd__mux4_1 _06379_ (.A0(\reg_module.gprf[232] ),
    .A1(\reg_module.gprf[200] ),
    .A2(\reg_module.gprf[168] ),
    .A3(\reg_module.gprf[136] ),
    .S0(net1044),
    .S1(net1010),
    .X(_01450_));
 sky130_fd_sc_hd__mux4_1 _06380_ (.A0(_01447_),
    .A1(_01448_),
    .A2(_01449_),
    .A3(_01450_),
    .S0(net827),
    .S1(net986),
    .X(_01451_));
 sky130_fd_sc_hd__mux4_1 _06381_ (.A0(\reg_module.gprf[872] ),
    .A1(\reg_module.gprf[840] ),
    .A2(\reg_module.gprf[808] ),
    .A3(\reg_module.gprf[776] ),
    .S0(net1045),
    .S1(net1011),
    .X(_01452_));
 sky130_fd_sc_hd__or2_1 _06382_ (.A(net827),
    .B(_01452_),
    .X(_01453_));
 sky130_fd_sc_hd__mux4_1 _06383_ (.A0(\reg_module.gprf[1000] ),
    .A1(\reg_module.gprf[968] ),
    .A2(\reg_module.gprf[936] ),
    .A3(\reg_module.gprf[904] ),
    .S0(net1043),
    .S1(net1010),
    .X(_01454_));
 sky130_fd_sc_hd__o21a_1 _06384_ (.A1(\brancher.imm21_j[17] ),
    .A2(_01454_),
    .B1(net820),
    .X(_01455_));
 sky130_fd_sc_hd__mux4_1 _06385_ (.A0(\reg_module.gprf[744] ),
    .A1(\reg_module.gprf[712] ),
    .A2(\reg_module.gprf[680] ),
    .A3(\reg_module.gprf[648] ),
    .S0(net1043),
    .S1(net1009),
    .X(_01456_));
 sky130_fd_sc_hd__mux4_1 _06386_ (.A0(\reg_module.gprf[616] ),
    .A1(\reg_module.gprf[584] ),
    .A2(\reg_module.gprf[552] ),
    .A3(\reg_module.gprf[520] ),
    .S0(net1044),
    .S1(net1010),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _06387_ (.A0(_01456_),
    .A1(_01457_),
    .S(\brancher.imm21_j[17] ),
    .X(_01458_));
 sky130_fd_sc_hd__a221o_1 _06388_ (.A1(_01453_),
    .A2(_01455_),
    .B1(_01458_),
    .B2(net987),
    .C1(net1070),
    .X(_01459_));
 sky130_fd_sc_hd__o21a_1 _06389_ (.A1(net815),
    .A2(_01451_),
    .B1(_01459_),
    .X(_01460_));
 sky130_fd_sc_hd__o211a_1 _06390_ (.A1(net815),
    .A2(_01451_),
    .B1(_01459_),
    .C1(net595),
    .X(_01461_));
 sky130_fd_sc_hd__a21o_1 _06391_ (.A1(\rWrDataWB[8] ),
    .A2(net589),
    .B1(net623),
    .X(_01462_));
 sky130_fd_sc_hd__o21a_1 _06392_ (.A1(_01461_),
    .A2(_01462_),
    .B1(_01446_),
    .X(_01463_));
 sky130_fd_sc_hd__nand2_1 _06393_ (.A(\brancher.imm12_i_s[8] ),
    .B(_01463_),
    .Y(_01464_));
 sky130_fd_sc_hd__or2_1 _06394_ (.A(\brancher.imm12_i_s[8] ),
    .B(_01463_),
    .X(_01465_));
 sky130_fd_sc_hd__nand2_1 _06395_ (.A(_01464_),
    .B(_01465_),
    .Y(_01466_));
 sky130_fd_sc_hd__o21ba_1 _06396_ (.A1(_01442_),
    .A2(_01444_),
    .B1_N(_01441_),
    .X(_01467_));
 sky130_fd_sc_hd__a21oi_1 _06397_ (.A1(_01466_),
    .A2(_01467_),
    .B1(net773),
    .Y(_01468_));
 sky130_fd_sc_hd__o21a_1 _06398_ (.A1(_01466_),
    .A2(_01467_),
    .B1(_01468_),
    .X(net101));
 sky130_fd_sc_hd__or2_2 _06399_ (.A(\rWrData[9] ),
    .B(net616),
    .X(_01469_));
 sky130_fd_sc_hd__mux4_1 _06400_ (.A0(\reg_module.gprf[233] ),
    .A1(\reg_module.gprf[201] ),
    .A2(\reg_module.gprf[169] ),
    .A3(\reg_module.gprf[137] ),
    .S0(net1037),
    .S1(net1003),
    .X(_01470_));
 sky130_fd_sc_hd__mux4_1 _06401_ (.A0(\reg_module.gprf[105] ),
    .A1(\reg_module.gprf[73] ),
    .A2(\reg_module.gprf[41] ),
    .A3(\reg_module.gprf[9] ),
    .S0(net1037),
    .S1(net1003),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _06402_ (.A0(_01470_),
    .A1(_01471_),
    .S(net994),
    .X(_01472_));
 sky130_fd_sc_hd__mux4_1 _06403_ (.A0(\reg_module.gprf[361] ),
    .A1(\reg_module.gprf[329] ),
    .A2(\reg_module.gprf[297] ),
    .A3(\reg_module.gprf[265] ),
    .S0(net1037),
    .S1(net1003),
    .X(_01473_));
 sky130_fd_sc_hd__mux4_1 _06404_ (.A0(\reg_module.gprf[489] ),
    .A1(\reg_module.gprf[457] ),
    .A2(\reg_module.gprf[425] ),
    .A3(\reg_module.gprf[393] ),
    .S0(net1032),
    .S1(net998),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _06405_ (.A0(_01473_),
    .A1(_01474_),
    .S(net823),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _06406_ (.A0(_01472_),
    .A1(_01475_),
    .S(net818),
    .X(_01476_));
 sky130_fd_sc_hd__mux4_1 _06407_ (.A0(\reg_module.gprf[873] ),
    .A1(\reg_module.gprf[841] ),
    .A2(\reg_module.gprf[809] ),
    .A3(\reg_module.gprf[777] ),
    .S0(net1032),
    .S1(net998),
    .X(_01477_));
 sky130_fd_sc_hd__mux4_1 _06408_ (.A0(\reg_module.gprf[1001] ),
    .A1(\reg_module.gprf[969] ),
    .A2(\reg_module.gprf[937] ),
    .A3(\reg_module.gprf[905] ),
    .S0(net1032),
    .S1(net998),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _06409_ (.A0(_01477_),
    .A1(_01478_),
    .S(net823),
    .X(_01479_));
 sky130_fd_sc_hd__mux4_1 _06410_ (.A0(\reg_module.gprf[745] ),
    .A1(\reg_module.gprf[713] ),
    .A2(\reg_module.gprf[681] ),
    .A3(\reg_module.gprf[649] ),
    .S0(net1032),
    .S1(net998),
    .X(_01480_));
 sky130_fd_sc_hd__mux4_1 _06411_ (.A0(\reg_module.gprf[617] ),
    .A1(\reg_module.gprf[585] ),
    .A2(\reg_module.gprf[553] ),
    .A3(\reg_module.gprf[521] ),
    .S0(net1036),
    .S1(net1002),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _06412_ (.A0(_01480_),
    .A1(_01481_),
    .S(net992),
    .X(_01482_));
 sky130_fd_sc_hd__nand2_1 _06413_ (.A(net984),
    .B(_01482_),
    .Y(_01483_));
 sky130_fd_sc_hd__a21oi_1 _06414_ (.A1(net818),
    .A2(_01479_),
    .B1(net1066),
    .Y(_01484_));
 sky130_fd_sc_hd__a2bb2o_2 _06415_ (.A1_N(net814),
    .A2_N(_01476_),
    .B1(_01483_),
    .B2(_01484_),
    .X(_01485_));
 sky130_fd_sc_hd__nand2_1 _06416_ (.A(\rWrDataWB[9] ),
    .B(net588),
    .Y(_01486_));
 sky130_fd_sc_hd__o21ai_1 _06417_ (.A1(net587),
    .A2(_01485_),
    .B1(_01486_),
    .Y(_01487_));
 sky130_fd_sc_hd__o21a_1 _06418_ (.A1(net622),
    .A2(_01487_),
    .B1(_01469_),
    .X(_01488_));
 sky130_fd_sc_hd__nand2_1 _06419_ (.A(\brancher.imm12_i_s[9] ),
    .B(_01488_),
    .Y(_01489_));
 sky130_fd_sc_hd__or2_1 _06420_ (.A(\brancher.imm12_i_s[9] ),
    .B(_01488_),
    .X(_01490_));
 sky130_fd_sc_hd__nand2_1 _06421_ (.A(_01489_),
    .B(_01490_),
    .Y(_01491_));
 sky130_fd_sc_hd__o21a_1 _06422_ (.A1(_01466_),
    .A2(_01467_),
    .B1(_01464_),
    .X(_01492_));
 sky130_fd_sc_hd__a21o_1 _06423_ (.A1(_01491_),
    .A2(_01492_),
    .B1(net773),
    .X(_01493_));
 sky130_fd_sc_hd__o21ba_1 _06424_ (.A1(_01491_),
    .A2(_01492_),
    .B1_N(_01493_),
    .X(net102));
 sky130_fd_sc_hd__mux4_1 _06425_ (.A0(\reg_module.gprf[362] ),
    .A1(\reg_module.gprf[330] ),
    .A2(\reg_module.gprf[298] ),
    .A3(\reg_module.gprf[266] ),
    .S0(net1032),
    .S1(net998),
    .X(_01494_));
 sky130_fd_sc_hd__mux4_1 _06426_ (.A0(\reg_module.gprf[490] ),
    .A1(\reg_module.gprf[458] ),
    .A2(\reg_module.gprf[426] ),
    .A3(\reg_module.gprf[394] ),
    .S0(net1032),
    .S1(net998),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _06427_ (.A0(_01494_),
    .A1(_01495_),
    .S(net823),
    .X(_01496_));
 sky130_fd_sc_hd__mux4_1 _06428_ (.A0(\reg_module.gprf[106] ),
    .A1(\reg_module.gprf[74] ),
    .A2(\reg_module.gprf[42] ),
    .A3(\reg_module.gprf[10] ),
    .S0(net1032),
    .S1(net998),
    .X(_01497_));
 sky130_fd_sc_hd__mux4_1 _06429_ (.A0(\reg_module.gprf[234] ),
    .A1(\reg_module.gprf[202] ),
    .A2(\reg_module.gprf[170] ),
    .A3(\reg_module.gprf[138] ),
    .S0(net1033),
    .S1(net999),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _06430_ (.A0(_01497_),
    .A1(_01498_),
    .S(net823),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _06431_ (.A0(_01496_),
    .A1(_01499_),
    .S(net984),
    .X(_01500_));
 sky130_fd_sc_hd__mux4_1 _06432_ (.A0(\reg_module.gprf[874] ),
    .A1(\reg_module.gprf[842] ),
    .A2(\reg_module.gprf[810] ),
    .A3(\reg_module.gprf[778] ),
    .S0(net1033),
    .S1(net999),
    .X(_01501_));
 sky130_fd_sc_hd__mux4_1 _06433_ (.A0(\reg_module.gprf[1002] ),
    .A1(\reg_module.gprf[970] ),
    .A2(\reg_module.gprf[938] ),
    .A3(\reg_module.gprf[906] ),
    .S0(net1033),
    .S1(net999),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _06434_ (.A0(_01501_),
    .A1(_01502_),
    .S(net823),
    .X(_01503_));
 sky130_fd_sc_hd__mux4_1 _06435_ (.A0(\reg_module.gprf[746] ),
    .A1(\reg_module.gprf[714] ),
    .A2(\reg_module.gprf[682] ),
    .A3(\reg_module.gprf[650] ),
    .S0(net1033),
    .S1(net999),
    .X(_01504_));
 sky130_fd_sc_hd__mux4_1 _06436_ (.A0(\reg_module.gprf[618] ),
    .A1(\reg_module.gprf[586] ),
    .A2(\reg_module.gprf[554] ),
    .A3(\reg_module.gprf[522] ),
    .S0(net1032),
    .S1(net998),
    .X(_01505_));
 sky130_fd_sc_hd__mux2_1 _06437_ (.A0(_01504_),
    .A1(_01505_),
    .S(net992),
    .X(_01506_));
 sky130_fd_sc_hd__nand2_1 _06438_ (.A(net984),
    .B(_01506_),
    .Y(_01507_));
 sky130_fd_sc_hd__a21oi_1 _06439_ (.A1(net818),
    .A2(_01503_),
    .B1(net1066),
    .Y(_01508_));
 sky130_fd_sc_hd__a2bb2o_2 _06440_ (.A1_N(net814),
    .A2_N(_01500_),
    .B1(_01507_),
    .B2(_01508_),
    .X(_01509_));
 sky130_fd_sc_hd__nor2_1 _06441_ (.A(net587),
    .B(_01509_),
    .Y(_01510_));
 sky130_fd_sc_hd__a21o_1 _06442_ (.A1(\rWrDataWB[10] ),
    .A2(net587),
    .B1(net622),
    .X(_01511_));
 sky130_fd_sc_hd__o22a_1 _06443_ (.A1(\rWrData[10] ),
    .A2(net616),
    .B1(_01510_),
    .B2(_01511_),
    .X(_01512_));
 sky130_fd_sc_hd__nand2_1 _06444_ (.A(\brancher.imm12_i_s[10] ),
    .B(_01512_),
    .Y(_01513_));
 sky130_fd_sc_hd__xnor2_1 _06445_ (.A(\brancher.imm12_i_s[10] ),
    .B(_01512_),
    .Y(_01514_));
 sky130_fd_sc_hd__o21a_1 _06446_ (.A1(_01491_),
    .A2(_01492_),
    .B1(_01489_),
    .X(_01515_));
 sky130_fd_sc_hd__a21o_1 _06447_ (.A1(_01514_),
    .A2(_01515_),
    .B1(net773),
    .X(_01516_));
 sky130_fd_sc_hd__o21ba_1 _06448_ (.A1(_01514_),
    .A2(_01515_),
    .B1_N(_01516_),
    .X(net72));
 sky130_fd_sc_hd__o21a_1 _06449_ (.A1(_01514_),
    .A2(_01515_),
    .B1(_01513_),
    .X(_01517_));
 sky130_fd_sc_hd__or2_1 _06450_ (.A(\rWrData[11] ),
    .B(net618),
    .X(_01518_));
 sky130_fd_sc_hd__mux4_1 _06451_ (.A0(\reg_module.gprf[363] ),
    .A1(\reg_module.gprf[331] ),
    .A2(\reg_module.gprf[299] ),
    .A3(\reg_module.gprf[267] ),
    .S0(net1038),
    .S1(net1004),
    .X(_01519_));
 sky130_fd_sc_hd__mux4_1 _06452_ (.A0(\reg_module.gprf[491] ),
    .A1(\reg_module.gprf[459] ),
    .A2(\reg_module.gprf[427] ),
    .A3(\reg_module.gprf[395] ),
    .S0(net1038),
    .S1(net1004),
    .X(_01520_));
 sky130_fd_sc_hd__mux2_1 _06453_ (.A0(_01519_),
    .A1(_01520_),
    .S(net825),
    .X(_01521_));
 sky130_fd_sc_hd__mux4_1 _06454_ (.A0(\reg_module.gprf[107] ),
    .A1(\reg_module.gprf[75] ),
    .A2(\reg_module.gprf[43] ),
    .A3(\reg_module.gprf[11] ),
    .S0(net1038),
    .S1(net1004),
    .X(_01522_));
 sky130_fd_sc_hd__mux4_1 _06455_ (.A0(\reg_module.gprf[235] ),
    .A1(\reg_module.gprf[203] ),
    .A2(\reg_module.gprf[171] ),
    .A3(\reg_module.gprf[139] ),
    .S0(net1038),
    .S1(net1004),
    .X(_01523_));
 sky130_fd_sc_hd__mux2_1 _06456_ (.A0(_01522_),
    .A1(_01523_),
    .S(net825),
    .X(_01524_));
 sky130_fd_sc_hd__mux2_1 _06457_ (.A0(_01521_),
    .A1(_01524_),
    .S(net985),
    .X(_01525_));
 sky130_fd_sc_hd__mux4_1 _06458_ (.A0(\reg_module.gprf[619] ),
    .A1(\reg_module.gprf[587] ),
    .A2(\reg_module.gprf[555] ),
    .A3(\reg_module.gprf[523] ),
    .S0(net1037),
    .S1(net1003),
    .X(_01526_));
 sky130_fd_sc_hd__mux4_1 _06459_ (.A0(\reg_module.gprf[747] ),
    .A1(\reg_module.gprf[715] ),
    .A2(\reg_module.gprf[683] ),
    .A3(\reg_module.gprf[651] ),
    .S0(net1037),
    .S1(net1003),
    .X(_01527_));
 sky130_fd_sc_hd__or2_1 _06460_ (.A(net993),
    .B(_01527_),
    .X(_01528_));
 sky130_fd_sc_hd__o21a_1 _06461_ (.A1(net825),
    .A2(_01526_),
    .B1(net985),
    .X(_01529_));
 sky130_fd_sc_hd__mux4_1 _06462_ (.A0(\reg_module.gprf[875] ),
    .A1(\reg_module.gprf[843] ),
    .A2(\reg_module.gprf[811] ),
    .A3(\reg_module.gprf[779] ),
    .S0(net1037),
    .S1(net1003),
    .X(_01530_));
 sky130_fd_sc_hd__mux4_1 _06463_ (.A0(\reg_module.gprf[1003] ),
    .A1(\reg_module.gprf[971] ),
    .A2(\reg_module.gprf[939] ),
    .A3(\reg_module.gprf[907] ),
    .S0(net1037),
    .S1(net1003),
    .X(_01531_));
 sky130_fd_sc_hd__mux2_1 _06464_ (.A0(_01530_),
    .A1(_01531_),
    .S(net825),
    .X(_01532_));
 sky130_fd_sc_hd__a221o_1 _06465_ (.A1(_01528_),
    .A2(_01529_),
    .B1(_01532_),
    .B2(net819),
    .C1(net1066),
    .X(_01533_));
 sky130_fd_sc_hd__o21a_2 _06466_ (.A1(net814),
    .A2(_01525_),
    .B1(_01533_),
    .X(_01534_));
 sky130_fd_sc_hd__nand2_1 _06467_ (.A(net596),
    .B(_01534_),
    .Y(_01535_));
 sky130_fd_sc_hd__a21oi_1 _06468_ (.A1(\rWrDataWB[11] ),
    .A2(net588),
    .B1(net623),
    .Y(_01536_));
 sky130_fd_sc_hd__a21bo_1 _06469_ (.A1(_01535_),
    .A2(_01536_),
    .B1_N(_01518_),
    .X(_01537_));
 sky130_fd_sc_hd__and2_1 _06470_ (.A(net812),
    .B(_01537_),
    .X(_01538_));
 sky130_fd_sc_hd__or2_1 _06471_ (.A(net812),
    .B(_01537_),
    .X(_01539_));
 sky130_fd_sc_hd__nand2b_1 _06472_ (.A_N(_01538_),
    .B(_01539_),
    .Y(_01540_));
 sky130_fd_sc_hd__a21oi_1 _06473_ (.A1(_01517_),
    .A2(_01540_),
    .B1(net773),
    .Y(_01541_));
 sky130_fd_sc_hd__o21a_1 _06474_ (.A1(_01517_),
    .A2(_01540_),
    .B1(_01541_),
    .X(net73));
 sky130_fd_sc_hd__or2_1 _06475_ (.A(\rWrData[12] ),
    .B(net618),
    .X(_01542_));
 sky130_fd_sc_hd__mux4_1 _06476_ (.A0(\reg_module.gprf[236] ),
    .A1(\reg_module.gprf[204] ),
    .A2(\reg_module.gprf[172] ),
    .A3(\reg_module.gprf[140] ),
    .S0(net1038),
    .S1(net1005),
    .X(_01543_));
 sky130_fd_sc_hd__mux4_1 _06477_ (.A0(\reg_module.gprf[108] ),
    .A1(\reg_module.gprf[76] ),
    .A2(\reg_module.gprf[44] ),
    .A3(\reg_module.gprf[12] ),
    .S0(net1039),
    .S1(net1005),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _06478_ (.A0(_01543_),
    .A1(_01544_),
    .S(net993),
    .X(_01545_));
 sky130_fd_sc_hd__mux4_1 _06479_ (.A0(\reg_module.gprf[364] ),
    .A1(\reg_module.gprf[332] ),
    .A2(\reg_module.gprf[300] ),
    .A3(\reg_module.gprf[268] ),
    .S0(net1038),
    .S1(net1004),
    .X(_01546_));
 sky130_fd_sc_hd__mux4_1 _06480_ (.A0(\reg_module.gprf[492] ),
    .A1(\reg_module.gprf[460] ),
    .A2(\reg_module.gprf[428] ),
    .A3(\reg_module.gprf[396] ),
    .S0(net1040),
    .S1(net1006),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_1 _06481_ (.A0(_01546_),
    .A1(_01547_),
    .S(net825),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _06482_ (.A0(_01545_),
    .A1(_01548_),
    .S(net819),
    .X(_01549_));
 sky130_fd_sc_hd__mux4_1 _06483_ (.A0(\reg_module.gprf[876] ),
    .A1(\reg_module.gprf[844] ),
    .A2(\reg_module.gprf[812] ),
    .A3(\reg_module.gprf[780] ),
    .S0(net1050),
    .S1(net1016),
    .X(_01550_));
 sky130_fd_sc_hd__mux4_1 _06484_ (.A0(\reg_module.gprf[1004] ),
    .A1(\reg_module.gprf[972] ),
    .A2(\reg_module.gprf[940] ),
    .A3(\reg_module.gprf[908] ),
    .S0(net1052),
    .S1(net1018),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _06485_ (.A0(_01550_),
    .A1(_01551_),
    .S(net829),
    .X(_01552_));
 sky130_fd_sc_hd__mux4_1 _06486_ (.A0(\reg_module.gprf[748] ),
    .A1(\reg_module.gprf[716] ),
    .A2(\reg_module.gprf[684] ),
    .A3(\reg_module.gprf[652] ),
    .S0(net1038),
    .S1(net1004),
    .X(_01553_));
 sky130_fd_sc_hd__mux4_1 _06487_ (.A0(\reg_module.gprf[620] ),
    .A1(\reg_module.gprf[588] ),
    .A2(\reg_module.gprf[556] ),
    .A3(\reg_module.gprf[524] ),
    .S0(net1039),
    .S1(net1004),
    .X(_01554_));
 sky130_fd_sc_hd__or2_1 _06488_ (.A(net825),
    .B(_01554_),
    .X(_01555_));
 sky130_fd_sc_hd__o211a_1 _06489_ (.A1(net994),
    .A2(_01553_),
    .B1(_01555_),
    .C1(net987),
    .X(_01556_));
 sky130_fd_sc_hd__a21o_1 _06490_ (.A1(net819),
    .A2(_01552_),
    .B1(net1067),
    .X(_01557_));
 sky130_fd_sc_hd__o22a_2 _06491_ (.A1(net814),
    .A2(_01549_),
    .B1(_01556_),
    .B2(_01557_),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _06492_ (.A0(\rWrDataWB[12] ),
    .A1(_01558_),
    .S(net596),
    .X(_01559_));
 sky130_fd_sc_hd__o21ai_2 _06493_ (.A1(net623),
    .A2(_01559_),
    .B1(_01542_),
    .Y(_01560_));
 sky130_fd_sc_hd__o211a_1 _06494_ (.A1(_01514_),
    .A2(_01515_),
    .B1(_01539_),
    .C1(_01513_),
    .X(_01561_));
 sky130_fd_sc_hd__o21ai_1 _06495_ (.A1(_01538_),
    .A2(_01561_),
    .B1(_01560_),
    .Y(_01562_));
 sky130_fd_sc_hd__or3_1 _06496_ (.A(_01538_),
    .B(_01560_),
    .C(_01561_),
    .X(_01563_));
 sky130_fd_sc_hd__and3_1 _06497_ (.A(net772),
    .B(_01562_),
    .C(_01563_),
    .X(net74));
 sky130_fd_sc_hd__or2_1 _06498_ (.A(\rWrData[13] ),
    .B(net618),
    .X(_01564_));
 sky130_fd_sc_hd__mux4_1 _06499_ (.A0(\reg_module.gprf[365] ),
    .A1(\reg_module.gprf[333] ),
    .A2(\reg_module.gprf[301] ),
    .A3(\reg_module.gprf[269] ),
    .S0(net1041),
    .S1(net1007),
    .X(_01565_));
 sky130_fd_sc_hd__mux4_1 _06500_ (.A0(\reg_module.gprf[493] ),
    .A1(\reg_module.gprf[461] ),
    .A2(\reg_module.gprf[429] ),
    .A3(\reg_module.gprf[397] ),
    .S0(net1037),
    .S1(net1003),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _06501_ (.A0(_01565_),
    .A1(_01566_),
    .S(net823),
    .X(_01567_));
 sky130_fd_sc_hd__mux4_1 _06502_ (.A0(\reg_module.gprf[109] ),
    .A1(\reg_module.gprf[77] ),
    .A2(\reg_module.gprf[45] ),
    .A3(\reg_module.gprf[13] ),
    .S0(net1037),
    .S1(net1003),
    .X(_01568_));
 sky130_fd_sc_hd__mux4_1 _06503_ (.A0(\reg_module.gprf[237] ),
    .A1(\reg_module.gprf[205] ),
    .A2(\reg_module.gprf[173] ),
    .A3(\reg_module.gprf[141] ),
    .S0(net1037),
    .S1(net1003),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _06504_ (.A0(_01568_),
    .A1(_01569_),
    .S(net825),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _06505_ (.A0(_01567_),
    .A1(_01570_),
    .S(net985),
    .X(_01571_));
 sky130_fd_sc_hd__mux4_1 _06506_ (.A0(\reg_module.gprf[877] ),
    .A1(\reg_module.gprf[845] ),
    .A2(\reg_module.gprf[813] ),
    .A3(\reg_module.gprf[781] ),
    .S0(net1036),
    .S1(net1002),
    .X(_01572_));
 sky130_fd_sc_hd__mux4_1 _06507_ (.A0(\reg_module.gprf[1005] ),
    .A1(\reg_module.gprf[973] ),
    .A2(\reg_module.gprf[941] ),
    .A3(\reg_module.gprf[909] ),
    .S0(net1032),
    .S1(net998),
    .X(_01573_));
 sky130_fd_sc_hd__or2_1 _06508_ (.A(net992),
    .B(_01573_),
    .X(_01574_));
 sky130_fd_sc_hd__o211a_1 _06509_ (.A1(net823),
    .A2(_01572_),
    .B1(_01574_),
    .C1(net818),
    .X(_01575_));
 sky130_fd_sc_hd__mux4_1 _06510_ (.A0(\reg_module.gprf[749] ),
    .A1(\reg_module.gprf[717] ),
    .A2(\reg_module.gprf[685] ),
    .A3(\reg_module.gprf[653] ),
    .S0(net1039),
    .S1(net1005),
    .X(_01576_));
 sky130_fd_sc_hd__mux4_1 _06511_ (.A0(\reg_module.gprf[621] ),
    .A1(\reg_module.gprf[589] ),
    .A2(\reg_module.gprf[557] ),
    .A3(\reg_module.gprf[525] ),
    .S0(net1041),
    .S1(net1007),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _06512_ (.A0(_01576_),
    .A1(_01577_),
    .S(net994),
    .X(_01578_));
 sky130_fd_sc_hd__a21o_1 _06513_ (.A1(net985),
    .A2(_01578_),
    .B1(net1067),
    .X(_01579_));
 sky130_fd_sc_hd__o22a_2 _06514_ (.A1(net814),
    .A2(_01571_),
    .B1(_01575_),
    .B2(_01579_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _06515_ (.A0(\rWrDataWB[13] ),
    .A1(_01580_),
    .S(net596),
    .X(_01581_));
 sky130_fd_sc_hd__o21ai_1 _06516_ (.A1(net622),
    .A2(_01581_),
    .B1(_01564_),
    .Y(_01582_));
 sky130_fd_sc_hd__nand2_1 _06517_ (.A(_01563_),
    .B(_01582_),
    .Y(_01583_));
 sky130_fd_sc_hd__or4_4 _06518_ (.A(_01538_),
    .B(_01560_),
    .C(_01561_),
    .D(_01582_),
    .X(_01584_));
 sky130_fd_sc_hd__and3_1 _06519_ (.A(net772),
    .B(_01583_),
    .C(_01584_),
    .X(net75));
 sky130_fd_sc_hd__or2_1 _06520_ (.A(\rWrData[14] ),
    .B(net618),
    .X(_01585_));
 sky130_fd_sc_hd__mux4_1 _06521_ (.A0(\reg_module.gprf[238] ),
    .A1(\reg_module.gprf[206] ),
    .A2(\reg_module.gprf[174] ),
    .A3(\reg_module.gprf[142] ),
    .S0(net1041),
    .S1(net1007),
    .X(_01586_));
 sky130_fd_sc_hd__mux4_1 _06522_ (.A0(\reg_module.gprf[110] ),
    .A1(\reg_module.gprf[78] ),
    .A2(\reg_module.gprf[46] ),
    .A3(\reg_module.gprf[14] ),
    .S0(net1042),
    .S1(net1008),
    .X(_01587_));
 sky130_fd_sc_hd__or2_1 _06523_ (.A(net826),
    .B(_01587_),
    .X(_01588_));
 sky130_fd_sc_hd__o21a_1 _06524_ (.A1(net993),
    .A2(_01586_),
    .B1(net987),
    .X(_01589_));
 sky130_fd_sc_hd__mux4_1 _06525_ (.A0(\reg_module.gprf[366] ),
    .A1(\reg_module.gprf[334] ),
    .A2(\reg_module.gprf[302] ),
    .A3(\reg_module.gprf[270] ),
    .S0(net1052),
    .S1(net1018),
    .X(_01590_));
 sky130_fd_sc_hd__mux4_1 _06526_ (.A0(\reg_module.gprf[494] ),
    .A1(\reg_module.gprf[462] ),
    .A2(\reg_module.gprf[430] ),
    .A3(\reg_module.gprf[398] ),
    .S0(net1064),
    .S1(net1030),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _06527_ (.A0(_01590_),
    .A1(_01591_),
    .S(net826),
    .X(_01592_));
 sky130_fd_sc_hd__a221o_1 _06528_ (.A1(_01588_),
    .A2(_01589_),
    .B1(_01592_),
    .B2(net819),
    .C1(net814),
    .X(_01593_));
 sky130_fd_sc_hd__mux4_1 _06529_ (.A0(\reg_module.gprf[878] ),
    .A1(\reg_module.gprf[846] ),
    .A2(\reg_module.gprf[814] ),
    .A3(\reg_module.gprf[782] ),
    .S0(net1040),
    .S1(net1006),
    .X(_01594_));
 sky130_fd_sc_hd__or2_1 _06530_ (.A(net826),
    .B(_01594_),
    .X(_01595_));
 sky130_fd_sc_hd__mux4_1 _06531_ (.A0(\reg_module.gprf[1006] ),
    .A1(\reg_module.gprf[974] ),
    .A2(\reg_module.gprf[942] ),
    .A3(\reg_module.gprf[910] ),
    .S0(net1040),
    .S1(net1006),
    .X(_01596_));
 sky130_fd_sc_hd__o211a_1 _06532_ (.A1(net993),
    .A2(_01596_),
    .B1(_01595_),
    .C1(net819),
    .X(_01597_));
 sky130_fd_sc_hd__mux4_1 _06533_ (.A0(\reg_module.gprf[750] ),
    .A1(\reg_module.gprf[718] ),
    .A2(\reg_module.gprf[686] ),
    .A3(\reg_module.gprf[654] ),
    .S0(net1040),
    .S1(net1006),
    .X(_01598_));
 sky130_fd_sc_hd__mux4_1 _06534_ (.A0(\reg_module.gprf[622] ),
    .A1(\reg_module.gprf[590] ),
    .A2(\reg_module.gprf[558] ),
    .A3(\reg_module.gprf[526] ),
    .S0(net1042),
    .S1(net1008),
    .X(_01599_));
 sky130_fd_sc_hd__or2_1 _06535_ (.A(net826),
    .B(_01599_),
    .X(_01600_));
 sky130_fd_sc_hd__o211a_1 _06536_ (.A1(net993),
    .A2(_01598_),
    .B1(_01600_),
    .C1(net985),
    .X(_01601_));
 sky130_fd_sc_hd__o31a_1 _06537_ (.A1(net1067),
    .A2(_01597_),
    .A3(_01601_),
    .B1(_01593_),
    .X(_01602_));
 sky130_fd_sc_hd__o311ai_4 _06538_ (.A1(net1067),
    .A2(_01597_),
    .A3(_01601_),
    .B1(net596),
    .C1(_01593_),
    .Y(_01603_));
 sky130_fd_sc_hd__a21oi_1 _06539_ (.A1(\rWrDataWB[14] ),
    .A2(net588),
    .B1(net623),
    .Y(_01604_));
 sky130_fd_sc_hd__a21bo_2 _06540_ (.A1(_01603_),
    .A2(_01604_),
    .B1_N(_01585_),
    .X(_01605_));
 sky130_fd_sc_hd__nor2_1 _06541_ (.A(_01584_),
    .B(_01605_),
    .Y(_01606_));
 sky130_fd_sc_hd__or2_1 _06542_ (.A(net773),
    .B(_01606_),
    .X(_01607_));
 sky130_fd_sc_hd__a21oi_1 _06543_ (.A1(_01584_),
    .A2(_01605_),
    .B1(_01607_),
    .Y(net76));
 sky130_fd_sc_hd__or2_1 _06544_ (.A(\rWrData[15] ),
    .B(net621),
    .X(_01608_));
 sky130_fd_sc_hd__mux4_1 _06545_ (.A0(\reg_module.gprf[367] ),
    .A1(\reg_module.gprf[335] ),
    .A2(\reg_module.gprf[303] ),
    .A3(\reg_module.gprf[271] ),
    .S0(net1051),
    .S1(net1017),
    .X(_01609_));
 sky130_fd_sc_hd__mux4_1 _06546_ (.A0(\reg_module.gprf[495] ),
    .A1(\reg_module.gprf[463] ),
    .A2(\reg_module.gprf[431] ),
    .A3(\reg_module.gprf[399] ),
    .S0(net1051),
    .S1(net1017),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _06547_ (.A0(_01609_),
    .A1(_01610_),
    .S(net830),
    .X(_01611_));
 sky130_fd_sc_hd__mux4_1 _06548_ (.A0(\reg_module.gprf[111] ),
    .A1(\reg_module.gprf[79] ),
    .A2(\reg_module.gprf[47] ),
    .A3(\reg_module.gprf[15] ),
    .S0(net1052),
    .S1(net1018),
    .X(_01612_));
 sky130_fd_sc_hd__mux4_1 _06549_ (.A0(\reg_module.gprf[239] ),
    .A1(\reg_module.gprf[207] ),
    .A2(\reg_module.gprf[175] ),
    .A3(\reg_module.gprf[143] ),
    .S0(net1052),
    .S1(net1018),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _06550_ (.A0(_01612_),
    .A1(_01613_),
    .S(net830),
    .X(_01614_));
 sky130_fd_sc_hd__mux2_1 _06551_ (.A0(_01611_),
    .A1(_01614_),
    .S(net989),
    .X(_01615_));
 sky130_fd_sc_hd__mux4_1 _06552_ (.A0(\reg_module.gprf[879] ),
    .A1(\reg_module.gprf[847] ),
    .A2(\reg_module.gprf[815] ),
    .A3(\reg_module.gprf[783] ),
    .S0(net1052),
    .S1(net1018),
    .X(_01616_));
 sky130_fd_sc_hd__mux4_1 _06553_ (.A0(\reg_module.gprf[1007] ),
    .A1(\reg_module.gprf[975] ),
    .A2(\reg_module.gprf[943] ),
    .A3(\reg_module.gprf[911] ),
    .S0(net1052),
    .S1(net1018),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _06554_ (.A0(_01616_),
    .A1(_01617_),
    .S(net830),
    .X(_01618_));
 sky130_fd_sc_hd__mux4_1 _06555_ (.A0(\reg_module.gprf[751] ),
    .A1(\reg_module.gprf[719] ),
    .A2(\reg_module.gprf[687] ),
    .A3(\reg_module.gprf[655] ),
    .S0(net1052),
    .S1(net1018),
    .X(_01619_));
 sky130_fd_sc_hd__mux4_1 _06556_ (.A0(\reg_module.gprf[623] ),
    .A1(\reg_module.gprf[591] ),
    .A2(\reg_module.gprf[559] ),
    .A3(\reg_module.gprf[527] ),
    .S0(net1052),
    .S1(net1018),
    .X(_01620_));
 sky130_fd_sc_hd__or2_1 _06557_ (.A(net830),
    .B(_01620_),
    .X(_01621_));
 sky130_fd_sc_hd__o211a_1 _06558_ (.A1(net995),
    .A2(_01619_),
    .B1(_01621_),
    .C1(net989),
    .X(_01622_));
 sky130_fd_sc_hd__a21o_1 _06559_ (.A1(net821),
    .A2(_01618_),
    .B1(net1068),
    .X(_01623_));
 sky130_fd_sc_hd__o22a_2 _06560_ (.A1(net816),
    .A2(_01615_),
    .B1(_01622_),
    .B2(_01623_),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_1 _06561_ (.A0(\rWrDataWB[15] ),
    .A1(_01624_),
    .S(net599),
    .X(_01625_));
 sky130_fd_sc_hd__o21a_1 _06562_ (.A1(net626),
    .A2(_01625_),
    .B1(_01608_),
    .X(_01626_));
 sky130_fd_sc_hd__and2_1 _06563_ (.A(_01606_),
    .B(_01626_),
    .X(_01627_));
 sky130_fd_sc_hd__o21ai_1 _06564_ (.A1(_01606_),
    .A2(_01626_),
    .B1(net772),
    .Y(_01628_));
 sky130_fd_sc_hd__nor2_1 _06565_ (.A(_01627_),
    .B(_01628_),
    .Y(net77));
 sky130_fd_sc_hd__or2_2 _06566_ (.A(\rWrData[16] ),
    .B(net620),
    .X(_01629_));
 sky130_fd_sc_hd__mux4_1 _06567_ (.A0(\reg_module.gprf[368] ),
    .A1(\reg_module.gprf[336] ),
    .A2(\reg_module.gprf[304] ),
    .A3(\reg_module.gprf[272] ),
    .S0(net1063),
    .S1(net1029),
    .X(_01630_));
 sky130_fd_sc_hd__mux4_1 _06568_ (.A0(\reg_module.gprf[496] ),
    .A1(\reg_module.gprf[464] ),
    .A2(\reg_module.gprf[432] ),
    .A3(\reg_module.gprf[400] ),
    .S0(net1063),
    .S1(net1029),
    .X(_01631_));
 sky130_fd_sc_hd__mux4_1 _06569_ (.A0(\reg_module.gprf[112] ),
    .A1(\reg_module.gprf[80] ),
    .A2(\reg_module.gprf[48] ),
    .A3(\reg_module.gprf[16] ),
    .S0(net1063),
    .S1(net1029),
    .X(_01632_));
 sky130_fd_sc_hd__mux4_1 _06570_ (.A0(\reg_module.gprf[240] ),
    .A1(\reg_module.gprf[208] ),
    .A2(\reg_module.gprf[176] ),
    .A3(\reg_module.gprf[144] ),
    .S0(net1063),
    .S1(net1029),
    .X(_01633_));
 sky130_fd_sc_hd__mux4_1 _06571_ (.A0(_01630_),
    .A1(_01631_),
    .A2(_01632_),
    .A3(_01633_),
    .S0(net833),
    .S1(net990),
    .X(_01634_));
 sky130_fd_sc_hd__nor2_1 _06572_ (.A(net817),
    .B(_01634_),
    .Y(_01635_));
 sky130_fd_sc_hd__mux4_1 _06573_ (.A0(\reg_module.gprf[624] ),
    .A1(\reg_module.gprf[592] ),
    .A2(\reg_module.gprf[560] ),
    .A3(\reg_module.gprf[528] ),
    .S0(net1063),
    .S1(net1029),
    .X(_01636_));
 sky130_fd_sc_hd__mux4_1 _06574_ (.A0(\reg_module.gprf[752] ),
    .A1(\reg_module.gprf[720] ),
    .A2(\reg_module.gprf[688] ),
    .A3(\reg_module.gprf[656] ),
    .S0(net1063),
    .S1(net1029),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _06575_ (.A0(_01636_),
    .A1(_01637_),
    .S(net833),
    .X(_01638_));
 sky130_fd_sc_hd__nand2_1 _06576_ (.A(net990),
    .B(_01638_),
    .Y(_01639_));
 sky130_fd_sc_hd__mux4_1 _06577_ (.A0(\reg_module.gprf[880] ),
    .A1(\reg_module.gprf[848] ),
    .A2(\reg_module.gprf[816] ),
    .A3(\reg_module.gprf[784] ),
    .S0(net1063),
    .S1(net1029),
    .X(_01640_));
 sky130_fd_sc_hd__mux4_1 _06578_ (.A0(\reg_module.gprf[1008] ),
    .A1(\reg_module.gprf[976] ),
    .A2(\reg_module.gprf[944] ),
    .A3(\reg_module.gprf[912] ),
    .S0(net1063),
    .S1(net1029),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _06579_ (.A0(_01640_),
    .A1(_01641_),
    .S(net833),
    .X(_01642_));
 sky130_fd_sc_hd__a21oi_1 _06580_ (.A1(net822),
    .A2(_01642_),
    .B1(net1069),
    .Y(_01643_));
 sky130_fd_sc_hd__a21oi_2 _06581_ (.A1(_01639_),
    .A2(_01643_),
    .B1(_01635_),
    .Y(_01644_));
 sky130_fd_sc_hd__a211o_1 _06582_ (.A1(_01639_),
    .A2(_01643_),
    .B1(net594),
    .C1(_01635_),
    .X(_01645_));
 sky130_fd_sc_hd__a21bo_1 _06583_ (.A1(\rWrDataWB[16] ),
    .A2(net594),
    .B1_N(_01645_),
    .X(_01646_));
 sky130_fd_sc_hd__o21a_2 _06584_ (.A1(net627),
    .A2(_01646_),
    .B1(_01629_),
    .X(_01647_));
 sky130_fd_sc_hd__and4bb_1 _06585_ (.A_N(_01584_),
    .B_N(_01605_),
    .C(_01626_),
    .D(_01647_),
    .X(_01648_));
 sky130_fd_sc_hd__nor2_1 _06586_ (.A(net773),
    .B(_01648_),
    .Y(_01649_));
 sky130_fd_sc_hd__o21a_1 _06587_ (.A1(_01627_),
    .A2(_01647_),
    .B1(_01649_),
    .X(net78));
 sky130_fd_sc_hd__or2_2 _06588_ (.A(\rWrData[17] ),
    .B(net621),
    .X(_01650_));
 sky130_fd_sc_hd__mux4_1 _06589_ (.A0(\reg_module.gprf[369] ),
    .A1(\reg_module.gprf[337] ),
    .A2(\reg_module.gprf[305] ),
    .A3(\reg_module.gprf[273] ),
    .S0(net1048),
    .S1(net1014),
    .X(_01651_));
 sky130_fd_sc_hd__mux4_1 _06590_ (.A0(\reg_module.gprf[497] ),
    .A1(\reg_module.gprf[465] ),
    .A2(\reg_module.gprf[433] ),
    .A3(\reg_module.gprf[401] ),
    .S0(net1048),
    .S1(net1014),
    .X(_01652_));
 sky130_fd_sc_hd__mux2_1 _06591_ (.A0(_01651_),
    .A1(_01652_),
    .S(net829),
    .X(_01653_));
 sky130_fd_sc_hd__mux4_1 _06592_ (.A0(\reg_module.gprf[113] ),
    .A1(\reg_module.gprf[81] ),
    .A2(\reg_module.gprf[49] ),
    .A3(\reg_module.gprf[17] ),
    .S0(net1048),
    .S1(net1014),
    .X(_01654_));
 sky130_fd_sc_hd__mux4_1 _06593_ (.A0(\reg_module.gprf[241] ),
    .A1(\reg_module.gprf[209] ),
    .A2(\reg_module.gprf[177] ),
    .A3(\reg_module.gprf[145] ),
    .S0(net1048),
    .S1(net1014),
    .X(_01655_));
 sky130_fd_sc_hd__mux2_1 _06594_ (.A0(_01654_),
    .A1(_01655_),
    .S(net829),
    .X(_01656_));
 sky130_fd_sc_hd__mux2_1 _06595_ (.A0(_01653_),
    .A1(_01656_),
    .S(net989),
    .X(_01657_));
 sky130_fd_sc_hd__mux4_1 _06596_ (.A0(\reg_module.gprf[881] ),
    .A1(\reg_module.gprf[849] ),
    .A2(\reg_module.gprf[817] ),
    .A3(\reg_module.gprf[785] ),
    .S0(net1049),
    .S1(net1015),
    .X(_01658_));
 sky130_fd_sc_hd__mux4_1 _06597_ (.A0(\reg_module.gprf[1009] ),
    .A1(\reg_module.gprf[977] ),
    .A2(\reg_module.gprf[945] ),
    .A3(\reg_module.gprf[913] ),
    .S0(net1049),
    .S1(net1015),
    .X(_01659_));
 sky130_fd_sc_hd__mux2_1 _06598_ (.A0(_01658_),
    .A1(_01659_),
    .S(net829),
    .X(_01660_));
 sky130_fd_sc_hd__mux4_1 _06599_ (.A0(\reg_module.gprf[753] ),
    .A1(\reg_module.gprf[721] ),
    .A2(\reg_module.gprf[689] ),
    .A3(\reg_module.gprf[657] ),
    .S0(net1049),
    .S1(net1015),
    .X(_01661_));
 sky130_fd_sc_hd__mux4_1 _06600_ (.A0(\reg_module.gprf[625] ),
    .A1(\reg_module.gprf[593] ),
    .A2(\reg_module.gprf[561] ),
    .A3(\reg_module.gprf[529] ),
    .S0(net1049),
    .S1(net1015),
    .X(_01662_));
 sky130_fd_sc_hd__mux2_1 _06601_ (.A0(_01661_),
    .A1(_01662_),
    .S(net995),
    .X(_01663_));
 sky130_fd_sc_hd__nand2_1 _06602_ (.A(net989),
    .B(_01663_),
    .Y(_01664_));
 sky130_fd_sc_hd__a21oi_1 _06603_ (.A1(net821),
    .A2(_01660_),
    .B1(net1068),
    .Y(_01665_));
 sky130_fd_sc_hd__a2bb2o_2 _06604_ (.A1_N(net816),
    .A2_N(_01657_),
    .B1(_01664_),
    .B2(_01665_),
    .X(_01666_));
 sky130_fd_sc_hd__nor2_1 _06605_ (.A(net593),
    .B(_01666_),
    .Y(_01667_));
 sky130_fd_sc_hd__a211o_1 _06606_ (.A1(\rWrDataWB[17] ),
    .A2(net593),
    .B1(_01667_),
    .C1(net626),
    .X(_01668_));
 sky130_fd_sc_hd__nand2_2 _06607_ (.A(_01650_),
    .B(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__inv_2 _06608_ (.A(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__and2_1 _06609_ (.A(_01648_),
    .B(_01670_),
    .X(_01671_));
 sky130_fd_sc_hd__o21ai_1 _06610_ (.A1(_01648_),
    .A2(_01670_),
    .B1(net771),
    .Y(_01672_));
 sky130_fd_sc_hd__nor2_1 _06611_ (.A(_01671_),
    .B(_01672_),
    .Y(net79));
 sky130_fd_sc_hd__or2_1 _06612_ (.A(\rWrData[18] ),
    .B(net621),
    .X(_01673_));
 sky130_fd_sc_hd__mux4_1 _06613_ (.A0(\reg_module.gprf[370] ),
    .A1(\reg_module.gprf[338] ),
    .A2(\reg_module.gprf[306] ),
    .A3(\reg_module.gprf[274] ),
    .S0(net1048),
    .S1(net1014),
    .X(_01674_));
 sky130_fd_sc_hd__mux4_1 _06614_ (.A0(\reg_module.gprf[498] ),
    .A1(\reg_module.gprf[466] ),
    .A2(\reg_module.gprf[434] ),
    .A3(\reg_module.gprf[402] ),
    .S0(net1048),
    .S1(net1014),
    .X(_01675_));
 sky130_fd_sc_hd__mux2_1 _06615_ (.A0(_01674_),
    .A1(_01675_),
    .S(net829),
    .X(_01676_));
 sky130_fd_sc_hd__mux4_1 _06616_ (.A0(\reg_module.gprf[114] ),
    .A1(\reg_module.gprf[82] ),
    .A2(\reg_module.gprf[50] ),
    .A3(\reg_module.gprf[18] ),
    .S0(net1038),
    .S1(net1004),
    .X(_01677_));
 sky130_fd_sc_hd__mux4_1 _06617_ (.A0(\reg_module.gprf[242] ),
    .A1(\reg_module.gprf[210] ),
    .A2(\reg_module.gprf[178] ),
    .A3(\reg_module.gprf[146] ),
    .S0(net1048),
    .S1(net1014),
    .X(_01678_));
 sky130_fd_sc_hd__mux2_1 _06618_ (.A0(_01677_),
    .A1(_01678_),
    .S(net829),
    .X(_01679_));
 sky130_fd_sc_hd__mux2_1 _06619_ (.A0(_01676_),
    .A1(_01679_),
    .S(net989),
    .X(_01680_));
 sky130_fd_sc_hd__mux4_1 _06620_ (.A0(\reg_module.gprf[882] ),
    .A1(\reg_module.gprf[850] ),
    .A2(\reg_module.gprf[818] ),
    .A3(\reg_module.gprf[786] ),
    .S0(net1048),
    .S1(net1014),
    .X(_01681_));
 sky130_fd_sc_hd__mux4_1 _06621_ (.A0(\reg_module.gprf[1010] ),
    .A1(\reg_module.gprf[978] ),
    .A2(\reg_module.gprf[946] ),
    .A3(\reg_module.gprf[914] ),
    .S0(net1038),
    .S1(net1004),
    .X(_01682_));
 sky130_fd_sc_hd__mux2_1 _06622_ (.A0(_01681_),
    .A1(_01682_),
    .S(net825),
    .X(_01683_));
 sky130_fd_sc_hd__mux4_1 _06623_ (.A0(\reg_module.gprf[754] ),
    .A1(\reg_module.gprf[722] ),
    .A2(\reg_module.gprf[690] ),
    .A3(\reg_module.gprf[658] ),
    .S0(net1038),
    .S1(net1004),
    .X(_01684_));
 sky130_fd_sc_hd__mux4_1 _06624_ (.A0(\reg_module.gprf[626] ),
    .A1(\reg_module.gprf[594] ),
    .A2(\reg_module.gprf[562] ),
    .A3(\reg_module.gprf[530] ),
    .S0(net1048),
    .S1(net1014),
    .X(_01685_));
 sky130_fd_sc_hd__or2_1 _06625_ (.A(net825),
    .B(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__o211a_1 _06626_ (.A1(net995),
    .A2(_01684_),
    .B1(_01686_),
    .C1(net989),
    .X(_01687_));
 sky130_fd_sc_hd__a21o_1 _06627_ (.A1(net821),
    .A2(_01683_),
    .B1(net1068),
    .X(_01688_));
 sky130_fd_sc_hd__o22a_2 _06628_ (.A1(net816),
    .A2(_01680_),
    .B1(_01687_),
    .B2(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__mux2_1 _06629_ (.A0(\rWrDataWB[18] ),
    .A1(_01689_),
    .S(net599),
    .X(_01690_));
 sky130_fd_sc_hd__o21a_2 _06630_ (.A1(net626),
    .A2(_01690_),
    .B1(_01673_),
    .X(_01691_));
 sky130_fd_sc_hd__or2_1 _06631_ (.A(_01671_),
    .B(_01691_),
    .X(_01692_));
 sky130_fd_sc_hd__nand2_1 _06632_ (.A(_01671_),
    .B(_01691_),
    .Y(_01693_));
 sky130_fd_sc_hd__and3_1 _06633_ (.A(net771),
    .B(_01692_),
    .C(_01693_),
    .X(net80));
 sky130_fd_sc_hd__nor2_1 _06634_ (.A(\rWrData[19] ),
    .B(net621),
    .Y(_01694_));
 sky130_fd_sc_hd__mux4_1 _06635_ (.A0(\reg_module.gprf[371] ),
    .A1(\reg_module.gprf[339] ),
    .A2(\reg_module.gprf[307] ),
    .A3(\reg_module.gprf[275] ),
    .S0(net1051),
    .S1(net1017),
    .X(_01695_));
 sky130_fd_sc_hd__mux4_1 _06636_ (.A0(\reg_module.gprf[499] ),
    .A1(\reg_module.gprf[467] ),
    .A2(\reg_module.gprf[435] ),
    .A3(\reg_module.gprf[403] ),
    .S0(net1049),
    .S1(net1015),
    .X(_01696_));
 sky130_fd_sc_hd__mux4_1 _06637_ (.A0(\reg_module.gprf[115] ),
    .A1(\reg_module.gprf[83] ),
    .A2(\reg_module.gprf[51] ),
    .A3(\reg_module.gprf[19] ),
    .S0(net1050),
    .S1(net1015),
    .X(_01697_));
 sky130_fd_sc_hd__mux4_1 _06638_ (.A0(\reg_module.gprf[243] ),
    .A1(\reg_module.gprf[211] ),
    .A2(\reg_module.gprf[179] ),
    .A3(\reg_module.gprf[147] ),
    .S0(net1050),
    .S1(net1016),
    .X(_01698_));
 sky130_fd_sc_hd__mux4_1 _06639_ (.A0(_01695_),
    .A1(_01696_),
    .A2(_01697_),
    .A3(_01698_),
    .S0(net829),
    .S1(net989),
    .X(_01699_));
 sky130_fd_sc_hd__nor2_1 _06640_ (.A(net816),
    .B(_01699_),
    .Y(_01700_));
 sky130_fd_sc_hd__mux4_1 _06641_ (.A0(\reg_module.gprf[883] ),
    .A1(\reg_module.gprf[851] ),
    .A2(\reg_module.gprf[819] ),
    .A3(\reg_module.gprf[787] ),
    .S0(net1051),
    .S1(net1017),
    .X(_01701_));
 sky130_fd_sc_hd__mux4_1 _06642_ (.A0(\reg_module.gprf[1011] ),
    .A1(\reg_module.gprf[979] ),
    .A2(\reg_module.gprf[947] ),
    .A3(\reg_module.gprf[915] ),
    .S0(net1051),
    .S1(net1017),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _06643_ (.A0(_01701_),
    .A1(_01702_),
    .S(net829),
    .X(_01703_));
 sky130_fd_sc_hd__mux4_1 _06644_ (.A0(\reg_module.gprf[755] ),
    .A1(\reg_module.gprf[723] ),
    .A2(\reg_module.gprf[691] ),
    .A3(\reg_module.gprf[659] ),
    .S0(net1049),
    .S1(net1016),
    .X(_01704_));
 sky130_fd_sc_hd__mux4_1 _06645_ (.A0(\reg_module.gprf[627] ),
    .A1(\reg_module.gprf[595] ),
    .A2(\reg_module.gprf[563] ),
    .A3(\reg_module.gprf[531] ),
    .S0(net1048),
    .S1(net1014),
    .X(_01705_));
 sky130_fd_sc_hd__mux2_1 _06646_ (.A0(_01704_),
    .A1(_01705_),
    .S(net995),
    .X(_01706_));
 sky130_fd_sc_hd__nand2_1 _06647_ (.A(net989),
    .B(_01706_),
    .Y(_01707_));
 sky130_fd_sc_hd__a21oi_1 _06648_ (.A1(net821),
    .A2(_01703_),
    .B1(net1068),
    .Y(_01708_));
 sky130_fd_sc_hd__a21oi_1 _06649_ (.A1(_01707_),
    .A2(_01708_),
    .B1(_01700_),
    .Y(_01709_));
 sky130_fd_sc_hd__a211o_1 _06650_ (.A1(_01707_),
    .A2(_01708_),
    .B1(net593),
    .C1(_01700_),
    .X(_01710_));
 sky130_fd_sc_hd__a21oi_1 _06651_ (.A1(\rWrDataWB[19] ),
    .A2(net593),
    .B1(net626),
    .Y(_01711_));
 sky130_fd_sc_hd__a21oi_2 _06652_ (.A1(_01710_),
    .A2(_01711_),
    .B1(_01694_),
    .Y(_01712_));
 sky130_fd_sc_hd__a31o_1 _06653_ (.A1(_01648_),
    .A2(_01670_),
    .A3(_01691_),
    .B1(_01712_),
    .X(_01713_));
 sky130_fd_sc_hd__nand4_1 _06654_ (.A(_01648_),
    .B(_01670_),
    .C(_01691_),
    .D(_01712_),
    .Y(_01714_));
 sky130_fd_sc_hd__and3_1 _06655_ (.A(net771),
    .B(_01713_),
    .C(_01714_),
    .X(net81));
 sky130_fd_sc_hd__or2_2 _06656_ (.A(\rWrData[20] ),
    .B(net621),
    .X(_01715_));
 sky130_fd_sc_hd__mux4_1 _06657_ (.A0(\reg_module.gprf[244] ),
    .A1(\reg_module.gprf[212] ),
    .A2(\reg_module.gprf[180] ),
    .A3(\reg_module.gprf[148] ),
    .S0(net1040),
    .S1(net1006),
    .X(_01716_));
 sky130_fd_sc_hd__mux4_1 _06658_ (.A0(\reg_module.gprf[116] ),
    .A1(\reg_module.gprf[84] ),
    .A2(\reg_module.gprf[52] ),
    .A3(\reg_module.gprf[20] ),
    .S0(net1040),
    .S1(net1006),
    .X(_01717_));
 sky130_fd_sc_hd__or2_1 _06659_ (.A(net826),
    .B(_01717_),
    .X(_01718_));
 sky130_fd_sc_hd__o21a_1 _06660_ (.A1(net994),
    .A2(_01716_),
    .B1(net985),
    .X(_01719_));
 sky130_fd_sc_hd__mux4_1 _06661_ (.A0(\reg_module.gprf[372] ),
    .A1(\reg_module.gprf[340] ),
    .A2(\reg_module.gprf[308] ),
    .A3(\reg_module.gprf[276] ),
    .S0(net1040),
    .S1(net1006),
    .X(_01720_));
 sky130_fd_sc_hd__mux4_1 _06662_ (.A0(\reg_module.gprf[500] ),
    .A1(\reg_module.gprf[468] ),
    .A2(\reg_module.gprf[436] ),
    .A3(\reg_module.gprf[404] ),
    .S0(net1052),
    .S1(net1018),
    .X(_01721_));
 sky130_fd_sc_hd__mux2_1 _06663_ (.A0(_01720_),
    .A1(_01721_),
    .S(net826),
    .X(_01722_));
 sky130_fd_sc_hd__a221o_1 _06664_ (.A1(_01718_),
    .A2(_01719_),
    .B1(_01722_),
    .B2(net819),
    .C1(net814),
    .X(_01723_));
 sky130_fd_sc_hd__mux4_1 _06665_ (.A0(\reg_module.gprf[884] ),
    .A1(\reg_module.gprf[852] ),
    .A2(\reg_module.gprf[820] ),
    .A3(\reg_module.gprf[788] ),
    .S0(net1040),
    .S1(net1006),
    .X(_01724_));
 sky130_fd_sc_hd__or2_1 _06666_ (.A(net825),
    .B(_01724_),
    .X(_01725_));
 sky130_fd_sc_hd__mux4_1 _06667_ (.A0(\reg_module.gprf[1012] ),
    .A1(\reg_module.gprf[980] ),
    .A2(\reg_module.gprf[948] ),
    .A3(\reg_module.gprf[916] ),
    .S0(net1040),
    .S1(net1006),
    .X(_01726_));
 sky130_fd_sc_hd__o21a_1 _06668_ (.A1(net995),
    .A2(_01726_),
    .B1(net821),
    .X(_01727_));
 sky130_fd_sc_hd__mux4_1 _06669_ (.A0(\reg_module.gprf[756] ),
    .A1(\reg_module.gprf[724] ),
    .A2(\reg_module.gprf[692] ),
    .A3(\reg_module.gprf[660] ),
    .S0(net1040),
    .S1(net1006),
    .X(_01728_));
 sky130_fd_sc_hd__mux4_1 _06670_ (.A0(\reg_module.gprf[628] ),
    .A1(\reg_module.gprf[596] ),
    .A2(\reg_module.gprf[564] ),
    .A3(\reg_module.gprf[532] ),
    .S0(net1042),
    .S1(net1008),
    .X(_01729_));
 sky130_fd_sc_hd__mux2_1 _06671_ (.A0(_01728_),
    .A1(_01729_),
    .S(net993),
    .X(_01730_));
 sky130_fd_sc_hd__a221o_1 _06672_ (.A1(_01725_),
    .A2(_01727_),
    .B1(_01730_),
    .B2(net985),
    .C1(net1066),
    .X(_01731_));
 sky130_fd_sc_hd__nand2_1 _06673_ (.A(_01723_),
    .B(_01731_),
    .Y(_01732_));
 sky130_fd_sc_hd__and3_1 _06674_ (.A(net599),
    .B(_01723_),
    .C(_01731_),
    .X(_01733_));
 sky130_fd_sc_hd__a211o_1 _06675_ (.A1(\rWrDataWB[20] ),
    .A2(net593),
    .B1(_01733_),
    .C1(net626),
    .X(_01734_));
 sky130_fd_sc_hd__nand2_2 _06676_ (.A(_01715_),
    .B(_01734_),
    .Y(_01735_));
 sky130_fd_sc_hd__nor2_1 _06677_ (.A(_01714_),
    .B(_01735_),
    .Y(_01736_));
 sky130_fd_sc_hd__or2_1 _06678_ (.A(net773),
    .B(_01736_),
    .X(_01737_));
 sky130_fd_sc_hd__a21oi_1 _06679_ (.A1(_01714_),
    .A2(_01735_),
    .B1(_01737_),
    .Y(net83));
 sky130_fd_sc_hd__or2_1 _06680_ (.A(\rWrData[21] ),
    .B(net620),
    .X(_01738_));
 sky130_fd_sc_hd__mux4_1 _06681_ (.A0(\reg_module.gprf[373] ),
    .A1(\reg_module.gprf[341] ),
    .A2(\reg_module.gprf[309] ),
    .A3(\reg_module.gprf[277] ),
    .S0(net1062),
    .S1(net1028),
    .X(_01739_));
 sky130_fd_sc_hd__mux4_1 _06682_ (.A0(\reg_module.gprf[501] ),
    .A1(\reg_module.gprf[469] ),
    .A2(\reg_module.gprf[437] ),
    .A3(\reg_module.gprf[405] ),
    .S0(net1062),
    .S1(net1027),
    .X(_01740_));
 sky130_fd_sc_hd__mux2_1 _06683_ (.A0(_01739_),
    .A1(_01740_),
    .S(net833),
    .X(_01741_));
 sky130_fd_sc_hd__mux4_1 _06684_ (.A0(\reg_module.gprf[117] ),
    .A1(\reg_module.gprf[85] ),
    .A2(\reg_module.gprf[53] ),
    .A3(\reg_module.gprf[21] ),
    .S0(net1062),
    .S1(net1028),
    .X(_01742_));
 sky130_fd_sc_hd__mux4_1 _06685_ (.A0(\reg_module.gprf[245] ),
    .A1(\reg_module.gprf[213] ),
    .A2(\reg_module.gprf[181] ),
    .A3(\reg_module.gprf[149] ),
    .S0(net1061),
    .S1(net1027),
    .X(_01743_));
 sky130_fd_sc_hd__mux2_1 _06686_ (.A0(_01742_),
    .A1(_01743_),
    .S(net834),
    .X(_01744_));
 sky130_fd_sc_hd__mux2_1 _06687_ (.A0(_01741_),
    .A1(_01744_),
    .S(net990),
    .X(_01745_));
 sky130_fd_sc_hd__mux4_1 _06688_ (.A0(\reg_module.gprf[629] ),
    .A1(\reg_module.gprf[597] ),
    .A2(\reg_module.gprf[565] ),
    .A3(\reg_module.gprf[533] ),
    .S0(net1062),
    .S1(net1028),
    .X(_01746_));
 sky130_fd_sc_hd__or2_1 _06689_ (.A(net834),
    .B(_01746_),
    .X(_01747_));
 sky130_fd_sc_hd__mux4_1 _06690_ (.A0(\reg_module.gprf[757] ),
    .A1(\reg_module.gprf[725] ),
    .A2(\reg_module.gprf[693] ),
    .A3(\reg_module.gprf[661] ),
    .S0(net1061),
    .S1(net1027),
    .X(_01748_));
 sky130_fd_sc_hd__o21a_1 _06691_ (.A1(net997),
    .A2(_01748_),
    .B1(net990),
    .X(_01749_));
 sky130_fd_sc_hd__mux4_1 _06692_ (.A0(\reg_module.gprf[885] ),
    .A1(\reg_module.gprf[853] ),
    .A2(\reg_module.gprf[821] ),
    .A3(\reg_module.gprf[789] ),
    .S0(net1061),
    .S1(net1028),
    .X(_01750_));
 sky130_fd_sc_hd__mux4_1 _06693_ (.A0(\reg_module.gprf[1013] ),
    .A1(\reg_module.gprf[981] ),
    .A2(\reg_module.gprf[949] ),
    .A3(\reg_module.gprf[917] ),
    .S0(net1062),
    .S1(net1028),
    .X(_01751_));
 sky130_fd_sc_hd__mux2_1 _06694_ (.A0(_01750_),
    .A1(_01751_),
    .S(net834),
    .X(_01752_));
 sky130_fd_sc_hd__a221o_1 _06695_ (.A1(_01747_),
    .A2(_01749_),
    .B1(_01752_),
    .B2(net822),
    .C1(net1069),
    .X(_01753_));
 sky130_fd_sc_hd__o21a_1 _06696_ (.A1(net817),
    .A2(_01745_),
    .B1(_01753_),
    .X(_01754_));
 sky130_fd_sc_hd__o211ai_1 _06697_ (.A1(net817),
    .A2(_01745_),
    .B1(_01753_),
    .C1(net598),
    .Y(_01755_));
 sky130_fd_sc_hd__a21bo_1 _06698_ (.A1(\rWrDataWB[21] ),
    .A2(net594),
    .B1_N(_01755_),
    .X(_01756_));
 sky130_fd_sc_hd__o21a_2 _06699_ (.A1(net627),
    .A2(_01756_),
    .B1(_01738_),
    .X(_01757_));
 sky130_fd_sc_hd__inv_2 _06700_ (.A(_01757_),
    .Y(_01758_));
 sky130_fd_sc_hd__or2_1 _06701_ (.A(_01736_),
    .B(_01757_),
    .X(_01759_));
 sky130_fd_sc_hd__nand2_1 _06702_ (.A(_01736_),
    .B(_01757_),
    .Y(_01760_));
 sky130_fd_sc_hd__and3_1 _06703_ (.A(net772),
    .B(_01759_),
    .C(_01760_),
    .X(net84));
 sky130_fd_sc_hd__or2_1 _06704_ (.A(\rWrData[22] ),
    .B(net620),
    .X(_01761_));
 sky130_fd_sc_hd__mux4_1 _06705_ (.A0(\reg_module.gprf[374] ),
    .A1(\reg_module.gprf[342] ),
    .A2(\reg_module.gprf[310] ),
    .A3(\reg_module.gprf[278] ),
    .S0(net1060),
    .S1(net1025),
    .X(_01762_));
 sky130_fd_sc_hd__mux4_1 _06706_ (.A0(\reg_module.gprf[502] ),
    .A1(\reg_module.gprf[470] ),
    .A2(\reg_module.gprf[438] ),
    .A3(\reg_module.gprf[406] ),
    .S0(net1060),
    .S1(net1026),
    .X(_01763_));
 sky130_fd_sc_hd__mux4_1 _06707_ (.A0(\reg_module.gprf[118] ),
    .A1(\reg_module.gprf[86] ),
    .A2(\reg_module.gprf[54] ),
    .A3(\reg_module.gprf[22] ),
    .S0(net1060),
    .S1(net1026),
    .X(_01764_));
 sky130_fd_sc_hd__mux4_1 _06708_ (.A0(\reg_module.gprf[246] ),
    .A1(\reg_module.gprf[214] ),
    .A2(\reg_module.gprf[182] ),
    .A3(\reg_module.gprf[150] ),
    .S0(net1059),
    .S1(net1025),
    .X(_01765_));
 sky130_fd_sc_hd__mux4_1 _06709_ (.A0(_01762_),
    .A1(_01763_),
    .A2(_01764_),
    .A3(_01765_),
    .S0(net833),
    .S1(net991),
    .X(_01766_));
 sky130_fd_sc_hd__nor2_1 _06710_ (.A(net817),
    .B(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__mux4_1 _06711_ (.A0(\reg_module.gprf[886] ),
    .A1(\reg_module.gprf[854] ),
    .A2(\reg_module.gprf[822] ),
    .A3(\reg_module.gprf[790] ),
    .S0(net1059),
    .S1(net1025),
    .X(_01768_));
 sky130_fd_sc_hd__mux4_1 _06712_ (.A0(\reg_module.gprf[1014] ),
    .A1(\reg_module.gprf[982] ),
    .A2(\reg_module.gprf[950] ),
    .A3(\reg_module.gprf[918] ),
    .S0(net1059),
    .S1(net1026),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _06713_ (.A0(_01768_),
    .A1(_01769_),
    .S(net833),
    .X(_01770_));
 sky130_fd_sc_hd__nand2_1 _06714_ (.A(net822),
    .B(_01770_),
    .Y(_01771_));
 sky130_fd_sc_hd__mux4_1 _06715_ (.A0(\reg_module.gprf[758] ),
    .A1(\reg_module.gprf[726] ),
    .A2(\reg_module.gprf[694] ),
    .A3(\reg_module.gprf[662] ),
    .S0(net1059),
    .S1(net1025),
    .X(_01772_));
 sky130_fd_sc_hd__mux4_1 _06716_ (.A0(\reg_module.gprf[630] ),
    .A1(\reg_module.gprf[598] ),
    .A2(\reg_module.gprf[566] ),
    .A3(\reg_module.gprf[534] ),
    .S0(net1060),
    .S1(net1026),
    .X(_01773_));
 sky130_fd_sc_hd__mux2_1 _06717_ (.A0(_01772_),
    .A1(_01773_),
    .S(net997),
    .X(_01774_));
 sky130_fd_sc_hd__a21oi_1 _06718_ (.A1(net990),
    .A2(_01774_),
    .B1(net1070),
    .Y(_01775_));
 sky130_fd_sc_hd__a21oi_2 _06719_ (.A1(_01771_),
    .A2(_01775_),
    .B1(_01767_),
    .Y(_01776_));
 sky130_fd_sc_hd__a211o_1 _06720_ (.A1(_01771_),
    .A2(_01775_),
    .B1(net592),
    .C1(_01767_),
    .X(_01777_));
 sky130_fd_sc_hd__a21oi_1 _06721_ (.A1(\rWrDataWB[22] ),
    .A2(net594),
    .B1(net627),
    .Y(_01778_));
 sky130_fd_sc_hd__a21bo_1 _06722_ (.A1(_01777_),
    .A2(_01778_),
    .B1_N(_01761_),
    .X(_01779_));
 sky130_fd_sc_hd__nand2_1 _06723_ (.A(_01760_),
    .B(_01779_),
    .Y(_01780_));
 sky130_fd_sc_hd__or4_1 _06724_ (.A(_01714_),
    .B(_01735_),
    .C(_01758_),
    .D(_01779_),
    .X(_01781_));
 sky130_fd_sc_hd__and3_1 _06725_ (.A(net771),
    .B(_01780_),
    .C(_01781_),
    .X(net85));
 sky130_fd_sc_hd__or2_2 _06726_ (.A(\rWrData[23] ),
    .B(net619),
    .X(_01782_));
 sky130_fd_sc_hd__mux4_1 _06727_ (.A0(\reg_module.gprf[247] ),
    .A1(\reg_module.gprf[215] ),
    .A2(\reg_module.gprf[183] ),
    .A3(\reg_module.gprf[151] ),
    .S0(net1054),
    .S1(net1020),
    .X(_01783_));
 sky130_fd_sc_hd__mux4_1 _06728_ (.A0(\reg_module.gprf[119] ),
    .A1(\reg_module.gprf[87] ),
    .A2(\reg_module.gprf[55] ),
    .A3(\reg_module.gprf[23] ),
    .S0(net1054),
    .S1(net1020),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _06729_ (.A0(_01783_),
    .A1(_01784_),
    .S(net996),
    .X(_01785_));
 sky130_fd_sc_hd__mux4_1 _06730_ (.A0(\reg_module.gprf[375] ),
    .A1(\reg_module.gprf[343] ),
    .A2(\reg_module.gprf[311] ),
    .A3(\reg_module.gprf[279] ),
    .S0(net1053),
    .S1(net1019),
    .X(_01786_));
 sky130_fd_sc_hd__mux4_1 _06731_ (.A0(\reg_module.gprf[503] ),
    .A1(\reg_module.gprf[471] ),
    .A2(\reg_module.gprf[439] ),
    .A3(\reg_module.gprf[407] ),
    .S0(net1054),
    .S1(net1020),
    .X(_01787_));
 sky130_fd_sc_hd__mux2_1 _06732_ (.A0(_01786_),
    .A1(_01787_),
    .S(net831),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _06733_ (.A0(_01785_),
    .A1(_01788_),
    .S(net821),
    .X(_01789_));
 sky130_fd_sc_hd__mux4_1 _06734_ (.A0(\reg_module.gprf[887] ),
    .A1(\reg_module.gprf[855] ),
    .A2(\reg_module.gprf[823] ),
    .A3(\reg_module.gprf[791] ),
    .S0(net1054),
    .S1(net1020),
    .X(_01790_));
 sky130_fd_sc_hd__mux4_1 _06735_ (.A0(\reg_module.gprf[1015] ),
    .A1(\reg_module.gprf[983] ),
    .A2(\reg_module.gprf[951] ),
    .A3(\reg_module.gprf[919] ),
    .S0(net1054),
    .S1(net1020),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _06736_ (.A0(_01790_),
    .A1(_01791_),
    .S(net831),
    .X(_01792_));
 sky130_fd_sc_hd__mux4_1 _06737_ (.A0(\reg_module.gprf[759] ),
    .A1(\reg_module.gprf[727] ),
    .A2(\reg_module.gprf[695] ),
    .A3(\reg_module.gprf[663] ),
    .S0(net1054),
    .S1(net1020),
    .X(_01793_));
 sky130_fd_sc_hd__mux4_1 _06738_ (.A0(\reg_module.gprf[631] ),
    .A1(\reg_module.gprf[599] ),
    .A2(\reg_module.gprf[567] ),
    .A3(\reg_module.gprf[535] ),
    .S0(net1054),
    .S1(net1020),
    .X(_01794_));
 sky130_fd_sc_hd__mux2_1 _06739_ (.A0(_01793_),
    .A1(_01794_),
    .S(net995),
    .X(_01795_));
 sky130_fd_sc_hd__nand2_1 _06740_ (.A(net988),
    .B(_01795_),
    .Y(_01796_));
 sky130_fd_sc_hd__a21oi_1 _06741_ (.A1(net821),
    .A2(_01792_),
    .B1(net1068),
    .Y(_01797_));
 sky130_fd_sc_hd__a2bb2o_2 _06742_ (.A1_N(net816),
    .A2_N(_01789_),
    .B1(_01796_),
    .B2(_01797_),
    .X(_01798_));
 sky130_fd_sc_hd__nor2_1 _06743_ (.A(net591),
    .B(_01798_),
    .Y(_01799_));
 sky130_fd_sc_hd__a211o_1 _06744_ (.A1(\rWrDataWB[23] ),
    .A2(net590),
    .B1(_01799_),
    .C1(net625),
    .X(_01800_));
 sky130_fd_sc_hd__nand2_1 _06745_ (.A(_01782_),
    .B(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__nor2_1 _06746_ (.A(_01781_),
    .B(_01801_),
    .Y(_01802_));
 sky130_fd_sc_hd__a21o_1 _06747_ (.A1(_01781_),
    .A2(_01801_),
    .B1(_01284_),
    .X(_01803_));
 sky130_fd_sc_hd__nor2_1 _06748_ (.A(_01802_),
    .B(_01803_),
    .Y(net86));
 sky130_fd_sc_hd__or2_2 _06749_ (.A(\rWrData[24] ),
    .B(net619),
    .X(_01804_));
 sky130_fd_sc_hd__mux4_1 _06750_ (.A0(\reg_module.gprf[376] ),
    .A1(\reg_module.gprf[344] ),
    .A2(\reg_module.gprf[312] ),
    .A3(\reg_module.gprf[280] ),
    .S0(net1055),
    .S1(net1021),
    .X(_01805_));
 sky130_fd_sc_hd__mux4_1 _06751_ (.A0(\reg_module.gprf[504] ),
    .A1(\reg_module.gprf[472] ),
    .A2(\reg_module.gprf[440] ),
    .A3(\reg_module.gprf[408] ),
    .S0(net1057),
    .S1(net1023),
    .X(_01806_));
 sky130_fd_sc_hd__mux2_1 _06752_ (.A0(_01805_),
    .A1(_01806_),
    .S(net832),
    .X(_01807_));
 sky130_fd_sc_hd__mux4_1 _06753_ (.A0(\reg_module.gprf[120] ),
    .A1(\reg_module.gprf[88] ),
    .A2(\reg_module.gprf[56] ),
    .A3(\reg_module.gprf[24] ),
    .S0(net1057),
    .S1(net1023),
    .X(_01808_));
 sky130_fd_sc_hd__mux4_1 _06754_ (.A0(\reg_module.gprf[248] ),
    .A1(\reg_module.gprf[216] ),
    .A2(\reg_module.gprf[184] ),
    .A3(\reg_module.gprf[152] ),
    .S0(net1055),
    .S1(net1021),
    .X(_01809_));
 sky130_fd_sc_hd__mux2_1 _06755_ (.A0(_01808_),
    .A1(_01809_),
    .S(net832),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _06756_ (.A0(_01807_),
    .A1(_01810_),
    .S(net988),
    .X(_01811_));
 sky130_fd_sc_hd__mux4_1 _06757_ (.A0(\reg_module.gprf[888] ),
    .A1(\reg_module.gprf[856] ),
    .A2(\reg_module.gprf[824] ),
    .A3(\reg_module.gprf[792] ),
    .S0(net1057),
    .S1(net1023),
    .X(_01812_));
 sky130_fd_sc_hd__mux4_1 _06758_ (.A0(\reg_module.gprf[1016] ),
    .A1(\reg_module.gprf[984] ),
    .A2(\reg_module.gprf[952] ),
    .A3(\reg_module.gprf[920] ),
    .S0(net1057),
    .S1(net1023),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _06759_ (.A0(_01812_),
    .A1(_01813_),
    .S(net832),
    .X(_01814_));
 sky130_fd_sc_hd__mux4_1 _06760_ (.A0(\reg_module.gprf[760] ),
    .A1(\reg_module.gprf[728] ),
    .A2(\reg_module.gprf[696] ),
    .A3(\reg_module.gprf[664] ),
    .S0(net1055),
    .S1(net1021),
    .X(_01815_));
 sky130_fd_sc_hd__mux4_1 _06761_ (.A0(\reg_module.gprf[632] ),
    .A1(\reg_module.gprf[600] ),
    .A2(\reg_module.gprf[568] ),
    .A3(\reg_module.gprf[536] ),
    .S0(net1055),
    .S1(net1021),
    .X(_01816_));
 sky130_fd_sc_hd__or2_1 _06762_ (.A(net832),
    .B(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__o211a_1 _06763_ (.A1(net996),
    .A2(_01815_),
    .B1(_01817_),
    .C1(net991),
    .X(_01818_));
 sky130_fd_sc_hd__a21o_1 _06764_ (.A1(net821),
    .A2(_01814_),
    .B1(net1068),
    .X(_01819_));
 sky130_fd_sc_hd__o22a_1 _06765_ (.A1(net816),
    .A2(_01811_),
    .B1(_01818_),
    .B2(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__mux2_1 _06766_ (.A0(\rWrDataWB[24] ),
    .A1(_01820_),
    .S(net598),
    .X(_01821_));
 sky130_fd_sc_hd__o21a_1 _06767_ (.A1(net625),
    .A2(_01821_),
    .B1(_01804_),
    .X(_01822_));
 sky130_fd_sc_hd__inv_2 _06768_ (.A(_01822_),
    .Y(_01823_));
 sky130_fd_sc_hd__or2_1 _06769_ (.A(_01802_),
    .B(_01822_),
    .X(_01824_));
 sky130_fd_sc_hd__nand2_1 _06770_ (.A(_01802_),
    .B(_01822_),
    .Y(_01825_));
 sky130_fd_sc_hd__and3_1 _06771_ (.A(net771),
    .B(_01824_),
    .C(_01825_),
    .X(net87));
 sky130_fd_sc_hd__or2_1 _06772_ (.A(\rWrData[25] ),
    .B(net621),
    .X(_01826_));
 sky130_fd_sc_hd__mux4_1 _06773_ (.A0(\reg_module.gprf[377] ),
    .A1(\reg_module.gprf[345] ),
    .A2(\reg_module.gprf[313] ),
    .A3(\reg_module.gprf[281] ),
    .S0(net1053),
    .S1(net1019),
    .X(_01827_));
 sky130_fd_sc_hd__mux4_1 _06774_ (.A0(\reg_module.gprf[505] ),
    .A1(\reg_module.gprf[473] ),
    .A2(\reg_module.gprf[441] ),
    .A3(\reg_module.gprf[409] ),
    .S0(net1055),
    .S1(net1021),
    .X(_01828_));
 sky130_fd_sc_hd__mux2_1 _06775_ (.A0(_01827_),
    .A1(_01828_),
    .S(net831),
    .X(_01829_));
 sky130_fd_sc_hd__mux4_1 _06776_ (.A0(\reg_module.gprf[121] ),
    .A1(\reg_module.gprf[89] ),
    .A2(\reg_module.gprf[57] ),
    .A3(\reg_module.gprf[25] ),
    .S0(net1058),
    .S1(net1024),
    .X(_01830_));
 sky130_fd_sc_hd__mux4_1 _06777_ (.A0(\reg_module.gprf[249] ),
    .A1(\reg_module.gprf[217] ),
    .A2(\reg_module.gprf[185] ),
    .A3(\reg_module.gprf[153] ),
    .S0(net1055),
    .S1(net1021),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _06778_ (.A0(_01830_),
    .A1(_01831_),
    .S(net831),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _06779_ (.A0(_01829_),
    .A1(_01832_),
    .S(net988),
    .X(_01833_));
 sky130_fd_sc_hd__mux4_1 _06780_ (.A0(\reg_module.gprf[633] ),
    .A1(\reg_module.gprf[601] ),
    .A2(\reg_module.gprf[569] ),
    .A3(\reg_module.gprf[537] ),
    .S0(net1055),
    .S1(net1021),
    .X(_01834_));
 sky130_fd_sc_hd__mux4_1 _06781_ (.A0(\reg_module.gprf[761] ),
    .A1(\reg_module.gprf[729] ),
    .A2(\reg_module.gprf[697] ),
    .A3(\reg_module.gprf[665] ),
    .S0(net1053),
    .S1(net1019),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _06782_ (.A0(_01834_),
    .A1(_01835_),
    .S(net832),
    .X(_01836_));
 sky130_fd_sc_hd__nand2_1 _06783_ (.A(net988),
    .B(_01836_),
    .Y(_01837_));
 sky130_fd_sc_hd__mux4_1 _06784_ (.A0(\reg_module.gprf[889] ),
    .A1(\reg_module.gprf[857] ),
    .A2(\reg_module.gprf[825] ),
    .A3(\reg_module.gprf[793] ),
    .S0(net1053),
    .S1(net1019),
    .X(_01838_));
 sky130_fd_sc_hd__mux4_1 _06785_ (.A0(\reg_module.gprf[1017] ),
    .A1(\reg_module.gprf[985] ),
    .A2(\reg_module.gprf[953] ),
    .A3(\reg_module.gprf[921] ),
    .S0(net1055),
    .S1(net1021),
    .X(_01839_));
 sky130_fd_sc_hd__mux2_1 _06786_ (.A0(_01838_),
    .A1(_01839_),
    .S(net831),
    .X(_01840_));
 sky130_fd_sc_hd__a21oi_1 _06787_ (.A1(net821),
    .A2(_01840_),
    .B1(net1068),
    .Y(_01841_));
 sky130_fd_sc_hd__a2bb2o_2 _06788_ (.A1_N(net816),
    .A2_N(_01833_),
    .B1(_01837_),
    .B2(_01841_),
    .X(_01842_));
 sky130_fd_sc_hd__nor2_1 _06789_ (.A(net590),
    .B(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__a211o_1 _06790_ (.A1(\rWrDataWB[25] ),
    .A2(net592),
    .B1(_01843_),
    .C1(net627),
    .X(_01844_));
 sky130_fd_sc_hd__nand2_1 _06791_ (.A(_01826_),
    .B(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__nand2_1 _06792_ (.A(_01825_),
    .B(_01845_),
    .Y(_01846_));
 sky130_fd_sc_hd__or4_2 _06793_ (.A(_01781_),
    .B(_01801_),
    .C(_01823_),
    .D(_01845_),
    .X(_01847_));
 sky130_fd_sc_hd__and3_1 _06794_ (.A(net771),
    .B(_01846_),
    .C(_01847_),
    .X(net88));
 sky130_fd_sc_hd__or2_2 _06795_ (.A(\rWrData[26] ),
    .B(net620),
    .X(_01848_));
 sky130_fd_sc_hd__mux4_1 _06796_ (.A0(\reg_module.gprf[378] ),
    .A1(\reg_module.gprf[346] ),
    .A2(\reg_module.gprf[314] ),
    .A3(\reg_module.gprf[282] ),
    .S0(net1065),
    .S1(net1031),
    .X(_01849_));
 sky130_fd_sc_hd__mux4_1 _06797_ (.A0(\reg_module.gprf[506] ),
    .A1(\reg_module.gprf[474] ),
    .A2(\reg_module.gprf[442] ),
    .A3(\reg_module.gprf[410] ),
    .S0(net1051),
    .S1(net1017),
    .X(_01850_));
 sky130_fd_sc_hd__mux4_1 _06798_ (.A0(\reg_module.gprf[122] ),
    .A1(\reg_module.gprf[90] ),
    .A2(\reg_module.gprf[58] ),
    .A3(\reg_module.gprf[26] ),
    .S0(net1051),
    .S1(net1017),
    .X(_01851_));
 sky130_fd_sc_hd__mux4_1 _06799_ (.A0(\reg_module.gprf[250] ),
    .A1(\reg_module.gprf[218] ),
    .A2(\reg_module.gprf[186] ),
    .A3(\reg_module.gprf[154] ),
    .S0(net1051),
    .S1(net1017),
    .X(_01852_));
 sky130_fd_sc_hd__mux4_1 _06800_ (.A0(_01849_),
    .A1(_01850_),
    .A2(_01851_),
    .A3(_01852_),
    .S0(net830),
    .S1(net989),
    .X(_01853_));
 sky130_fd_sc_hd__nor2_1 _06801_ (.A(net817),
    .B(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__mux4_1 _06802_ (.A0(\reg_module.gprf[890] ),
    .A1(\reg_module.gprf[858] ),
    .A2(\reg_module.gprf[826] ),
    .A3(\reg_module.gprf[794] ),
    .S0(net1056),
    .S1(net1022),
    .X(_01855_));
 sky130_fd_sc_hd__mux4_1 _06803_ (.A0(\reg_module.gprf[1018] ),
    .A1(\reg_module.gprf[986] ),
    .A2(\reg_module.gprf[954] ),
    .A3(\reg_module.gprf[922] ),
    .S0(net1056),
    .S1(net1022),
    .X(_01856_));
 sky130_fd_sc_hd__mux2_1 _06804_ (.A0(_01855_),
    .A1(_01856_),
    .S(net832),
    .X(_01857_));
 sky130_fd_sc_hd__mux4_1 _06805_ (.A0(\reg_module.gprf[762] ),
    .A1(\reg_module.gprf[730] ),
    .A2(\reg_module.gprf[698] ),
    .A3(\reg_module.gprf[666] ),
    .S0(net1051),
    .S1(net1017),
    .X(_01858_));
 sky130_fd_sc_hd__mux4_1 _06806_ (.A0(\reg_module.gprf[634] ),
    .A1(\reg_module.gprf[602] ),
    .A2(\reg_module.gprf[570] ),
    .A3(\reg_module.gprf[538] ),
    .S0(net1051),
    .S1(net1017),
    .X(_01859_));
 sky130_fd_sc_hd__mux2_1 _06807_ (.A0(_01858_),
    .A1(_01859_),
    .S(net995),
    .X(_01860_));
 sky130_fd_sc_hd__nand2_1 _06808_ (.A(net989),
    .B(_01860_),
    .Y(_01861_));
 sky130_fd_sc_hd__a21oi_1 _06809_ (.A1(net822),
    .A2(_01857_),
    .B1(net1069),
    .Y(_01862_));
 sky130_fd_sc_hd__a21oi_1 _06810_ (.A1(_01861_),
    .A2(_01862_),
    .B1(_01854_),
    .Y(_01863_));
 sky130_fd_sc_hd__a211o_1 _06811_ (.A1(_01861_),
    .A2(_01862_),
    .B1(net590),
    .C1(_01854_),
    .X(_01864_));
 sky130_fd_sc_hd__a21oi_1 _06812_ (.A1(\rWrDataWB[26] ),
    .A2(net590),
    .B1(net625),
    .Y(_01865_));
 sky130_fd_sc_hd__a21bo_2 _06813_ (.A1(_01864_),
    .A2(_01865_),
    .B1_N(_01848_),
    .X(_01866_));
 sky130_fd_sc_hd__o21ai_1 _06814_ (.A1(_01847_),
    .A2(_01866_),
    .B1(net771),
    .Y(_01867_));
 sky130_fd_sc_hd__a21oi_1 _06815_ (.A1(_01847_),
    .A2(_01866_),
    .B1(_01867_),
    .Y(net89));
 sky130_fd_sc_hd__nor2_1 _06816_ (.A(\rWrData[27] ),
    .B(net619),
    .Y(_01868_));
 sky130_fd_sc_hd__mux4_1 _06817_ (.A0(\reg_module.gprf[379] ),
    .A1(\reg_module.gprf[347] ),
    .A2(\reg_module.gprf[315] ),
    .A3(\reg_module.gprf[283] ),
    .S0(net1054),
    .S1(net1020),
    .X(_01869_));
 sky130_fd_sc_hd__mux4_1 _06818_ (.A0(\reg_module.gprf[507] ),
    .A1(\reg_module.gprf[475] ),
    .A2(\reg_module.gprf[443] ),
    .A3(\reg_module.gprf[411] ),
    .S0(net1049),
    .S1(net1015),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _06819_ (.A0(_01869_),
    .A1(_01870_),
    .S(net831),
    .X(_01871_));
 sky130_fd_sc_hd__mux4_1 _06820_ (.A0(\reg_module.gprf[123] ),
    .A1(\reg_module.gprf[91] ),
    .A2(\reg_module.gprf[59] ),
    .A3(\reg_module.gprf[27] ),
    .S0(net1054),
    .S1(net1020),
    .X(_01872_));
 sky130_fd_sc_hd__mux4_1 _06821_ (.A0(\reg_module.gprf[251] ),
    .A1(\reg_module.gprf[219] ),
    .A2(\reg_module.gprf[187] ),
    .A3(\reg_module.gprf[155] ),
    .S0(net1049),
    .S1(net1015),
    .X(_01873_));
 sky130_fd_sc_hd__mux2_1 _06822_ (.A0(_01872_),
    .A1(_01873_),
    .S(net831),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_1 _06823_ (.A0(_01871_),
    .A1(_01874_),
    .S(net988),
    .X(_01875_));
 sky130_fd_sc_hd__mux4_1 _06824_ (.A0(\reg_module.gprf[891] ),
    .A1(\reg_module.gprf[859] ),
    .A2(\reg_module.gprf[827] ),
    .A3(\reg_module.gprf[795] ),
    .S0(net1049),
    .S1(net1015),
    .X(_01876_));
 sky130_fd_sc_hd__mux4_1 _06825_ (.A0(\reg_module.gprf[1019] ),
    .A1(\reg_module.gprf[987] ),
    .A2(\reg_module.gprf[955] ),
    .A3(\reg_module.gprf[923] ),
    .S0(net1049),
    .S1(net1015),
    .X(_01877_));
 sky130_fd_sc_hd__mux2_1 _06826_ (.A0(_01876_),
    .A1(_01877_),
    .S(net829),
    .X(_01878_));
 sky130_fd_sc_hd__mux4_1 _06827_ (.A0(\reg_module.gprf[763] ),
    .A1(\reg_module.gprf[731] ),
    .A2(\reg_module.gprf[699] ),
    .A3(\reg_module.gprf[667] ),
    .S0(net1050),
    .S1(net1016),
    .X(_01879_));
 sky130_fd_sc_hd__mux4_1 _06828_ (.A0(\reg_module.gprf[635] ),
    .A1(\reg_module.gprf[603] ),
    .A2(\reg_module.gprf[571] ),
    .A3(\reg_module.gprf[539] ),
    .S0(net1054),
    .S1(net1020),
    .X(_01880_));
 sky130_fd_sc_hd__or2_1 _06829_ (.A(net829),
    .B(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__o211a_1 _06830_ (.A1(net996),
    .A2(_01879_),
    .B1(_01881_),
    .C1(net988),
    .X(_01882_));
 sky130_fd_sc_hd__a21o_1 _06831_ (.A1(net821),
    .A2(_01878_),
    .B1(net1068),
    .X(_01883_));
 sky130_fd_sc_hd__o22a_2 _06832_ (.A1(net816),
    .A2(_01875_),
    .B1(_01882_),
    .B2(_01883_),
    .X(_01884_));
 sky130_fd_sc_hd__nand2_1 _06833_ (.A(net598),
    .B(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__nand2_1 _06834_ (.A(\rWrDataWB[27] ),
    .B(net590),
    .Y(_01886_));
 sky130_fd_sc_hd__a31o_1 _06835_ (.A1(net619),
    .A2(_01885_),
    .A3(_01886_),
    .B1(_01868_),
    .X(_01887_));
 sky130_fd_sc_hd__o21ai_1 _06836_ (.A1(_01847_),
    .A2(_01866_),
    .B1(_01887_),
    .Y(_01888_));
 sky130_fd_sc_hd__or3_1 _06837_ (.A(_01847_),
    .B(_01866_),
    .C(_01887_),
    .X(_01889_));
 sky130_fd_sc_hd__and3_1 _06838_ (.A(net771),
    .B(_01888_),
    .C(_01889_),
    .X(net90));
 sky130_fd_sc_hd__or2_2 _06839_ (.A(\rWrData[28] ),
    .B(net619),
    .X(_01890_));
 sky130_fd_sc_hd__mux4_1 _06840_ (.A0(\reg_module.gprf[380] ),
    .A1(\reg_module.gprf[348] ),
    .A2(\reg_module.gprf[316] ),
    .A3(\reg_module.gprf[284] ),
    .S0(net1053),
    .S1(net1019),
    .X(_01891_));
 sky130_fd_sc_hd__mux4_1 _06841_ (.A0(\reg_module.gprf[508] ),
    .A1(\reg_module.gprf[476] ),
    .A2(\reg_module.gprf[444] ),
    .A3(\reg_module.gprf[412] ),
    .S0(net1058),
    .S1(net1024),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _06842_ (.A0(_01891_),
    .A1(_01892_),
    .S(net831),
    .X(_01893_));
 sky130_fd_sc_hd__mux4_1 _06843_ (.A0(\reg_module.gprf[124] ),
    .A1(\reg_module.gprf[92] ),
    .A2(\reg_module.gprf[60] ),
    .A3(\reg_module.gprf[28] ),
    .S0(net1053),
    .S1(net1019),
    .X(_01894_));
 sky130_fd_sc_hd__mux4_1 _06844_ (.A0(\reg_module.gprf[252] ),
    .A1(\reg_module.gprf[220] ),
    .A2(\reg_module.gprf[188] ),
    .A3(\reg_module.gprf[156] ),
    .S0(net1053),
    .S1(net1019),
    .X(_01895_));
 sky130_fd_sc_hd__mux2_1 _06845_ (.A0(_01894_),
    .A1(_01895_),
    .S(net831),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_1 _06846_ (.A0(_01893_),
    .A1(_01896_),
    .S(net988),
    .X(_01897_));
 sky130_fd_sc_hd__mux4_1 _06847_ (.A0(\reg_module.gprf[892] ),
    .A1(\reg_module.gprf[860] ),
    .A2(\reg_module.gprf[828] ),
    .A3(\reg_module.gprf[796] ),
    .S0(net1053),
    .S1(net1019),
    .X(_01898_));
 sky130_fd_sc_hd__mux4_1 _06848_ (.A0(\reg_module.gprf[1020] ),
    .A1(\reg_module.gprf[988] ),
    .A2(\reg_module.gprf[956] ),
    .A3(\reg_module.gprf[924] ),
    .S0(net1053),
    .S1(net1019),
    .X(_01899_));
 sky130_fd_sc_hd__mux2_1 _06849_ (.A0(_01898_),
    .A1(_01899_),
    .S(net831),
    .X(_01900_));
 sky130_fd_sc_hd__mux4_1 _06850_ (.A0(\reg_module.gprf[764] ),
    .A1(\reg_module.gprf[732] ),
    .A2(\reg_module.gprf[700] ),
    .A3(\reg_module.gprf[668] ),
    .S0(net1053),
    .S1(net1019),
    .X(_01901_));
 sky130_fd_sc_hd__mux4_1 _06851_ (.A0(\reg_module.gprf[636] ),
    .A1(\reg_module.gprf[604] ),
    .A2(\reg_module.gprf[572] ),
    .A3(\reg_module.gprf[540] ),
    .S0(net1058),
    .S1(net1024),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_1 _06852_ (.A0(_01901_),
    .A1(_01902_),
    .S(net996),
    .X(_01903_));
 sky130_fd_sc_hd__nand2_1 _06853_ (.A(net988),
    .B(_01903_),
    .Y(_01904_));
 sky130_fd_sc_hd__a21oi_1 _06854_ (.A1(net822),
    .A2(_01900_),
    .B1(net1068),
    .Y(_01905_));
 sky130_fd_sc_hd__a2bb2o_2 _06855_ (.A1_N(net816),
    .A2_N(_01897_),
    .B1(_01904_),
    .B2(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__nor2_1 _06856_ (.A(net591),
    .B(_01906_),
    .Y(_01907_));
 sky130_fd_sc_hd__a211o_1 _06857_ (.A1(\rWrDataWB[28] ),
    .A2(net591),
    .B1(_01907_),
    .C1(net625),
    .X(_01908_));
 sky130_fd_sc_hd__nand2_1 _06858_ (.A(_01890_),
    .B(_01908_),
    .Y(_01909_));
 sky130_fd_sc_hd__nand2_1 _06859_ (.A(_01889_),
    .B(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hd__or2_1 _06860_ (.A(_01889_),
    .B(_01909_),
    .X(_01911_));
 sky130_fd_sc_hd__and3_1 _06861_ (.A(net771),
    .B(_01910_),
    .C(_01911_),
    .X(net91));
 sky130_fd_sc_hd__nor2_1 _06862_ (.A(\rWrData[29] ),
    .B(net619),
    .Y(_01912_));
 sky130_fd_sc_hd__mux4_1 _06863_ (.A0(\reg_module.gprf[253] ),
    .A1(\reg_module.gprf[221] ),
    .A2(\reg_module.gprf[189] ),
    .A3(\reg_module.gprf[157] ),
    .S0(net1056),
    .S1(net1022),
    .X(_01913_));
 sky130_fd_sc_hd__mux4_1 _06864_ (.A0(\reg_module.gprf[125] ),
    .A1(\reg_module.gprf[93] ),
    .A2(\reg_module.gprf[61] ),
    .A3(\reg_module.gprf[29] ),
    .S0(net1056),
    .S1(net1022),
    .X(_01914_));
 sky130_fd_sc_hd__mux2_1 _06865_ (.A0(_01913_),
    .A1(_01914_),
    .S(net996),
    .X(_01915_));
 sky130_fd_sc_hd__mux4_1 _06866_ (.A0(\reg_module.gprf[381] ),
    .A1(\reg_module.gprf[349] ),
    .A2(\reg_module.gprf[317] ),
    .A3(\reg_module.gprf[285] ),
    .S0(net1056),
    .S1(net1022),
    .X(_01916_));
 sky130_fd_sc_hd__mux4_1 _06867_ (.A0(\reg_module.gprf[509] ),
    .A1(\reg_module.gprf[477] ),
    .A2(\reg_module.gprf[445] ),
    .A3(\reg_module.gprf[413] ),
    .S0(net1056),
    .S1(net1022),
    .X(_01917_));
 sky130_fd_sc_hd__mux2_1 _06868_ (.A0(_01916_),
    .A1(_01917_),
    .S(net832),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_1 _06869_ (.A0(_01915_),
    .A1(_01918_),
    .S(net822),
    .X(_01919_));
 sky130_fd_sc_hd__mux4_1 _06870_ (.A0(\reg_module.gprf[893] ),
    .A1(\reg_module.gprf[861] ),
    .A2(\reg_module.gprf[829] ),
    .A3(\reg_module.gprf[797] ),
    .S0(net1056),
    .S1(net1022),
    .X(_01920_));
 sky130_fd_sc_hd__or2_1 _06871_ (.A(net832),
    .B(_01920_),
    .X(_01921_));
 sky130_fd_sc_hd__mux4_1 _06872_ (.A0(\reg_module.gprf[1021] ),
    .A1(\reg_module.gprf[989] ),
    .A2(\reg_module.gprf[957] ),
    .A3(\reg_module.gprf[925] ),
    .S0(net1056),
    .S1(net1022),
    .X(_01922_));
 sky130_fd_sc_hd__o21a_1 _06873_ (.A1(net995),
    .A2(_01922_),
    .B1(net822),
    .X(_01923_));
 sky130_fd_sc_hd__mux4_1 _06874_ (.A0(\reg_module.gprf[765] ),
    .A1(\reg_module.gprf[733] ),
    .A2(\reg_module.gprf[701] ),
    .A3(\reg_module.gprf[669] ),
    .S0(net1056),
    .S1(net1022),
    .X(_01924_));
 sky130_fd_sc_hd__mux4_1 _06875_ (.A0(\reg_module.gprf[637] ),
    .A1(\reg_module.gprf[605] ),
    .A2(\reg_module.gprf[573] ),
    .A3(\reg_module.gprf[541] ),
    .S0(net1056),
    .S1(net1022),
    .X(_01925_));
 sky130_fd_sc_hd__mux2_1 _06876_ (.A0(_01924_),
    .A1(_01925_),
    .S(net995),
    .X(_01926_));
 sky130_fd_sc_hd__a221o_1 _06877_ (.A1(_01921_),
    .A2(_01923_),
    .B1(_01926_),
    .B2(net988),
    .C1(net1068),
    .X(_01927_));
 sky130_fd_sc_hd__o21a_1 _06878_ (.A1(net816),
    .A2(_01919_),
    .B1(_01927_),
    .X(_01928_));
 sky130_fd_sc_hd__o211ai_1 _06879_ (.A1(net817),
    .A2(_01919_),
    .B1(_01927_),
    .C1(net598),
    .Y(_01929_));
 sky130_fd_sc_hd__nand2_1 _06880_ (.A(\rWrDataWB[29] ),
    .B(net590),
    .Y(_01930_));
 sky130_fd_sc_hd__a31o_1 _06881_ (.A1(net619),
    .A2(_01929_),
    .A3(_01930_),
    .B1(_01912_),
    .X(_01931_));
 sky130_fd_sc_hd__nor2_1 _06882_ (.A(_01911_),
    .B(_01931_),
    .Y(_01932_));
 sky130_fd_sc_hd__or2_1 _06883_ (.A(_01284_),
    .B(_01932_),
    .X(_01933_));
 sky130_fd_sc_hd__a21oi_1 _06884_ (.A1(_01911_),
    .A2(_01931_),
    .B1(_01933_),
    .Y(net92));
 sky130_fd_sc_hd__mux4_1 _06885_ (.A0(\reg_module.gprf[382] ),
    .A1(\reg_module.gprf[350] ),
    .A2(\reg_module.gprf[318] ),
    .A3(\reg_module.gprf[286] ),
    .S0(net1059),
    .S1(net1025),
    .X(_01934_));
 sky130_fd_sc_hd__mux4_1 _06886_ (.A0(\reg_module.gprf[510] ),
    .A1(\reg_module.gprf[478] ),
    .A2(\reg_module.gprf[446] ),
    .A3(\reg_module.gprf[414] ),
    .S0(net1059),
    .S1(net1025),
    .X(_01935_));
 sky130_fd_sc_hd__mux4_1 _06887_ (.A0(\reg_module.gprf[126] ),
    .A1(\reg_module.gprf[94] ),
    .A2(\reg_module.gprf[62] ),
    .A3(\reg_module.gprf[30] ),
    .S0(net1059),
    .S1(net1025),
    .X(_01936_));
 sky130_fd_sc_hd__mux4_1 _06888_ (.A0(\reg_module.gprf[254] ),
    .A1(\reg_module.gprf[222] ),
    .A2(\reg_module.gprf[190] ),
    .A3(\reg_module.gprf[158] ),
    .S0(net1055),
    .S1(net1021),
    .X(_01937_));
 sky130_fd_sc_hd__mux4_1 _06889_ (.A0(_01934_),
    .A1(_01935_),
    .A2(_01936_),
    .A3(_01937_),
    .S0(net833),
    .S1(net991),
    .X(_01938_));
 sky130_fd_sc_hd__mux4_1 _06890_ (.A0(\reg_module.gprf[638] ),
    .A1(\reg_module.gprf[606] ),
    .A2(\reg_module.gprf[574] ),
    .A3(\reg_module.gprf[542] ),
    .S0(net1059),
    .S1(net1025),
    .X(_01939_));
 sky130_fd_sc_hd__or2_1 _06891_ (.A(net833),
    .B(_01939_),
    .X(_01940_));
 sky130_fd_sc_hd__mux4_1 _06892_ (.A0(\reg_module.gprf[766] ),
    .A1(\reg_module.gprf[734] ),
    .A2(\reg_module.gprf[702] ),
    .A3(\reg_module.gprf[670] ),
    .S0(net1055),
    .S1(net1021),
    .X(_01941_));
 sky130_fd_sc_hd__o21a_1 _06893_ (.A1(net995),
    .A2(_01941_),
    .B1(net988),
    .X(_01942_));
 sky130_fd_sc_hd__mux4_1 _06894_ (.A0(\reg_module.gprf[894] ),
    .A1(\reg_module.gprf[862] ),
    .A2(\reg_module.gprf[830] ),
    .A3(\reg_module.gprf[798] ),
    .S0(net1059),
    .S1(net1025),
    .X(_01943_));
 sky130_fd_sc_hd__mux4_1 _06895_ (.A0(\reg_module.gprf[1022] ),
    .A1(\reg_module.gprf[990] ),
    .A2(\reg_module.gprf[958] ),
    .A3(\reg_module.gprf[926] ),
    .S0(net1059),
    .S1(net1025),
    .X(_01944_));
 sky130_fd_sc_hd__mux2_1 _06896_ (.A0(_01943_),
    .A1(_01944_),
    .S(net833),
    .X(_01945_));
 sky130_fd_sc_hd__a221o_1 _06897_ (.A1(_01940_),
    .A2(_01942_),
    .B1(_01945_),
    .B2(net822),
    .C1(net1069),
    .X(_01946_));
 sky130_fd_sc_hd__o21a_1 _06898_ (.A1(net817),
    .A2(_01938_),
    .B1(_01946_),
    .X(_01947_));
 sky130_fd_sc_hd__o211a_1 _06899_ (.A1(net817),
    .A2(_01938_),
    .B1(_01946_),
    .C1(net598),
    .X(_01948_));
 sky130_fd_sc_hd__a21o_1 _06900_ (.A1(\rWrDataWB[30] ),
    .A2(net591),
    .B1(net625),
    .X(_01949_));
 sky130_fd_sc_hd__o22a_1 _06901_ (.A1(\rWrData[30] ),
    .A2(net619),
    .B1(_01948_),
    .B2(_01949_),
    .X(_01950_));
 sky130_fd_sc_hd__and2_1 _06902_ (.A(_01932_),
    .B(_01950_),
    .X(_01951_));
 sky130_fd_sc_hd__nor2_1 _06903_ (.A(_01284_),
    .B(_01951_),
    .Y(_01952_));
 sky130_fd_sc_hd__o21a_1 _06904_ (.A1(_01932_),
    .A2(_01950_),
    .B1(_01952_),
    .X(net94));
 sky130_fd_sc_hd__nor2_1 _06905_ (.A(\rWrData[31] ),
    .B(net620),
    .Y(_01953_));
 sky130_fd_sc_hd__mux4_1 _06906_ (.A0(\reg_module.gprf[383] ),
    .A1(\reg_module.gprf[351] ),
    .A2(\reg_module.gprf[319] ),
    .A3(\reg_module.gprf[287] ),
    .S0(net1061),
    .S1(net1027),
    .X(_01954_));
 sky130_fd_sc_hd__mux4_1 _06907_ (.A0(\reg_module.gprf[511] ),
    .A1(\reg_module.gprf[479] ),
    .A2(\reg_module.gprf[447] ),
    .A3(\reg_module.gprf[415] ),
    .S0(net1061),
    .S1(net1027),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _06908_ (.A0(_01954_),
    .A1(_01955_),
    .S(net834),
    .X(_01956_));
 sky130_fd_sc_hd__mux4_1 _06909_ (.A0(\reg_module.gprf[127] ),
    .A1(\reg_module.gprf[95] ),
    .A2(\reg_module.gprf[63] ),
    .A3(\reg_module.gprf[31] ),
    .S0(net1061),
    .S1(net1027),
    .X(_01957_));
 sky130_fd_sc_hd__mux4_1 _06910_ (.A0(\reg_module.gprf[255] ),
    .A1(\reg_module.gprf[223] ),
    .A2(\reg_module.gprf[191] ),
    .A3(\reg_module.gprf[159] ),
    .S0(net1061),
    .S1(net1027),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_1 _06911_ (.A0(_01957_),
    .A1(_01958_),
    .S(net833),
    .X(_01959_));
 sky130_fd_sc_hd__mux2_1 _06912_ (.A0(_01956_),
    .A1(_01959_),
    .S(net990),
    .X(_01960_));
 sky130_fd_sc_hd__mux4_1 _06913_ (.A0(\reg_module.gprf[895] ),
    .A1(\reg_module.gprf[863] ),
    .A2(\reg_module.gprf[831] ),
    .A3(\reg_module.gprf[799] ),
    .S0(net1061),
    .S1(net1027),
    .X(_01961_));
 sky130_fd_sc_hd__mux4_1 _06914_ (.A0(\reg_module.gprf[1023] ),
    .A1(\reg_module.gprf[991] ),
    .A2(\reg_module.gprf[959] ),
    .A3(\reg_module.gprf[927] ),
    .S0(net1061),
    .S1(net1027),
    .X(_01962_));
 sky130_fd_sc_hd__mux2_1 _06915_ (.A0(_01961_),
    .A1(_01962_),
    .S(net834),
    .X(_01963_));
 sky130_fd_sc_hd__mux4_1 _06916_ (.A0(\reg_module.gprf[767] ),
    .A1(\reg_module.gprf[735] ),
    .A2(\reg_module.gprf[703] ),
    .A3(\reg_module.gprf[671] ),
    .S0(net1060),
    .S1(net1026),
    .X(_01964_));
 sky130_fd_sc_hd__mux4_1 _06917_ (.A0(\reg_module.gprf[639] ),
    .A1(\reg_module.gprf[607] ),
    .A2(\reg_module.gprf[575] ),
    .A3(\reg_module.gprf[543] ),
    .S0(net1061),
    .S1(net1027),
    .X(_01965_));
 sky130_fd_sc_hd__mux2_1 _06918_ (.A0(_01964_),
    .A1(_01965_),
    .S(net997),
    .X(_01966_));
 sky130_fd_sc_hd__nand2_1 _06919_ (.A(net991),
    .B(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__a21oi_1 _06920_ (.A1(net822),
    .A2(_01963_),
    .B1(net1069),
    .Y(_01968_));
 sky130_fd_sc_hd__a2bb2o_1 _06921_ (.A1_N(net817),
    .A2_N(_01960_),
    .B1(_01967_),
    .B2(_01968_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _06922_ (.A0(_01215_),
    .A1(_01969_),
    .S(net600),
    .X(_01970_));
 sky130_fd_sc_hd__a21oi_2 _06923_ (.A1(net620),
    .A2(_01970_),
    .B1(_01953_),
    .Y(_01971_));
 sky130_fd_sc_hd__o21ai_1 _06924_ (.A1(_01951_),
    .A2(_01971_),
    .B1(net771),
    .Y(_01972_));
 sky130_fd_sc_hd__a21oi_1 _06925_ (.A1(_01951_),
    .A2(_01971_),
    .B1(_01972_),
    .Y(net95));
 sky130_fd_sc_hd__nor2_2 _06926_ (.A(\rWrData[0] ),
    .B(net602),
    .Y(_01973_));
 sky130_fd_sc_hd__o21a_2 _06927_ (.A1(\rReg_d2[4] ),
    .A2(_01254_),
    .B1(rRegWrEn2),
    .X(_01974_));
 sky130_fd_sc_hd__xor2_1 _06928_ (.A(\rReg_d2[0] ),
    .B(net917),
    .X(_01975_));
 sky130_fd_sc_hd__xnor2_1 _06929_ (.A(net968),
    .B(net860),
    .Y(_01976_));
 sky130_fd_sc_hd__or2_1 _06930_ (.A(net969),
    .B(net880),
    .X(_01977_));
 sky130_fd_sc_hd__nand2_1 _06931_ (.A(net969),
    .B(net880),
    .Y(_01978_));
 sky130_fd_sc_hd__nor2_1 _06932_ (.A(net966),
    .B(net851),
    .Y(_01979_));
 sky130_fd_sc_hd__and2_1 _06933_ (.A(net966),
    .B(net851),
    .X(_01980_));
 sky130_fd_sc_hd__nor2_1 _06934_ (.A(\rReg_d2[4] ),
    .B(net939),
    .Y(_01981_));
 sky130_fd_sc_hd__and2_1 _06935_ (.A(\rReg_d2[4] ),
    .B(net939),
    .X(_01982_));
 sky130_fd_sc_hd__o221a_1 _06936_ (.A1(_01979_),
    .A2(_01980_),
    .B1(_01981_),
    .B2(_01982_),
    .C1(_01976_),
    .X(_01983_));
 sky130_fd_sc_hd__a21oi_2 _06937_ (.A1(_01977_),
    .A2(_01978_),
    .B1(_01975_),
    .Y(_01984_));
 sky130_fd_sc_hd__a31oi_4 _06938_ (.A1(_01974_),
    .A2(_01983_),
    .A3(_01984_),
    .B1(rHazardStallRs2),
    .Y(_01985_));
 sky130_fd_sc_hd__a31o_1 _06939_ (.A1(_01974_),
    .A2(_01983_),
    .A3(_01984_),
    .B1(rHazardStallRs2),
    .X(_01986_));
 sky130_fd_sc_hd__mux4_1 _06940_ (.A0(\reg_module.gprf[480] ),
    .A1(\reg_module.gprf[448] ),
    .A2(\reg_module.gprf[416] ),
    .A3(\reg_module.gprf[384] ),
    .S0(net915),
    .S1(net878),
    .X(_01987_));
 sky130_fd_sc_hd__mux4_1 _06941_ (.A0(\reg_module.gprf[352] ),
    .A1(\reg_module.gprf[320] ),
    .A2(\reg_module.gprf[288] ),
    .A3(\reg_module.gprf[256] ),
    .S0(net915),
    .S1(net878),
    .X(_01988_));
 sky130_fd_sc_hd__mux2_1 _06942_ (.A0(_01987_),
    .A1(_01988_),
    .S(net857),
    .X(_01989_));
 sky130_fd_sc_hd__mux2_1 _06943_ (.A0(\reg_module.gprf[32] ),
    .A1(\reg_module.gprf[0] ),
    .S(net905),
    .X(_01990_));
 sky130_fd_sc_hd__nand2b_1 _06944_ (.A_N(\reg_module.gprf[64] ),
    .B(net906),
    .Y(_01991_));
 sky130_fd_sc_hd__o21ba_1 _06945_ (.A1(\reg_module.gprf[96] ),
    .A2(net905),
    .B1_N(net868),
    .X(_01992_));
 sky130_fd_sc_hd__a221o_1 _06946_ (.A1(net869),
    .A2(_01990_),
    .B1(_01991_),
    .B2(_01992_),
    .C1(net797),
    .X(_01993_));
 sky130_fd_sc_hd__mux4_1 _06947_ (.A0(\reg_module.gprf[224] ),
    .A1(\reg_module.gprf[192] ),
    .A2(\reg_module.gprf[160] ),
    .A3(\reg_module.gprf[128] ),
    .S0(net905),
    .S1(net868),
    .X(_01994_));
 sky130_fd_sc_hd__o21a_1 _06948_ (.A1(net858),
    .A2(_01994_),
    .B1(net848),
    .X(_01995_));
 sky130_fd_sc_hd__a221o_1 _06949_ (.A1(net788),
    .A2(_01989_),
    .B1(_01993_),
    .B2(_01995_),
    .C1(net783),
    .X(_01996_));
 sky130_fd_sc_hd__mux4_1 _06950_ (.A0(\reg_module.gprf[992] ),
    .A1(\reg_module.gprf[960] ),
    .A2(\reg_module.gprf[928] ),
    .A3(\reg_module.gprf[896] ),
    .S0(net915),
    .S1(net878),
    .X(_01997_));
 sky130_fd_sc_hd__mux4_1 _06951_ (.A0(\reg_module.gprf[864] ),
    .A1(\reg_module.gprf[832] ),
    .A2(\reg_module.gprf[800] ),
    .A3(\reg_module.gprf[768] ),
    .S0(net915),
    .S1(net878),
    .X(_01998_));
 sky130_fd_sc_hd__mux2_1 _06952_ (.A0(_01997_),
    .A1(_01998_),
    .S(net860),
    .X(_01999_));
 sky130_fd_sc_hd__mux4_1 _06953_ (.A0(\reg_module.gprf[736] ),
    .A1(\reg_module.gprf[704] ),
    .A2(\reg_module.gprf[672] ),
    .A3(\reg_module.gprf[640] ),
    .S0(net906),
    .S1(net869),
    .X(_02000_));
 sky130_fd_sc_hd__mux4_1 _06954_ (.A0(\reg_module.gprf[608] ),
    .A1(\reg_module.gprf[576] ),
    .A2(\reg_module.gprf[544] ),
    .A3(\reg_module.gprf[512] ),
    .S0(net912),
    .S1(net875),
    .X(_02001_));
 sky130_fd_sc_hd__or2_1 _06955_ (.A(net798),
    .B(_02001_),
    .X(_02002_));
 sky130_fd_sc_hd__o21a_1 _06956_ (.A1(net858),
    .A2(_02000_),
    .B1(net848),
    .X(_02003_));
 sky130_fd_sc_hd__a221o_1 _06957_ (.A1(net787),
    .A2(_01999_),
    .B1(_02002_),
    .B2(_02003_),
    .C1(net938),
    .X(_02004_));
 sky130_fd_sc_hd__a21o_1 _06958_ (.A1(_01996_),
    .A2(_02004_),
    .B1(net575),
    .X(_02005_));
 sky130_fd_sc_hd__o21ai_1 _06959_ (.A1(\rWrDataWB[0] ),
    .A2(net584),
    .B1(_02005_),
    .Y(_02006_));
 sky130_fd_sc_hd__a21oi_2 _06960_ (.A1(net602),
    .A2(_02006_),
    .B1(_01973_),
    .Y(net103));
 sky130_fd_sc_hd__and2_1 _06961_ (.A(\rWrData[1] ),
    .B(net610),
    .X(_02007_));
 sky130_fd_sc_hd__mux4_1 _06962_ (.A0(\reg_module.gprf[865] ),
    .A1(\reg_module.gprf[833] ),
    .A2(\reg_module.gprf[801] ),
    .A3(\reg_module.gprf[769] ),
    .S0(net916),
    .S1(net879),
    .X(_02008_));
 sky130_fd_sc_hd__mux4_1 _06963_ (.A0(\reg_module.gprf[993] ),
    .A1(\reg_module.gprf[961] ),
    .A2(\reg_module.gprf[929] ),
    .A3(\reg_module.gprf[897] ),
    .S0(net917),
    .S1(net880),
    .X(_02009_));
 sky130_fd_sc_hd__or2_1 _06964_ (.A(net860),
    .B(_02009_),
    .X(_02010_));
 sky130_fd_sc_hd__o21a_1 _06965_ (.A1(net802),
    .A2(_02008_),
    .B1(net790),
    .X(_02011_));
 sky130_fd_sc_hd__mux4_1 _06966_ (.A0(\reg_module.gprf[609] ),
    .A1(\reg_module.gprf[577] ),
    .A2(\reg_module.gprf[545] ),
    .A3(\reg_module.gprf[513] ),
    .S0(net917),
    .S1(net881),
    .X(_02012_));
 sky130_fd_sc_hd__mux4_1 _06967_ (.A0(\reg_module.gprf[737] ),
    .A1(\reg_module.gprf[705] ),
    .A2(\reg_module.gprf[673] ),
    .A3(\reg_module.gprf[641] ),
    .S0(net918),
    .S1(net881),
    .X(_02013_));
 sky130_fd_sc_hd__mux2_1 _06968_ (.A0(_02012_),
    .A1(_02013_),
    .S(net802),
    .X(_02014_));
 sky130_fd_sc_hd__a221o_1 _06969_ (.A1(_02010_),
    .A2(_02011_),
    .B1(_02014_),
    .B2(net852),
    .C1(net939),
    .X(_02015_));
 sky130_fd_sc_hd__mux4_1 _06970_ (.A0(\reg_module.gprf[353] ),
    .A1(\reg_module.gprf[321] ),
    .A2(\reg_module.gprf[289] ),
    .A3(\reg_module.gprf[257] ),
    .S0(net916),
    .S1(net879),
    .X(_02016_));
 sky130_fd_sc_hd__or2_1 _06971_ (.A(net801),
    .B(_02016_),
    .X(_02017_));
 sky130_fd_sc_hd__mux4_1 _06972_ (.A0(\reg_module.gprf[481] ),
    .A1(\reg_module.gprf[449] ),
    .A2(\reg_module.gprf[417] ),
    .A3(\reg_module.gprf[385] ),
    .S0(net917),
    .S1(net881),
    .X(_02018_));
 sky130_fd_sc_hd__o211a_1 _06973_ (.A1(net860),
    .A2(_02018_),
    .B1(_02017_),
    .C1(net790),
    .X(_02019_));
 sky130_fd_sc_hd__mux4_1 _06974_ (.A0(\reg_module.gprf[97] ),
    .A1(\reg_module.gprf[65] ),
    .A2(\reg_module.gprf[33] ),
    .A3(\reg_module.gprf[1] ),
    .S0(net916),
    .S1(net879),
    .X(_02020_));
 sky130_fd_sc_hd__mux4_1 _06975_ (.A0(\reg_module.gprf[225] ),
    .A1(\reg_module.gprf[193] ),
    .A2(\reg_module.gprf[161] ),
    .A3(\reg_module.gprf[129] ),
    .S0(net917),
    .S1(net879),
    .X(_02021_));
 sky130_fd_sc_hd__mux2_1 _06976_ (.A0(_02020_),
    .A1(_02021_),
    .S(net802),
    .X(_02022_));
 sky130_fd_sc_hd__a21o_1 _06977_ (.A1(net852),
    .A2(_02022_),
    .B1(net784),
    .X(_02023_));
 sky130_fd_sc_hd__o211a_1 _06978_ (.A1(_02019_),
    .A2(_02023_),
    .B1(net584),
    .C1(_02015_),
    .X(_02024_));
 sky130_fd_sc_hd__a21o_1 _06979_ (.A1(\rWrDataWB[1] ),
    .A2(net577),
    .B1(_02024_),
    .X(_02025_));
 sky130_fd_sc_hd__a21o_1 _06980_ (.A1(net602),
    .A2(_02025_),
    .B1(_02007_),
    .X(net114));
 sky130_fd_sc_hd__nand2_1 _06981_ (.A(\rWrData[2] ),
    .B(net610),
    .Y(_02026_));
 sky130_fd_sc_hd__mux4_1 _06982_ (.A0(\reg_module.gprf[866] ),
    .A1(\reg_module.gprf[834] ),
    .A2(\reg_module.gprf[802] ),
    .A3(\reg_module.gprf[770] ),
    .S0(net912),
    .S1(net875),
    .X(_02027_));
 sky130_fd_sc_hd__or2_1 _06983_ (.A(net797),
    .B(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__mux4_1 _06984_ (.A0(\reg_module.gprf[994] ),
    .A1(\reg_module.gprf[962] ),
    .A2(\reg_module.gprf[930] ),
    .A3(\reg_module.gprf[898] ),
    .S0(net912),
    .S1(net875),
    .X(_02029_));
 sky130_fd_sc_hd__o21a_1 _06985_ (.A1(net858),
    .A2(_02029_),
    .B1(net788),
    .X(_02030_));
 sky130_fd_sc_hd__mux4_1 _06986_ (.A0(\reg_module.gprf[610] ),
    .A1(\reg_module.gprf[578] ),
    .A2(\reg_module.gprf[546] ),
    .A3(\reg_module.gprf[514] ),
    .S0(net905),
    .S1(net868),
    .X(_02031_));
 sky130_fd_sc_hd__mux4_1 _06987_ (.A0(\reg_module.gprf[738] ),
    .A1(\reg_module.gprf[706] ),
    .A2(\reg_module.gprf[674] ),
    .A3(\reg_module.gprf[642] ),
    .S0(net905),
    .S1(net868),
    .X(_02032_));
 sky130_fd_sc_hd__mux2_1 _06988_ (.A0(_02031_),
    .A1(_02032_),
    .S(net797),
    .X(_02033_));
 sky130_fd_sc_hd__a221oi_1 _06989_ (.A1(_02028_),
    .A2(_02030_),
    .B1(_02033_),
    .B2(net850),
    .C1(net938),
    .Y(_02034_));
 sky130_fd_sc_hd__mux4_1 _06990_ (.A0(\reg_module.gprf[226] ),
    .A1(\reg_module.gprf[194] ),
    .A2(\reg_module.gprf[162] ),
    .A3(\reg_module.gprf[130] ),
    .S0(net912),
    .S1(net875),
    .X(_02035_));
 sky130_fd_sc_hd__mux4_1 _06991_ (.A0(\reg_module.gprf[98] ),
    .A1(\reg_module.gprf[66] ),
    .A2(\reg_module.gprf[34] ),
    .A3(\reg_module.gprf[2] ),
    .S0(net912),
    .S1(net875),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _06992_ (.A0(_02035_),
    .A1(_02036_),
    .S(net859),
    .X(_02037_));
 sky130_fd_sc_hd__nand2_1 _06993_ (.A(net849),
    .B(_02037_),
    .Y(_02038_));
 sky130_fd_sc_hd__mux4_1 _06994_ (.A0(\reg_module.gprf[354] ),
    .A1(\reg_module.gprf[322] ),
    .A2(\reg_module.gprf[290] ),
    .A3(\reg_module.gprf[258] ),
    .S0(net912),
    .S1(net875),
    .X(_02039_));
 sky130_fd_sc_hd__mux4_1 _06995_ (.A0(\reg_module.gprf[482] ),
    .A1(\reg_module.gprf[450] ),
    .A2(\reg_module.gprf[418] ),
    .A3(\reg_module.gprf[386] ),
    .S0(net912),
    .S1(net875),
    .X(_02040_));
 sky130_fd_sc_hd__mux2_1 _06996_ (.A0(_02039_),
    .A1(_02040_),
    .S(net800),
    .X(_02041_));
 sky130_fd_sc_hd__nand2_1 _06997_ (.A(net789),
    .B(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__a311o_2 _06998_ (.A1(net939),
    .A2(_02038_),
    .A3(_02042_),
    .B1(net576),
    .C1(_02034_),
    .X(_02043_));
 sky130_fd_sc_hd__nand2_1 _06999_ (.A(\rWrDataWB[2] ),
    .B(net577),
    .Y(_02044_));
 sky130_fd_sc_hd__a21o_1 _07000_ (.A1(_02043_),
    .A2(_02044_),
    .B1(net611),
    .X(_02045_));
 sky130_fd_sc_hd__nand2_1 _07001_ (.A(_02026_),
    .B(_02045_),
    .Y(net125));
 sky130_fd_sc_hd__mux4_1 _07002_ (.A0(\reg_module.gprf[867] ),
    .A1(\reg_module.gprf[835] ),
    .A2(\reg_module.gprf[803] ),
    .A3(\reg_module.gprf[771] ),
    .S0(net905),
    .S1(net868),
    .X(_02046_));
 sky130_fd_sc_hd__mux4_1 _07003_ (.A0(\reg_module.gprf[995] ),
    .A1(\reg_module.gprf[963] ),
    .A2(\reg_module.gprf[931] ),
    .A3(\reg_module.gprf[899] ),
    .S0(net906),
    .S1(net868),
    .X(_02047_));
 sky130_fd_sc_hd__or2_1 _07004_ (.A(net858),
    .B(_02047_),
    .X(_02048_));
 sky130_fd_sc_hd__o21a_1 _07005_ (.A1(net797),
    .A2(_02046_),
    .B1(net787),
    .X(_02049_));
 sky130_fd_sc_hd__mux4_1 _07006_ (.A0(\reg_module.gprf[611] ),
    .A1(\reg_module.gprf[579] ),
    .A2(\reg_module.gprf[547] ),
    .A3(\reg_module.gprf[515] ),
    .S0(net905),
    .S1(net868),
    .X(_02050_));
 sky130_fd_sc_hd__mux4_1 _07007_ (.A0(\reg_module.gprf[739] ),
    .A1(\reg_module.gprf[707] ),
    .A2(\reg_module.gprf[675] ),
    .A3(\reg_module.gprf[643] ),
    .S0(net905),
    .S1(net868),
    .X(_02051_));
 sky130_fd_sc_hd__mux2_1 _07008_ (.A0(_02050_),
    .A1(_02051_),
    .S(net797),
    .X(_02052_));
 sky130_fd_sc_hd__a221o_1 _07009_ (.A1(_02048_),
    .A2(_02049_),
    .B1(_02052_),
    .B2(net850),
    .C1(net938),
    .X(_02053_));
 sky130_fd_sc_hd__mux4_1 _07010_ (.A0(\reg_module.gprf[355] ),
    .A1(\reg_module.gprf[323] ),
    .A2(\reg_module.gprf[291] ),
    .A3(\reg_module.gprf[259] ),
    .S0(net905),
    .S1(net868),
    .X(_02054_));
 sky130_fd_sc_hd__or2_1 _07011_ (.A(net798),
    .B(_02054_),
    .X(_02055_));
 sky130_fd_sc_hd__mux4_1 _07012_ (.A0(\reg_module.gprf[483] ),
    .A1(\reg_module.gprf[451] ),
    .A2(\reg_module.gprf[419] ),
    .A3(\reg_module.gprf[387] ),
    .S0(net905),
    .S1(net868),
    .X(_02056_));
 sky130_fd_sc_hd__o211a_1 _07013_ (.A1(net858),
    .A2(_02056_),
    .B1(_02055_),
    .C1(net788),
    .X(_02057_));
 sky130_fd_sc_hd__mux4_1 _07014_ (.A0(\reg_module.gprf[99] ),
    .A1(\reg_module.gprf[67] ),
    .A2(\reg_module.gprf[35] ),
    .A3(\reg_module.gprf[3] ),
    .S0(net907),
    .S1(net866),
    .X(_02058_));
 sky130_fd_sc_hd__mux4_1 _07015_ (.A0(\reg_module.gprf[227] ),
    .A1(\reg_module.gprf[195] ),
    .A2(\reg_module.gprf[163] ),
    .A3(\reg_module.gprf[131] ),
    .S0(net907),
    .S1(net870),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _07016_ (.A0(_02058_),
    .A1(_02059_),
    .S(net796),
    .X(_02060_));
 sky130_fd_sc_hd__a21o_1 _07017_ (.A1(net848),
    .A2(_02060_),
    .B1(net783),
    .X(_02061_));
 sky130_fd_sc_hd__o211a_1 _07018_ (.A1(_02057_),
    .A2(_02061_),
    .B1(net583),
    .C1(_02053_),
    .X(_02062_));
 sky130_fd_sc_hd__a21o_1 _07019_ (.A1(\rWrDataWB[3] ),
    .A2(net577),
    .B1(_02062_),
    .X(_02063_));
 sky130_fd_sc_hd__mux2_1 _07020_ (.A0(\rWrData[3] ),
    .A1(_02063_),
    .S(net602),
    .X(net128));
 sky130_fd_sc_hd__nand2_2 _07021_ (.A(\rWrData[4] ),
    .B(net610),
    .Y(_02064_));
 sky130_fd_sc_hd__mux4_1 _07022_ (.A0(\reg_module.gprf[868] ),
    .A1(\reg_module.gprf[836] ),
    .A2(\reg_module.gprf[804] ),
    .A3(\reg_module.gprf[772] ),
    .S0(net916),
    .S1(net880),
    .X(_02065_));
 sky130_fd_sc_hd__mux4_1 _07023_ (.A0(\reg_module.gprf[996] ),
    .A1(\reg_module.gprf[964] ),
    .A2(\reg_module.gprf[932] ),
    .A3(\reg_module.gprf[900] ),
    .S0(net917),
    .S1(net880),
    .X(_02066_));
 sky130_fd_sc_hd__mux2_1 _07024_ (.A0(_02065_),
    .A1(_02066_),
    .S(net801),
    .X(_02067_));
 sky130_fd_sc_hd__mux4_1 _07025_ (.A0(\reg_module.gprf[612] ),
    .A1(\reg_module.gprf[580] ),
    .A2(\reg_module.gprf[548] ),
    .A3(\reg_module.gprf[516] ),
    .S0(net916),
    .S1(net879),
    .X(_02068_));
 sky130_fd_sc_hd__mux4_1 _07026_ (.A0(\reg_module.gprf[740] ),
    .A1(\reg_module.gprf[708] ),
    .A2(\reg_module.gprf[676] ),
    .A3(\reg_module.gprf[644] ),
    .S0(net916),
    .S1(net879),
    .X(_02069_));
 sky130_fd_sc_hd__mux2_1 _07027_ (.A0(_02068_),
    .A1(_02069_),
    .S(net801),
    .X(_02070_));
 sky130_fd_sc_hd__a21o_1 _07028_ (.A1(net790),
    .A2(_02067_),
    .B1(net939),
    .X(_02071_));
 sky130_fd_sc_hd__a21o_1 _07029_ (.A1(net852),
    .A2(_02070_),
    .B1(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__mux4_1 _07030_ (.A0(\reg_module.gprf[228] ),
    .A1(\reg_module.gprf[196] ),
    .A2(\reg_module.gprf[164] ),
    .A3(\reg_module.gprf[132] ),
    .S0(net916),
    .S1(net879),
    .X(_02073_));
 sky130_fd_sc_hd__mux4_1 _07031_ (.A0(\reg_module.gprf[100] ),
    .A1(\reg_module.gprf[68] ),
    .A2(\reg_module.gprf[36] ),
    .A3(\reg_module.gprf[4] ),
    .S0(net916),
    .S1(net879),
    .X(_02074_));
 sky130_fd_sc_hd__mux2_1 _07032_ (.A0(_02073_),
    .A1(_02074_),
    .S(net860),
    .X(_02075_));
 sky130_fd_sc_hd__mux4_1 _07033_ (.A0(\reg_module.gprf[356] ),
    .A1(\reg_module.gprf[324] ),
    .A2(\reg_module.gprf[292] ),
    .A3(\reg_module.gprf[260] ),
    .S0(net916),
    .S1(net879),
    .X(_02076_));
 sky130_fd_sc_hd__mux4_1 _07034_ (.A0(\reg_module.gprf[484] ),
    .A1(\reg_module.gprf[452] ),
    .A2(\reg_module.gprf[420] ),
    .A3(\reg_module.gprf[388] ),
    .S0(net917),
    .S1(net880),
    .X(_02077_));
 sky130_fd_sc_hd__mux2_1 _07035_ (.A0(_02076_),
    .A1(_02077_),
    .S(net802),
    .X(_02078_));
 sky130_fd_sc_hd__a21o_1 _07036_ (.A1(net790),
    .A2(_02078_),
    .B1(net784),
    .X(_02079_));
 sky130_fd_sc_hd__a21o_1 _07037_ (.A1(net852),
    .A2(_02075_),
    .B1(_02079_),
    .X(_02080_));
 sky130_fd_sc_hd__and3_1 _07038_ (.A(net584),
    .B(_02072_),
    .C(_02080_),
    .X(_02081_));
 sky130_fd_sc_hd__a21o_1 _07039_ (.A1(\rWrDataWB[4] ),
    .A2(net577),
    .B1(_02081_),
    .X(_02082_));
 sky130_fd_sc_hd__a21bo_1 _07040_ (.A1(net602),
    .A2(_02082_),
    .B1_N(_02064_),
    .X(net129));
 sky130_fd_sc_hd__mux4_1 _07041_ (.A0(\reg_module.gprf[869] ),
    .A1(\reg_module.gprf[837] ),
    .A2(\reg_module.gprf[805] ),
    .A3(\reg_module.gprf[773] ),
    .S0(net914),
    .S1(net877),
    .X(_02083_));
 sky130_fd_sc_hd__or2_1 _07042_ (.A(net801),
    .B(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__mux4_1 _07043_ (.A0(\reg_module.gprf[997] ),
    .A1(\reg_module.gprf[965] ),
    .A2(\reg_module.gprf[933] ),
    .A3(\reg_module.gprf[901] ),
    .S0(net914),
    .S1(net877),
    .X(_02085_));
 sky130_fd_sc_hd__o21a_1 _07044_ (.A1(net860),
    .A2(_02085_),
    .B1(net790),
    .X(_02086_));
 sky130_fd_sc_hd__mux4_1 _07045_ (.A0(\reg_module.gprf[613] ),
    .A1(\reg_module.gprf[581] ),
    .A2(\reg_module.gprf[549] ),
    .A3(\reg_module.gprf[517] ),
    .S0(net914),
    .S1(net877),
    .X(_02087_));
 sky130_fd_sc_hd__mux4_1 _07046_ (.A0(\reg_module.gprf[741] ),
    .A1(\reg_module.gprf[709] ),
    .A2(\reg_module.gprf[677] ),
    .A3(\reg_module.gprf[645] ),
    .S0(net904),
    .S1(net867),
    .X(_02088_));
 sky130_fd_sc_hd__mux2_1 _07047_ (.A0(_02087_),
    .A1(_02088_),
    .S(net797),
    .X(_02089_));
 sky130_fd_sc_hd__a221o_1 _07048_ (.A1(_02084_),
    .A2(_02086_),
    .B1(_02089_),
    .B2(net851),
    .C1(net940),
    .X(_02090_));
 sky130_fd_sc_hd__mux4_1 _07049_ (.A0(\reg_module.gprf[357] ),
    .A1(\reg_module.gprf[325] ),
    .A2(\reg_module.gprf[293] ),
    .A3(\reg_module.gprf[261] ),
    .S0(net914),
    .S1(net877),
    .X(_02091_));
 sky130_fd_sc_hd__mux4_1 _07050_ (.A0(\reg_module.gprf[485] ),
    .A1(\reg_module.gprf[453] ),
    .A2(\reg_module.gprf[421] ),
    .A3(\reg_module.gprf[389] ),
    .S0(net914),
    .S1(net877),
    .X(_02092_));
 sky130_fd_sc_hd__mux2_1 _07051_ (.A0(_02091_),
    .A1(_02092_),
    .S(net801),
    .X(_02093_));
 sky130_fd_sc_hd__mux4_1 _07052_ (.A0(\reg_module.gprf[101] ),
    .A1(\reg_module.gprf[69] ),
    .A2(\reg_module.gprf[37] ),
    .A3(\reg_module.gprf[5] ),
    .S0(net914),
    .S1(net877),
    .X(_02094_));
 sky130_fd_sc_hd__or2_1 _07053_ (.A(net801),
    .B(_02094_),
    .X(_02095_));
 sky130_fd_sc_hd__mux4_1 _07054_ (.A0(\reg_module.gprf[229] ),
    .A1(\reg_module.gprf[197] ),
    .A2(\reg_module.gprf[165] ),
    .A3(\reg_module.gprf[133] ),
    .S0(net914),
    .S1(net877),
    .X(_02096_));
 sky130_fd_sc_hd__o211a_1 _07055_ (.A1(net860),
    .A2(_02096_),
    .B1(_02095_),
    .C1(net851),
    .X(_02097_));
 sky130_fd_sc_hd__a21o_1 _07056_ (.A1(net790),
    .A2(_02093_),
    .B1(net784),
    .X(_02098_));
 sky130_fd_sc_hd__o211a_1 _07057_ (.A1(_02097_),
    .A2(_02098_),
    .B1(net584),
    .C1(_02090_),
    .X(_02099_));
 sky130_fd_sc_hd__a21o_1 _07058_ (.A1(\rWrDataWB[5] ),
    .A2(net577),
    .B1(net610),
    .X(_02100_));
 sky130_fd_sc_hd__o22a_1 _07059_ (.A1(\rWrData[5] ),
    .A2(net602),
    .B1(_02099_),
    .B2(_02100_),
    .X(net130));
 sky130_fd_sc_hd__mux4_1 _07060_ (.A0(\reg_module.gprf[870] ),
    .A1(\reg_module.gprf[838] ),
    .A2(\reg_module.gprf[806] ),
    .A3(\reg_module.gprf[774] ),
    .S0(net904),
    .S1(net867),
    .X(_02101_));
 sky130_fd_sc_hd__mux4_1 _07061_ (.A0(\reg_module.gprf[998] ),
    .A1(\reg_module.gprf[966] ),
    .A2(\reg_module.gprf[934] ),
    .A3(\reg_module.gprf[902] ),
    .S0(net904),
    .S1(net867),
    .X(_02102_));
 sky130_fd_sc_hd__or2_1 _07062_ (.A(net857),
    .B(_02102_),
    .X(_02103_));
 sky130_fd_sc_hd__o21a_1 _07063_ (.A1(net795),
    .A2(_02101_),
    .B1(net787),
    .X(_02104_));
 sky130_fd_sc_hd__mux4_1 _07064_ (.A0(\reg_module.gprf[614] ),
    .A1(\reg_module.gprf[582] ),
    .A2(\reg_module.gprf[550] ),
    .A3(\reg_module.gprf[518] ),
    .S0(net903),
    .S1(net866),
    .X(_02105_));
 sky130_fd_sc_hd__mux4_1 _07065_ (.A0(\reg_module.gprf[742] ),
    .A1(\reg_module.gprf[710] ),
    .A2(\reg_module.gprf[678] ),
    .A3(\reg_module.gprf[646] ),
    .S0(net903),
    .S1(net866),
    .X(_02106_));
 sky130_fd_sc_hd__mux2_1 _07066_ (.A0(_02105_),
    .A1(_02106_),
    .S(net795),
    .X(_02107_));
 sky130_fd_sc_hd__a221o_1 _07067_ (.A1(_02103_),
    .A2(_02104_),
    .B1(_02107_),
    .B2(net848),
    .C1(net938),
    .X(_02108_));
 sky130_fd_sc_hd__mux4_1 _07068_ (.A0(\reg_module.gprf[358] ),
    .A1(\reg_module.gprf[326] ),
    .A2(\reg_module.gprf[294] ),
    .A3(\reg_module.gprf[262] ),
    .S0(net903),
    .S1(net866),
    .X(_02109_));
 sky130_fd_sc_hd__mux4_1 _07069_ (.A0(\reg_module.gprf[486] ),
    .A1(\reg_module.gprf[454] ),
    .A2(\reg_module.gprf[422] ),
    .A3(\reg_module.gprf[390] ),
    .S0(net904),
    .S1(net867),
    .X(_02110_));
 sky130_fd_sc_hd__mux2_1 _07070_ (.A0(_02109_),
    .A1(_02110_),
    .S(net795),
    .X(_02111_));
 sky130_fd_sc_hd__mux4_1 _07071_ (.A0(\reg_module.gprf[102] ),
    .A1(\reg_module.gprf[70] ),
    .A2(\reg_module.gprf[38] ),
    .A3(\reg_module.gprf[6] ),
    .S0(net903),
    .S1(net866),
    .X(_02112_));
 sky130_fd_sc_hd__mux4_1 _07072_ (.A0(\reg_module.gprf[230] ),
    .A1(\reg_module.gprf[198] ),
    .A2(\reg_module.gprf[166] ),
    .A3(\reg_module.gprf[134] ),
    .S0(net903),
    .S1(net866),
    .X(_02113_));
 sky130_fd_sc_hd__or2_1 _07073_ (.A(net857),
    .B(_02113_),
    .X(_02114_));
 sky130_fd_sc_hd__o211a_1 _07074_ (.A1(net795),
    .A2(_02112_),
    .B1(_02114_),
    .C1(net848),
    .X(_02115_));
 sky130_fd_sc_hd__a21o_1 _07075_ (.A1(net787),
    .A2(_02111_),
    .B1(net783),
    .X(_02116_));
 sky130_fd_sc_hd__o211a_1 _07076_ (.A1(_02115_),
    .A2(_02116_),
    .B1(net583),
    .C1(_02108_),
    .X(_02117_));
 sky130_fd_sc_hd__a21o_1 _07077_ (.A1(\rWrDataWB[6] ),
    .A2(net575),
    .B1(net609),
    .X(_02118_));
 sky130_fd_sc_hd__o22a_1 _07078_ (.A1(\rWrData[6] ),
    .A2(net601),
    .B1(_02117_),
    .B2(_02118_),
    .X(net131));
 sky130_fd_sc_hd__mux4_1 _07079_ (.A0(\reg_module.gprf[871] ),
    .A1(\reg_module.gprf[839] ),
    .A2(\reg_module.gprf[807] ),
    .A3(\reg_module.gprf[775] ),
    .S0(net906),
    .S1(net869),
    .X(_02119_));
 sky130_fd_sc_hd__mux4_1 _07080_ (.A0(\reg_module.gprf[999] ),
    .A1(\reg_module.gprf[967] ),
    .A2(\reg_module.gprf[935] ),
    .A3(\reg_module.gprf[903] ),
    .S0(net904),
    .S1(net867),
    .X(_02120_));
 sky130_fd_sc_hd__or2_1 _07081_ (.A(net858),
    .B(_02120_),
    .X(_02121_));
 sky130_fd_sc_hd__o21a_1 _07082_ (.A1(net797),
    .A2(_02119_),
    .B1(net788),
    .X(_02122_));
 sky130_fd_sc_hd__mux4_1 _07083_ (.A0(\reg_module.gprf[615] ),
    .A1(\reg_module.gprf[583] ),
    .A2(\reg_module.gprf[551] ),
    .A3(\reg_module.gprf[519] ),
    .S0(net904),
    .S1(net867),
    .X(_02123_));
 sky130_fd_sc_hd__mux4_1 _07084_ (.A0(\reg_module.gprf[743] ),
    .A1(\reg_module.gprf[711] ),
    .A2(\reg_module.gprf[679] ),
    .A3(\reg_module.gprf[647] ),
    .S0(net904),
    .S1(net867),
    .X(_02124_));
 sky130_fd_sc_hd__mux2_1 _07085_ (.A0(_02123_),
    .A1(_02124_),
    .S(net797),
    .X(_02125_));
 sky130_fd_sc_hd__a221o_1 _07086_ (.A1(_02121_),
    .A2(_02122_),
    .B1(_02125_),
    .B2(net850),
    .C1(net938),
    .X(_02126_));
 sky130_fd_sc_hd__mux4_1 _07087_ (.A0(\reg_module.gprf[359] ),
    .A1(\reg_module.gprf[327] ),
    .A2(\reg_module.gprf[295] ),
    .A3(\reg_module.gprf[263] ),
    .S0(net906),
    .S1(net869),
    .X(_02127_));
 sky130_fd_sc_hd__mux4_1 _07088_ (.A0(\reg_module.gprf[487] ),
    .A1(\reg_module.gprf[455] ),
    .A2(\reg_module.gprf[423] ),
    .A3(\reg_module.gprf[391] ),
    .S0(net904),
    .S1(net867),
    .X(_02128_));
 sky130_fd_sc_hd__mux2_1 _07089_ (.A0(_02127_),
    .A1(_02128_),
    .S(net797),
    .X(_02129_));
 sky130_fd_sc_hd__mux4_1 _07090_ (.A0(\reg_module.gprf[103] ),
    .A1(\reg_module.gprf[71] ),
    .A2(\reg_module.gprf[39] ),
    .A3(\reg_module.gprf[7] ),
    .S0(net904),
    .S1(net867),
    .X(_02130_));
 sky130_fd_sc_hd__or2_1 _07091_ (.A(net797),
    .B(_02130_),
    .X(_02131_));
 sky130_fd_sc_hd__mux4_1 _07092_ (.A0(\reg_module.gprf[231] ),
    .A1(\reg_module.gprf[199] ),
    .A2(\reg_module.gprf[167] ),
    .A3(\reg_module.gprf[135] ),
    .S0(net904),
    .S1(net867),
    .X(_02132_));
 sky130_fd_sc_hd__o211a_1 _07093_ (.A1(net857),
    .A2(_02132_),
    .B1(_02131_),
    .C1(net850),
    .X(_02133_));
 sky130_fd_sc_hd__a21o_1 _07094_ (.A1(net788),
    .A2(_02129_),
    .B1(net783),
    .X(_02134_));
 sky130_fd_sc_hd__o211a_1 _07095_ (.A1(_02133_),
    .A2(_02134_),
    .B1(net583),
    .C1(_02126_),
    .X(_02135_));
 sky130_fd_sc_hd__a21o_1 _07096_ (.A1(\rWrDataWB[7] ),
    .A2(net575),
    .B1(net609),
    .X(_02136_));
 sky130_fd_sc_hd__o22a_1 _07097_ (.A1(\rWrData[7] ),
    .A2(net601),
    .B1(_02135_),
    .B2(_02136_),
    .X(net132));
 sky130_fd_sc_hd__mux4_1 _07098_ (.A0(\reg_module.gprf[872] ),
    .A1(\reg_module.gprf[840] ),
    .A2(\reg_module.gprf[808] ),
    .A3(\reg_module.gprf[776] ),
    .S0(net916),
    .S1(net879),
    .X(_02137_));
 sky130_fd_sc_hd__or2_1 _07099_ (.A(net801),
    .B(_02137_),
    .X(_02138_));
 sky130_fd_sc_hd__mux4_1 _07100_ (.A0(\reg_module.gprf[1000] ),
    .A1(\reg_module.gprf[968] ),
    .A2(\reg_module.gprf[936] ),
    .A3(\reg_module.gprf[904] ),
    .S0(net915),
    .S1(net877),
    .X(_02139_));
 sky130_fd_sc_hd__o21a_1 _07101_ (.A1(net860),
    .A2(_02139_),
    .B1(net790),
    .X(_02140_));
 sky130_fd_sc_hd__mux4_1 _07102_ (.A0(\reg_module.gprf[616] ),
    .A1(\reg_module.gprf[584] ),
    .A2(\reg_module.gprf[552] ),
    .A3(\reg_module.gprf[520] ),
    .S0(net915),
    .S1(net878),
    .X(_02141_));
 sky130_fd_sc_hd__mux4_1 _07103_ (.A0(\reg_module.gprf[744] ),
    .A1(\reg_module.gprf[712] ),
    .A2(\reg_module.gprf[680] ),
    .A3(\reg_module.gprf[648] ),
    .S0(net914),
    .S1(net877),
    .X(_02142_));
 sky130_fd_sc_hd__mux2_1 _07104_ (.A0(_02141_),
    .A1(_02142_),
    .S(net801),
    .X(_02143_));
 sky130_fd_sc_hd__a221o_1 _07105_ (.A1(_02138_),
    .A2(_02140_),
    .B1(_02143_),
    .B2(net851),
    .C1(net940),
    .X(_02144_));
 sky130_fd_sc_hd__mux4_1 _07106_ (.A0(\reg_module.gprf[360] ),
    .A1(\reg_module.gprf[328] ),
    .A2(\reg_module.gprf[296] ),
    .A3(\reg_module.gprf[264] ),
    .S0(net914),
    .S1(net877),
    .X(_02145_));
 sky130_fd_sc_hd__mux4_1 _07107_ (.A0(\reg_module.gprf[488] ),
    .A1(\reg_module.gprf[456] ),
    .A2(\reg_module.gprf[424] ),
    .A3(\reg_module.gprf[392] ),
    .S0(net915),
    .S1(net878),
    .X(_02146_));
 sky130_fd_sc_hd__mux2_1 _07108_ (.A0(_02145_),
    .A1(_02146_),
    .S(net801),
    .X(_02147_));
 sky130_fd_sc_hd__mux4_1 _07109_ (.A0(\reg_module.gprf[104] ),
    .A1(\reg_module.gprf[72] ),
    .A2(\reg_module.gprf[40] ),
    .A3(\reg_module.gprf[8] ),
    .S0(net914),
    .S1(net878),
    .X(_02148_));
 sky130_fd_sc_hd__or2_1 _07110_ (.A(net801),
    .B(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__mux4_1 _07111_ (.A0(\reg_module.gprf[232] ),
    .A1(\reg_module.gprf[200] ),
    .A2(\reg_module.gprf[168] ),
    .A3(\reg_module.gprf[136] ),
    .S0(net915),
    .S1(net878),
    .X(_02150_));
 sky130_fd_sc_hd__o211a_1 _07112_ (.A1(net860),
    .A2(_02150_),
    .B1(_02149_),
    .C1(net851),
    .X(_02151_));
 sky130_fd_sc_hd__a21o_1 _07113_ (.A1(net794),
    .A2(_02147_),
    .B1(net784),
    .X(_02152_));
 sky130_fd_sc_hd__o211a_1 _07114_ (.A1(_02151_),
    .A2(_02152_),
    .B1(net584),
    .C1(_02144_),
    .X(_02153_));
 sky130_fd_sc_hd__a21o_1 _07115_ (.A1(\rWrDataWB[8] ),
    .A2(net577),
    .B1(net610),
    .X(_02154_));
 sky130_fd_sc_hd__o22a_1 _07116_ (.A1(\rWrData[8] ),
    .A2(net602),
    .B1(_02153_),
    .B2(_02154_),
    .X(net133));
 sky130_fd_sc_hd__mux4_1 _07117_ (.A0(\reg_module.gprf[873] ),
    .A1(\reg_module.gprf[841] ),
    .A2(\reg_module.gprf[809] ),
    .A3(\reg_module.gprf[777] ),
    .S0(net902),
    .S1(net865),
    .X(_02155_));
 sky130_fd_sc_hd__or2_1 _07118_ (.A(net796),
    .B(_02155_),
    .X(_02156_));
 sky130_fd_sc_hd__mux4_1 _07119_ (.A0(\reg_module.gprf[1001] ),
    .A1(\reg_module.gprf[969] ),
    .A2(\reg_module.gprf[937] ),
    .A3(\reg_module.gprf[905] ),
    .S0(net902),
    .S1(net865),
    .X(_02157_));
 sky130_fd_sc_hd__o21a_1 _07120_ (.A1(net857),
    .A2(_02157_),
    .B1(net787),
    .X(_02158_));
 sky130_fd_sc_hd__mux4_1 _07121_ (.A0(\reg_module.gprf[617] ),
    .A1(\reg_module.gprf[585] ),
    .A2(\reg_module.gprf[553] ),
    .A3(\reg_module.gprf[521] ),
    .S0(net907),
    .S1(net870),
    .X(_02159_));
 sky130_fd_sc_hd__mux4_1 _07122_ (.A0(\reg_module.gprf[745] ),
    .A1(\reg_module.gprf[713] ),
    .A2(\reg_module.gprf[681] ),
    .A3(\reg_module.gprf[649] ),
    .S0(net902),
    .S1(net865),
    .X(_02160_));
 sky130_fd_sc_hd__mux2_1 _07123_ (.A0(_02159_),
    .A1(_02160_),
    .S(net796),
    .X(_02161_));
 sky130_fd_sc_hd__a221o_1 _07124_ (.A1(_02156_),
    .A2(_02158_),
    .B1(_02161_),
    .B2(net848),
    .C1(net938),
    .X(_02162_));
 sky130_fd_sc_hd__mux4_1 _07125_ (.A0(\reg_module.gprf[361] ),
    .A1(\reg_module.gprf[329] ),
    .A2(\reg_module.gprf[297] ),
    .A3(\reg_module.gprf[265] ),
    .S0(net908),
    .S1(net871),
    .X(_02163_));
 sky130_fd_sc_hd__mux4_1 _07126_ (.A0(\reg_module.gprf[489] ),
    .A1(\reg_module.gprf[457] ),
    .A2(\reg_module.gprf[425] ),
    .A3(\reg_module.gprf[393] ),
    .S0(net902),
    .S1(net865),
    .X(_02164_));
 sky130_fd_sc_hd__mux2_1 _07127_ (.A0(_02163_),
    .A1(_02164_),
    .S(net796),
    .X(_02165_));
 sky130_fd_sc_hd__mux4_1 _07128_ (.A0(\reg_module.gprf[105] ),
    .A1(\reg_module.gprf[73] ),
    .A2(\reg_module.gprf[41] ),
    .A3(\reg_module.gprf[9] ),
    .S0(net908),
    .S1(net871),
    .X(_02166_));
 sky130_fd_sc_hd__mux4_1 _07129_ (.A0(\reg_module.gprf[233] ),
    .A1(\reg_module.gprf[201] ),
    .A2(\reg_module.gprf[169] ),
    .A3(\reg_module.gprf[137] ),
    .S0(net908),
    .S1(net871),
    .X(_02167_));
 sky130_fd_sc_hd__or2_1 _07130_ (.A(net857),
    .B(_02167_),
    .X(_02168_));
 sky130_fd_sc_hd__o211a_1 _07131_ (.A1(net795),
    .A2(_02166_),
    .B1(_02168_),
    .C1(net849),
    .X(_02169_));
 sky130_fd_sc_hd__a21o_1 _07132_ (.A1(net787),
    .A2(_02165_),
    .B1(net783),
    .X(_02170_));
 sky130_fd_sc_hd__o211a_1 _07133_ (.A1(_02169_),
    .A2(_02170_),
    .B1(net583),
    .C1(_02162_),
    .X(_02171_));
 sky130_fd_sc_hd__a21o_1 _07134_ (.A1(\rWrDataWB[9] ),
    .A2(net575),
    .B1(net609),
    .X(_02172_));
 sky130_fd_sc_hd__o22a_1 _07135_ (.A1(\rWrData[9] ),
    .A2(net601),
    .B1(_02171_),
    .B2(_02172_),
    .X(net134));
 sky130_fd_sc_hd__mux4_1 _07136_ (.A0(\reg_module.gprf[874] ),
    .A1(\reg_module.gprf[842] ),
    .A2(\reg_module.gprf[810] ),
    .A3(\reg_module.gprf[778] ),
    .S0(net902),
    .S1(net865),
    .X(_02173_));
 sky130_fd_sc_hd__mux4_1 _07137_ (.A0(\reg_module.gprf[1002] ),
    .A1(\reg_module.gprf[970] ),
    .A2(\reg_module.gprf[938] ),
    .A3(\reg_module.gprf[906] ),
    .S0(net903),
    .S1(net866),
    .X(_02174_));
 sky130_fd_sc_hd__or2_1 _07138_ (.A(net857),
    .B(_02174_),
    .X(_02175_));
 sky130_fd_sc_hd__o21a_1 _07139_ (.A1(net795),
    .A2(_02173_),
    .B1(net787),
    .X(_02176_));
 sky130_fd_sc_hd__mux4_1 _07140_ (.A0(\reg_module.gprf[618] ),
    .A1(\reg_module.gprf[586] ),
    .A2(\reg_module.gprf[554] ),
    .A3(\reg_module.gprf[522] ),
    .S0(net902),
    .S1(net865),
    .X(_02177_));
 sky130_fd_sc_hd__mux4_1 _07141_ (.A0(\reg_module.gprf[746] ),
    .A1(\reg_module.gprf[714] ),
    .A2(\reg_module.gprf[682] ),
    .A3(\reg_module.gprf[650] ),
    .S0(net903),
    .S1(net866),
    .X(_02178_));
 sky130_fd_sc_hd__mux2_1 _07142_ (.A0(_02177_),
    .A1(_02178_),
    .S(net795),
    .X(_02179_));
 sky130_fd_sc_hd__a221o_1 _07143_ (.A1(_02175_),
    .A2(_02176_),
    .B1(_02179_),
    .B2(net848),
    .C1(net938),
    .X(_02180_));
 sky130_fd_sc_hd__mux4_1 _07144_ (.A0(\reg_module.gprf[362] ),
    .A1(\reg_module.gprf[330] ),
    .A2(\reg_module.gprf[298] ),
    .A3(\reg_module.gprf[266] ),
    .S0(net902),
    .S1(net865),
    .X(_02181_));
 sky130_fd_sc_hd__mux4_1 _07145_ (.A0(\reg_module.gprf[490] ),
    .A1(\reg_module.gprf[458] ),
    .A2(\reg_module.gprf[426] ),
    .A3(\reg_module.gprf[394] ),
    .S0(net902),
    .S1(net865),
    .X(_02182_));
 sky130_fd_sc_hd__mux2_1 _07146_ (.A0(_02181_),
    .A1(_02182_),
    .S(net795),
    .X(_02183_));
 sky130_fd_sc_hd__mux4_1 _07147_ (.A0(\reg_module.gprf[106] ),
    .A1(\reg_module.gprf[74] ),
    .A2(\reg_module.gprf[42] ),
    .A3(\reg_module.gprf[10] ),
    .S0(net902),
    .S1(net865),
    .X(_02184_));
 sky130_fd_sc_hd__mux4_1 _07148_ (.A0(\reg_module.gprf[234] ),
    .A1(\reg_module.gprf[202] ),
    .A2(\reg_module.gprf[170] ),
    .A3(\reg_module.gprf[138] ),
    .S0(net903),
    .S1(net866),
    .X(_02185_));
 sky130_fd_sc_hd__or2_1 _07149_ (.A(net857),
    .B(_02185_),
    .X(_02186_));
 sky130_fd_sc_hd__o211a_1 _07150_ (.A1(net795),
    .A2(_02184_),
    .B1(_02186_),
    .C1(net848),
    .X(_02187_));
 sky130_fd_sc_hd__a21o_1 _07151_ (.A1(net787),
    .A2(_02183_),
    .B1(net783),
    .X(_02188_));
 sky130_fd_sc_hd__o211a_2 _07152_ (.A1(_02187_),
    .A2(_02188_),
    .B1(net583),
    .C1(_02180_),
    .X(_02189_));
 sky130_fd_sc_hd__a21o_1 _07153_ (.A1(\rWrDataWB[10] ),
    .A2(net575),
    .B1(net609),
    .X(_02190_));
 sky130_fd_sc_hd__o22a_1 _07154_ (.A1(\rWrData[10] ),
    .A2(net601),
    .B1(_02189_),
    .B2(_02190_),
    .X(net104));
 sky130_fd_sc_hd__mux4_1 _07155_ (.A0(\reg_module.gprf[875] ),
    .A1(\reg_module.gprf[843] ),
    .A2(\reg_module.gprf[811] ),
    .A3(\reg_module.gprf[779] ),
    .S0(net908),
    .S1(net871),
    .X(_02191_));
 sky130_fd_sc_hd__mux4_1 _07156_ (.A0(\reg_module.gprf[1003] ),
    .A1(\reg_module.gprf[971] ),
    .A2(\reg_module.gprf[939] ),
    .A3(\reg_module.gprf[907] ),
    .S0(net908),
    .S1(net871),
    .X(_02192_));
 sky130_fd_sc_hd__or2_1 _07157_ (.A(net859),
    .B(_02192_),
    .X(_02193_));
 sky130_fd_sc_hd__o21a_1 _07158_ (.A1(net799),
    .A2(_02191_),
    .B1(net790),
    .X(_02194_));
 sky130_fd_sc_hd__mux4_1 _07159_ (.A0(\reg_module.gprf[619] ),
    .A1(\reg_module.gprf[587] ),
    .A2(\reg_module.gprf[555] ),
    .A3(\reg_module.gprf[523] ),
    .S0(net908),
    .S1(net871),
    .X(_02195_));
 sky130_fd_sc_hd__mux4_1 _07160_ (.A0(\reg_module.gprf[747] ),
    .A1(\reg_module.gprf[715] ),
    .A2(\reg_module.gprf[683] ),
    .A3(\reg_module.gprf[651] ),
    .S0(net908),
    .S1(net871),
    .X(_02196_));
 sky130_fd_sc_hd__mux2_1 _07161_ (.A0(_02195_),
    .A1(_02196_),
    .S(net799),
    .X(_02197_));
 sky130_fd_sc_hd__a221o_1 _07162_ (.A1(_02193_),
    .A2(_02194_),
    .B1(_02197_),
    .B2(net849),
    .C1(net939),
    .X(_02198_));
 sky130_fd_sc_hd__mux4_1 _07163_ (.A0(\reg_module.gprf[363] ),
    .A1(\reg_module.gprf[331] ),
    .A2(\reg_module.gprf[299] ),
    .A3(\reg_module.gprf[267] ),
    .S0(net909),
    .S1(net872),
    .X(_02199_));
 sky130_fd_sc_hd__mux4_1 _07164_ (.A0(\reg_module.gprf[491] ),
    .A1(\reg_module.gprf[459] ),
    .A2(\reg_module.gprf[427] ),
    .A3(\reg_module.gprf[395] ),
    .S0(net909),
    .S1(net872),
    .X(_02200_));
 sky130_fd_sc_hd__mux2_1 _07165_ (.A0(_02199_),
    .A1(_02200_),
    .S(net799),
    .X(_02201_));
 sky130_fd_sc_hd__mux4_1 _07166_ (.A0(\reg_module.gprf[107] ),
    .A1(\reg_module.gprf[75] ),
    .A2(\reg_module.gprf[43] ),
    .A3(\reg_module.gprf[11] ),
    .S0(net909),
    .S1(net872),
    .X(_02202_));
 sky130_fd_sc_hd__or2_1 _07167_ (.A(net799),
    .B(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__mux4_1 _07168_ (.A0(\reg_module.gprf[235] ),
    .A1(\reg_module.gprf[203] ),
    .A2(\reg_module.gprf[171] ),
    .A3(\reg_module.gprf[139] ),
    .S0(net909),
    .S1(net872),
    .X(_02204_));
 sky130_fd_sc_hd__o211a_1 _07169_ (.A1(net859),
    .A2(_02204_),
    .B1(_02203_),
    .C1(net849),
    .X(_02205_));
 sky130_fd_sc_hd__a21o_1 _07170_ (.A1(net789),
    .A2(_02201_),
    .B1(net783),
    .X(_02206_));
 sky130_fd_sc_hd__o211a_1 _07171_ (.A1(_02205_),
    .A2(_02206_),
    .B1(net583),
    .C1(_02198_),
    .X(_02207_));
 sky130_fd_sc_hd__a21o_1 _07172_ (.A1(\rWrDataWB[11] ),
    .A2(net575),
    .B1(net611),
    .X(_02208_));
 sky130_fd_sc_hd__o22a_1 _07173_ (.A1(\rWrData[11] ),
    .A2(net604),
    .B1(_02207_),
    .B2(_02208_),
    .X(net105));
 sky130_fd_sc_hd__or2_1 _07174_ (.A(\rWrData[12] ),
    .B(net604),
    .X(_02209_));
 sky130_fd_sc_hd__mux4_1 _07175_ (.A0(\reg_module.gprf[748] ),
    .A1(\reg_module.gprf[716] ),
    .A2(\reg_module.gprf[684] ),
    .A3(\reg_module.gprf[652] ),
    .S0(net909),
    .S1(net872),
    .X(_02210_));
 sky130_fd_sc_hd__mux4_1 _07176_ (.A0(\reg_module.gprf[620] ),
    .A1(\reg_module.gprf[588] ),
    .A2(\reg_module.gprf[556] ),
    .A3(\reg_module.gprf[524] ),
    .S0(net910),
    .S1(net873),
    .X(_02211_));
 sky130_fd_sc_hd__mux2_1 _07177_ (.A0(_02210_),
    .A1(_02211_),
    .S(net859),
    .X(_02212_));
 sky130_fd_sc_hd__mux4_1 _07178_ (.A0(\reg_module.gprf[876] ),
    .A1(\reg_module.gprf[844] ),
    .A2(\reg_module.gprf[812] ),
    .A3(\reg_module.gprf[780] ),
    .S0(net921),
    .S1(net885),
    .X(_02213_));
 sky130_fd_sc_hd__mux4_1 _07179_ (.A0(\reg_module.gprf[1004] ),
    .A1(\reg_module.gprf[972] ),
    .A2(\reg_module.gprf[940] ),
    .A3(\reg_module.gprf[908] ),
    .S0(net923),
    .S1(net887),
    .X(_02214_));
 sky130_fd_sc_hd__mux2_1 _07180_ (.A0(_02213_),
    .A1(_02214_),
    .S(net804),
    .X(_02215_));
 sky130_fd_sc_hd__a21o_1 _07181_ (.A1(net789),
    .A2(_02215_),
    .B1(net938),
    .X(_02216_));
 sky130_fd_sc_hd__a21o_1 _07182_ (.A1(net849),
    .A2(_02212_),
    .B1(_02216_),
    .X(_02217_));
 sky130_fd_sc_hd__mux4_1 _07183_ (.A0(\reg_module.gprf[364] ),
    .A1(\reg_module.gprf[332] ),
    .A2(\reg_module.gprf[300] ),
    .A3(\reg_module.gprf[268] ),
    .S0(net909),
    .S1(net872),
    .X(_02218_));
 sky130_fd_sc_hd__mux4_1 _07184_ (.A0(\reg_module.gprf[492] ),
    .A1(\reg_module.gprf[460] ),
    .A2(\reg_module.gprf[428] ),
    .A3(\reg_module.gprf[396] ),
    .S0(net911),
    .S1(net874),
    .X(_02219_));
 sky130_fd_sc_hd__mux2_1 _07185_ (.A0(_02218_),
    .A1(_02219_),
    .S(net799),
    .X(_02220_));
 sky130_fd_sc_hd__mux4_1 _07186_ (.A0(\reg_module.gprf[108] ),
    .A1(\reg_module.gprf[76] ),
    .A2(\reg_module.gprf[44] ),
    .A3(\reg_module.gprf[12] ),
    .S0(net909),
    .S1(net872),
    .X(_02221_));
 sky130_fd_sc_hd__mux4_1 _07187_ (.A0(\reg_module.gprf[236] ),
    .A1(\reg_module.gprf[204] ),
    .A2(\reg_module.gprf[172] ),
    .A3(\reg_module.gprf[140] ),
    .S0(net910),
    .S1(net873),
    .X(_02222_));
 sky130_fd_sc_hd__mux2_1 _07188_ (.A0(_02221_),
    .A1(_02222_),
    .S(net799),
    .X(_02223_));
 sky130_fd_sc_hd__a21o_1 _07189_ (.A1(net849),
    .A2(_02223_),
    .B1(net784),
    .X(_02224_));
 sky130_fd_sc_hd__a21o_1 _07190_ (.A1(net789),
    .A2(_02220_),
    .B1(_02224_),
    .X(_02225_));
 sky130_fd_sc_hd__and2_1 _07191_ (.A(\rWrDataWB[12] ),
    .B(net576),
    .X(_02226_));
 sky130_fd_sc_hd__a31o_1 _07192_ (.A1(net583),
    .A2(_02217_),
    .A3(_02225_),
    .B1(_02226_),
    .X(_02227_));
 sky130_fd_sc_hd__o21a_2 _07193_ (.A1(net611),
    .A2(_02227_),
    .B1(_02209_),
    .X(net106));
 sky130_fd_sc_hd__mux4_1 _07194_ (.A0(\reg_module.gprf[877] ),
    .A1(\reg_module.gprf[845] ),
    .A2(\reg_module.gprf[813] ),
    .A3(\reg_module.gprf[781] ),
    .S0(net903),
    .S1(net870),
    .X(_02228_));
 sky130_fd_sc_hd__or2_1 _07195_ (.A(net796),
    .B(_02228_),
    .X(_02229_));
 sky130_fd_sc_hd__mux4_1 _07196_ (.A0(\reg_module.gprf[1005] ),
    .A1(\reg_module.gprf[973] ),
    .A2(\reg_module.gprf[941] ),
    .A3(\reg_module.gprf[909] ),
    .S0(net902),
    .S1(net865),
    .X(_02230_));
 sky130_fd_sc_hd__o21a_1 _07197_ (.A1(net857),
    .A2(_02230_),
    .B1(net787),
    .X(_02231_));
 sky130_fd_sc_hd__mux4_1 _07198_ (.A0(\reg_module.gprf[621] ),
    .A1(\reg_module.gprf[589] ),
    .A2(\reg_module.gprf[557] ),
    .A3(\reg_module.gprf[525] ),
    .S0(net912),
    .S1(net875),
    .X(_02232_));
 sky130_fd_sc_hd__mux4_1 _07199_ (.A0(\reg_module.gprf[749] ),
    .A1(\reg_module.gprf[717] ),
    .A2(\reg_module.gprf[685] ),
    .A3(\reg_module.gprf[653] ),
    .S0(net908),
    .S1(net871),
    .X(_02233_));
 sky130_fd_sc_hd__mux2_1 _07200_ (.A0(_02232_),
    .A1(_02233_),
    .S(net799),
    .X(_02234_));
 sky130_fd_sc_hd__a221o_1 _07201_ (.A1(_02229_),
    .A2(_02231_),
    .B1(_02234_),
    .B2(net848),
    .C1(net938),
    .X(_02235_));
 sky130_fd_sc_hd__mux4_1 _07202_ (.A0(\reg_module.gprf[365] ),
    .A1(\reg_module.gprf[333] ),
    .A2(\reg_module.gprf[301] ),
    .A3(\reg_module.gprf[269] ),
    .S0(net912),
    .S1(net875),
    .X(_02236_));
 sky130_fd_sc_hd__mux4_1 _07203_ (.A0(\reg_module.gprf[493] ),
    .A1(\reg_module.gprf[461] ),
    .A2(\reg_module.gprf[429] ),
    .A3(\reg_module.gprf[397] ),
    .S0(net908),
    .S1(net873),
    .X(_02237_));
 sky130_fd_sc_hd__mux2_1 _07204_ (.A0(_02236_),
    .A1(_02237_),
    .S(net795),
    .X(_02238_));
 sky130_fd_sc_hd__mux4_1 _07205_ (.A0(\reg_module.gprf[109] ),
    .A1(\reg_module.gprf[77] ),
    .A2(\reg_module.gprf[45] ),
    .A3(\reg_module.gprf[13] ),
    .S0(net910),
    .S1(net871),
    .X(_02239_));
 sky130_fd_sc_hd__or2_1 _07206_ (.A(net799),
    .B(_02239_),
    .X(_02240_));
 sky130_fd_sc_hd__mux4_1 _07207_ (.A0(\reg_module.gprf[237] ),
    .A1(\reg_module.gprf[205] ),
    .A2(\reg_module.gprf[173] ),
    .A3(\reg_module.gprf[141] ),
    .S0(net908),
    .S1(net871),
    .X(_02241_));
 sky130_fd_sc_hd__o211a_1 _07208_ (.A1(net859),
    .A2(_02241_),
    .B1(_02240_),
    .C1(net849),
    .X(_02242_));
 sky130_fd_sc_hd__a21o_1 _07209_ (.A1(net787),
    .A2(_02238_),
    .B1(net783),
    .X(_02243_));
 sky130_fd_sc_hd__o211a_1 _07210_ (.A1(_02242_),
    .A2(_02243_),
    .B1(net583),
    .C1(_02235_),
    .X(_02244_));
 sky130_fd_sc_hd__a21o_1 _07211_ (.A1(\rWrDataWB[13] ),
    .A2(net576),
    .B1(net611),
    .X(_02245_));
 sky130_fd_sc_hd__o22a_1 _07212_ (.A1(\rWrData[13] ),
    .A2(net601),
    .B1(_02244_),
    .B2(_02245_),
    .X(net107));
 sky130_fd_sc_hd__mux4_1 _07213_ (.A0(\reg_module.gprf[750] ),
    .A1(\reg_module.gprf[718] ),
    .A2(\reg_module.gprf[686] ),
    .A3(\reg_module.gprf[654] ),
    .S0(net911),
    .S1(net874),
    .X(_02246_));
 sky130_fd_sc_hd__mux4_1 _07214_ (.A0(\reg_module.gprf[622] ),
    .A1(\reg_module.gprf[590] ),
    .A2(\reg_module.gprf[558] ),
    .A3(\reg_module.gprf[526] ),
    .S0(net913),
    .S1(net876),
    .X(_02247_));
 sky130_fd_sc_hd__or2_1 _07215_ (.A(net800),
    .B(_02247_),
    .X(_02248_));
 sky130_fd_sc_hd__o21a_1 _07216_ (.A1(net861),
    .A2(_02246_),
    .B1(net849),
    .X(_02249_));
 sky130_fd_sc_hd__mux4_1 _07217_ (.A0(\reg_module.gprf[878] ),
    .A1(\reg_module.gprf[846] ),
    .A2(\reg_module.gprf[814] ),
    .A3(\reg_module.gprf[782] ),
    .S0(net911),
    .S1(net874),
    .X(_02250_));
 sky130_fd_sc_hd__mux4_1 _07218_ (.A0(\reg_module.gprf[1006] ),
    .A1(\reg_module.gprf[974] ),
    .A2(\reg_module.gprf[942] ),
    .A3(\reg_module.gprf[910] ),
    .S0(net911),
    .S1(net874),
    .X(_02251_));
 sky130_fd_sc_hd__mux2_1 _07219_ (.A0(_02250_),
    .A1(_02251_),
    .S(net800),
    .X(_02252_));
 sky130_fd_sc_hd__a221o_1 _07220_ (.A1(_02248_),
    .A2(_02249_),
    .B1(_02252_),
    .B2(net789),
    .C1(net939),
    .X(_02253_));
 sky130_fd_sc_hd__mux4_1 _07221_ (.A0(\reg_module.gprf[366] ),
    .A1(\reg_module.gprf[334] ),
    .A2(\reg_module.gprf[302] ),
    .A3(\reg_module.gprf[270] ),
    .S0(net923),
    .S1(net887),
    .X(_02254_));
 sky130_fd_sc_hd__mux4_1 _07222_ (.A0(\reg_module.gprf[494] ),
    .A1(\reg_module.gprf[462] ),
    .A2(\reg_module.gprf[430] ),
    .A3(\reg_module.gprf[398] ),
    .S0(net936),
    .S1(net900),
    .X(_02255_));
 sky130_fd_sc_hd__mux2_1 _07223_ (.A0(_02254_),
    .A1(_02255_),
    .S(net800),
    .X(_02256_));
 sky130_fd_sc_hd__mux4_1 _07224_ (.A0(\reg_module.gprf[110] ),
    .A1(\reg_module.gprf[78] ),
    .A2(\reg_module.gprf[46] ),
    .A3(\reg_module.gprf[14] ),
    .S0(net913),
    .S1(net876),
    .X(_02257_));
 sky130_fd_sc_hd__mux4_1 _07225_ (.A0(\reg_module.gprf[238] ),
    .A1(\reg_module.gprf[206] ),
    .A2(\reg_module.gprf[174] ),
    .A3(\reg_module.gprf[142] ),
    .S0(net912),
    .S1(net875),
    .X(_02258_));
 sky130_fd_sc_hd__or2_1 _07226_ (.A(net861),
    .B(_02258_),
    .X(_02259_));
 sky130_fd_sc_hd__o211a_1 _07227_ (.A1(net800),
    .A2(_02257_),
    .B1(_02259_),
    .C1(net849),
    .X(_02260_));
 sky130_fd_sc_hd__a21o_1 _07228_ (.A1(net789),
    .A2(_02256_),
    .B1(net783),
    .X(_02261_));
 sky130_fd_sc_hd__o211a_1 _07229_ (.A1(_02260_),
    .A2(_02261_),
    .B1(net583),
    .C1(_02253_),
    .X(_02262_));
 sky130_fd_sc_hd__a21o_1 _07230_ (.A1(\rWrDataWB[14] ),
    .A2(net581),
    .B1(net615),
    .X(_02263_));
 sky130_fd_sc_hd__o22a_2 _07231_ (.A1(\rWrData[14] ),
    .A2(net608),
    .B1(_02262_),
    .B2(_02263_),
    .X(net108));
 sky130_fd_sc_hd__mux4_1 _07232_ (.A0(\reg_module.gprf[879] ),
    .A1(\reg_module.gprf[847] ),
    .A2(\reg_module.gprf[815] ),
    .A3(\reg_module.gprf[783] ),
    .S0(net923),
    .S1(net887),
    .X(_02264_));
 sky130_fd_sc_hd__or2_1 _07233_ (.A(net806),
    .B(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__mux4_1 _07234_ (.A0(\reg_module.gprf[1007] ),
    .A1(\reg_module.gprf[975] ),
    .A2(\reg_module.gprf[943] ),
    .A3(\reg_module.gprf[911] ),
    .S0(net923),
    .S1(net887),
    .X(_02266_));
 sky130_fd_sc_hd__o21a_1 _07235_ (.A1(net862),
    .A2(_02266_),
    .B1(net791),
    .X(_02267_));
 sky130_fd_sc_hd__mux4_1 _07236_ (.A0(\reg_module.gprf[623] ),
    .A1(\reg_module.gprf[591] ),
    .A2(\reg_module.gprf[559] ),
    .A3(\reg_module.gprf[527] ),
    .S0(net923),
    .S1(net887),
    .X(_02268_));
 sky130_fd_sc_hd__mux4_1 _07237_ (.A0(\reg_module.gprf[751] ),
    .A1(\reg_module.gprf[719] ),
    .A2(\reg_module.gprf[687] ),
    .A3(\reg_module.gprf[655] ),
    .S0(net923),
    .S1(net887),
    .X(_02269_));
 sky130_fd_sc_hd__mux2_1 _07238_ (.A0(_02268_),
    .A1(_02269_),
    .S(net806),
    .X(_02270_));
 sky130_fd_sc_hd__a221o_1 _07239_ (.A1(_02265_),
    .A2(_02267_),
    .B1(_02270_),
    .B2(net853),
    .C1(net941),
    .X(_02271_));
 sky130_fd_sc_hd__mux4_1 _07240_ (.A0(\reg_module.gprf[367] ),
    .A1(\reg_module.gprf[335] ),
    .A2(\reg_module.gprf[303] ),
    .A3(\reg_module.gprf[271] ),
    .S0(net922),
    .S1(net886),
    .X(_02272_));
 sky130_fd_sc_hd__mux4_1 _07241_ (.A0(\reg_module.gprf[495] ),
    .A1(\reg_module.gprf[463] ),
    .A2(\reg_module.gprf[431] ),
    .A3(\reg_module.gprf[399] ),
    .S0(net922),
    .S1(net886),
    .X(_02273_));
 sky130_fd_sc_hd__mux2_1 _07242_ (.A0(_02272_),
    .A1(_02273_),
    .S(net806),
    .X(_02274_));
 sky130_fd_sc_hd__mux4_1 _07243_ (.A0(\reg_module.gprf[111] ),
    .A1(\reg_module.gprf[79] ),
    .A2(\reg_module.gprf[47] ),
    .A3(\reg_module.gprf[15] ),
    .S0(net923),
    .S1(net887),
    .X(_02275_));
 sky130_fd_sc_hd__mux4_1 _07244_ (.A0(\reg_module.gprf[239] ),
    .A1(\reg_module.gprf[207] ),
    .A2(\reg_module.gprf[175] ),
    .A3(\reg_module.gprf[143] ),
    .S0(net923),
    .S1(net887),
    .X(_02276_));
 sky130_fd_sc_hd__or2_1 _07245_ (.A(net862),
    .B(_02276_),
    .X(_02277_));
 sky130_fd_sc_hd__o211a_1 _07246_ (.A1(net806),
    .A2(_02275_),
    .B1(_02277_),
    .C1(net853),
    .X(_02278_));
 sky130_fd_sc_hd__a21o_1 _07247_ (.A1(net791),
    .A2(_02274_),
    .B1(net785),
    .X(_02279_));
 sky130_fd_sc_hd__o211a_1 _07248_ (.A1(_02278_),
    .A2(_02279_),
    .B1(net585),
    .C1(_02271_),
    .X(_02280_));
 sky130_fd_sc_hd__a21o_1 _07249_ (.A1(\rWrDataWB[15] ),
    .A2(net581),
    .B1(net613),
    .X(_02281_));
 sky130_fd_sc_hd__o22a_2 _07250_ (.A1(\rWrData[15] ),
    .A2(net605),
    .B1(_02280_),
    .B2(_02281_),
    .X(net109));
 sky130_fd_sc_hd__or2_1 _07251_ (.A(\rWrData[16] ),
    .B(net607),
    .X(_02282_));
 sky130_fd_sc_hd__mux4_1 _07252_ (.A0(\reg_module.gprf[880] ),
    .A1(\reg_module.gprf[848] ),
    .A2(\reg_module.gprf[816] ),
    .A3(\reg_module.gprf[784] ),
    .S0(net935),
    .S1(net899),
    .X(_02283_));
 sky130_fd_sc_hd__mux4_1 _07253_ (.A0(\reg_module.gprf[1008] ),
    .A1(\reg_module.gprf[976] ),
    .A2(\reg_module.gprf[944] ),
    .A3(\reg_module.gprf[912] ),
    .S0(net935),
    .S1(net899),
    .X(_02284_));
 sky130_fd_sc_hd__mux2_1 _07254_ (.A0(_02283_),
    .A1(_02284_),
    .S(net809),
    .X(_02285_));
 sky130_fd_sc_hd__mux4_1 _07255_ (.A0(\reg_module.gprf[624] ),
    .A1(\reg_module.gprf[592] ),
    .A2(\reg_module.gprf[560] ),
    .A3(\reg_module.gprf[528] ),
    .S0(net935),
    .S1(net899),
    .X(_02286_));
 sky130_fd_sc_hd__mux4_1 _07256_ (.A0(\reg_module.gprf[752] ),
    .A1(\reg_module.gprf[720] ),
    .A2(\reg_module.gprf[688] ),
    .A3(\reg_module.gprf[656] ),
    .S0(net935),
    .S1(net899),
    .X(_02287_));
 sky130_fd_sc_hd__or2_1 _07257_ (.A(net864),
    .B(_02287_),
    .X(_02288_));
 sky130_fd_sc_hd__o211a_1 _07258_ (.A1(net809),
    .A2(_02286_),
    .B1(_02288_),
    .C1(net855),
    .X(_02289_));
 sky130_fd_sc_hd__a211o_1 _07259_ (.A1(net794),
    .A2(_02285_),
    .B1(_02289_),
    .C1(net942),
    .X(_02290_));
 sky130_fd_sc_hd__mux4_1 _07260_ (.A0(\reg_module.gprf[368] ),
    .A1(\reg_module.gprf[336] ),
    .A2(\reg_module.gprf[304] ),
    .A3(\reg_module.gprf[272] ),
    .S0(net935),
    .S1(net899),
    .X(_02291_));
 sky130_fd_sc_hd__mux4_1 _07261_ (.A0(\reg_module.gprf[496] ),
    .A1(\reg_module.gprf[464] ),
    .A2(\reg_module.gprf[432] ),
    .A3(\reg_module.gprf[400] ),
    .S0(net935),
    .S1(net899),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _07262_ (.A0(_02291_),
    .A1(_02292_),
    .S(net809),
    .X(_02293_));
 sky130_fd_sc_hd__mux4_1 _07263_ (.A0(\reg_module.gprf[112] ),
    .A1(\reg_module.gprf[80] ),
    .A2(\reg_module.gprf[48] ),
    .A3(\reg_module.gprf[16] ),
    .S0(net935),
    .S1(net899),
    .X(_02294_));
 sky130_fd_sc_hd__mux4_1 _07264_ (.A0(\reg_module.gprf[240] ),
    .A1(\reg_module.gprf[208] ),
    .A2(\reg_module.gprf[176] ),
    .A3(\reg_module.gprf[144] ),
    .S0(net935),
    .S1(net899),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _07265_ (.A0(_02294_),
    .A1(_02295_),
    .S(net809),
    .X(_02296_));
 sky130_fd_sc_hd__a21o_1 _07266_ (.A1(net855),
    .A2(_02296_),
    .B1(net786),
    .X(_02297_));
 sky130_fd_sc_hd__a21o_1 _07267_ (.A1(net794),
    .A2(_02293_),
    .B1(_02297_),
    .X(_02298_));
 sky130_fd_sc_hd__a21o_1 _07268_ (.A1(\rWrDataWB[16] ),
    .A2(net580),
    .B1(net614),
    .X(_02299_));
 sky130_fd_sc_hd__a31o_1 _07269_ (.A1(net586),
    .A2(_02290_),
    .A3(_02298_),
    .B1(_02299_),
    .X(_02300_));
 sky130_fd_sc_hd__and2_1 _07270_ (.A(_02282_),
    .B(_02300_),
    .X(net110));
 sky130_fd_sc_hd__mux4_1 _07271_ (.A0(\reg_module.gprf[881] ),
    .A1(\reg_module.gprf[849] ),
    .A2(\reg_module.gprf[817] ),
    .A3(\reg_module.gprf[785] ),
    .S0(net920),
    .S1(net884),
    .X(_02301_));
 sky130_fd_sc_hd__or2_1 _07272_ (.A(net804),
    .B(_02301_),
    .X(_02302_));
 sky130_fd_sc_hd__mux4_1 _07273_ (.A0(\reg_module.gprf[1009] ),
    .A1(\reg_module.gprf[977] ),
    .A2(\reg_module.gprf[945] ),
    .A3(\reg_module.gprf[913] ),
    .S0(net920),
    .S1(net884),
    .X(_02303_));
 sky130_fd_sc_hd__o21a_1 _07274_ (.A1(net862),
    .A2(_02303_),
    .B1(net791),
    .X(_02304_));
 sky130_fd_sc_hd__mux4_1 _07275_ (.A0(\reg_module.gprf[625] ),
    .A1(\reg_module.gprf[593] ),
    .A2(\reg_module.gprf[561] ),
    .A3(\reg_module.gprf[529] ),
    .S0(net920),
    .S1(net884),
    .X(_02305_));
 sky130_fd_sc_hd__mux4_1 _07276_ (.A0(\reg_module.gprf[753] ),
    .A1(\reg_module.gprf[721] ),
    .A2(\reg_module.gprf[689] ),
    .A3(\reg_module.gprf[657] ),
    .S0(net920),
    .S1(net884),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _07277_ (.A0(_02305_),
    .A1(_02306_),
    .S(net805),
    .X(_02307_));
 sky130_fd_sc_hd__a221o_1 _07278_ (.A1(_02302_),
    .A2(_02304_),
    .B1(_02307_),
    .B2(net853),
    .C1(net941),
    .X(_02308_));
 sky130_fd_sc_hd__mux4_1 _07279_ (.A0(\reg_module.gprf[369] ),
    .A1(\reg_module.gprf[337] ),
    .A2(\reg_module.gprf[305] ),
    .A3(\reg_module.gprf[273] ),
    .S0(net919),
    .S1(net883),
    .X(_02309_));
 sky130_fd_sc_hd__mux4_1 _07280_ (.A0(\reg_module.gprf[497] ),
    .A1(\reg_module.gprf[465] ),
    .A2(\reg_module.gprf[433] ),
    .A3(\reg_module.gprf[401] ),
    .S0(net919),
    .S1(net883),
    .X(_02310_));
 sky130_fd_sc_hd__mux2_1 _07281_ (.A0(_02309_),
    .A1(_02310_),
    .S(net804),
    .X(_02311_));
 sky130_fd_sc_hd__mux4_1 _07282_ (.A0(\reg_module.gprf[113] ),
    .A1(\reg_module.gprf[81] ),
    .A2(\reg_module.gprf[49] ),
    .A3(\reg_module.gprf[17] ),
    .S0(net919),
    .S1(net883),
    .X(_02312_));
 sky130_fd_sc_hd__or2_1 _07283_ (.A(net804),
    .B(_02312_),
    .X(_02313_));
 sky130_fd_sc_hd__mux4_1 _07284_ (.A0(\reg_module.gprf[241] ),
    .A1(\reg_module.gprf[209] ),
    .A2(\reg_module.gprf[177] ),
    .A3(\reg_module.gprf[145] ),
    .S0(net919),
    .S1(net883),
    .X(_02314_));
 sky130_fd_sc_hd__o211a_1 _07285_ (.A1(net862),
    .A2(_02314_),
    .B1(_02313_),
    .C1(net853),
    .X(_02315_));
 sky130_fd_sc_hd__a21o_1 _07286_ (.A1(net791),
    .A2(_02311_),
    .B1(net785),
    .X(_02316_));
 sky130_fd_sc_hd__o211a_1 _07287_ (.A1(_02315_),
    .A2(_02316_),
    .B1(net585),
    .C1(_02308_),
    .X(_02317_));
 sky130_fd_sc_hd__a21o_1 _07288_ (.A1(\rWrDataWB[17] ),
    .A2(net579),
    .B1(net613),
    .X(_02318_));
 sky130_fd_sc_hd__o22a_1 _07289_ (.A1(\rWrData[17] ),
    .A2(net605),
    .B1(_02317_),
    .B2(_02318_),
    .X(net111));
 sky130_fd_sc_hd__mux4_1 _07290_ (.A0(\reg_module.gprf[882] ),
    .A1(\reg_module.gprf[850] ),
    .A2(\reg_module.gprf[818] ),
    .A3(\reg_module.gprf[786] ),
    .S0(net919),
    .S1(net883),
    .X(_02319_));
 sky130_fd_sc_hd__mux4_1 _07291_ (.A0(\reg_module.gprf[1010] ),
    .A1(\reg_module.gprf[978] ),
    .A2(\reg_module.gprf[946] ),
    .A3(\reg_module.gprf[914] ),
    .S0(net909),
    .S1(net872),
    .X(_02320_));
 sky130_fd_sc_hd__or2_1 _07292_ (.A(net859),
    .B(_02320_),
    .X(_02321_));
 sky130_fd_sc_hd__o21a_1 _07293_ (.A1(net799),
    .A2(_02319_),
    .B1(net791),
    .X(_02322_));
 sky130_fd_sc_hd__mux4_1 _07294_ (.A0(\reg_module.gprf[626] ),
    .A1(\reg_module.gprf[594] ),
    .A2(\reg_module.gprf[562] ),
    .A3(\reg_module.gprf[530] ),
    .S0(net919),
    .S1(net883),
    .X(_02323_));
 sky130_fd_sc_hd__mux4_1 _07295_ (.A0(\reg_module.gprf[754] ),
    .A1(\reg_module.gprf[722] ),
    .A2(\reg_module.gprf[690] ),
    .A3(\reg_module.gprf[658] ),
    .S0(net909),
    .S1(net872),
    .X(_02324_));
 sky130_fd_sc_hd__mux2_1 _07296_ (.A0(_02323_),
    .A1(_02324_),
    .S(net799),
    .X(_02325_));
 sky130_fd_sc_hd__a221o_1 _07297_ (.A1(_02321_),
    .A2(_02322_),
    .B1(_02325_),
    .B2(net853),
    .C1(net941),
    .X(_02326_));
 sky130_fd_sc_hd__mux4_1 _07298_ (.A0(\reg_module.gprf[370] ),
    .A1(\reg_module.gprf[338] ),
    .A2(\reg_module.gprf[306] ),
    .A3(\reg_module.gprf[274] ),
    .S0(net919),
    .S1(net883),
    .X(_02327_));
 sky130_fd_sc_hd__or2_1 _07299_ (.A(net804),
    .B(_02327_),
    .X(_02328_));
 sky130_fd_sc_hd__mux4_1 _07300_ (.A0(\reg_module.gprf[498] ),
    .A1(\reg_module.gprf[466] ),
    .A2(\reg_module.gprf[434] ),
    .A3(\reg_module.gprf[402] ),
    .S0(net919),
    .S1(net883),
    .X(_02329_));
 sky130_fd_sc_hd__o211a_1 _07301_ (.A1(net862),
    .A2(_02329_),
    .B1(_02328_),
    .C1(net791),
    .X(_02330_));
 sky130_fd_sc_hd__mux4_1 _07302_ (.A0(\reg_module.gprf[114] ),
    .A1(\reg_module.gprf[82] ),
    .A2(\reg_module.gprf[50] ),
    .A3(\reg_module.gprf[18] ),
    .S0(net909),
    .S1(net872),
    .X(_02331_));
 sky130_fd_sc_hd__mux4_1 _07303_ (.A0(\reg_module.gprf[242] ),
    .A1(\reg_module.gprf[210] ),
    .A2(\reg_module.gprf[178] ),
    .A3(\reg_module.gprf[146] ),
    .S0(net919),
    .S1(net883),
    .X(_02332_));
 sky130_fd_sc_hd__mux2_1 _07304_ (.A0(_02331_),
    .A1(_02332_),
    .S(net804),
    .X(_02333_));
 sky130_fd_sc_hd__a21o_1 _07305_ (.A1(net853),
    .A2(_02333_),
    .B1(net785),
    .X(_02334_));
 sky130_fd_sc_hd__o211ai_1 _07306_ (.A1(_02330_),
    .A2(_02334_),
    .B1(net585),
    .C1(_02326_),
    .Y(_02335_));
 sky130_fd_sc_hd__a21oi_1 _07307_ (.A1(\rWrDataWB[18] ),
    .A2(net579),
    .B1(net613),
    .Y(_02336_));
 sky130_fd_sc_hd__o2bb2a_1 _07308_ (.A1_N(_02336_),
    .A2_N(_02335_),
    .B1(net605),
    .B2(\rWrData[18] ),
    .X(net112));
 sky130_fd_sc_hd__mux4_1 _07309_ (.A0(\reg_module.gprf[883] ),
    .A1(\reg_module.gprf[851] ),
    .A2(\reg_module.gprf[819] ),
    .A3(\reg_module.gprf[787] ),
    .S0(net922),
    .S1(net886),
    .X(_02337_));
 sky130_fd_sc_hd__or2_1 _07310_ (.A(net804),
    .B(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__mux4_1 _07311_ (.A0(\reg_module.gprf[1011] ),
    .A1(\reg_module.gprf[979] ),
    .A2(\reg_module.gprf[947] ),
    .A3(\reg_module.gprf[915] ),
    .S0(net922),
    .S1(net886),
    .X(_02339_));
 sky130_fd_sc_hd__o21a_1 _07312_ (.A1(net862),
    .A2(_02339_),
    .B1(net791),
    .X(_02340_));
 sky130_fd_sc_hd__mux4_1 _07313_ (.A0(\reg_module.gprf[627] ),
    .A1(\reg_module.gprf[595] ),
    .A2(\reg_module.gprf[563] ),
    .A3(\reg_module.gprf[531] ),
    .S0(net919),
    .S1(net883),
    .X(_02341_));
 sky130_fd_sc_hd__mux4_1 _07314_ (.A0(\reg_module.gprf[755] ),
    .A1(\reg_module.gprf[723] ),
    .A2(\reg_module.gprf[691] ),
    .A3(\reg_module.gprf[659] ),
    .S0(net920),
    .S1(net884),
    .X(_02342_));
 sky130_fd_sc_hd__mux2_1 _07315_ (.A0(_02341_),
    .A1(_02342_),
    .S(net804),
    .X(_02343_));
 sky130_fd_sc_hd__a221o_1 _07316_ (.A1(_02338_),
    .A2(_02340_),
    .B1(_02343_),
    .B2(net853),
    .C1(net941),
    .X(_02344_));
 sky130_fd_sc_hd__mux4_1 _07317_ (.A0(\reg_module.gprf[371] ),
    .A1(\reg_module.gprf[339] ),
    .A2(\reg_module.gprf[307] ),
    .A3(\reg_module.gprf[275] ),
    .S0(net922),
    .S1(net886),
    .X(_02345_));
 sky130_fd_sc_hd__or2_1 _07318_ (.A(net804),
    .B(_02345_),
    .X(_02346_));
 sky130_fd_sc_hd__mux4_1 _07319_ (.A0(\reg_module.gprf[499] ),
    .A1(\reg_module.gprf[467] ),
    .A2(\reg_module.gprf[435] ),
    .A3(\reg_module.gprf[403] ),
    .S0(net922),
    .S1(net886),
    .X(_02347_));
 sky130_fd_sc_hd__o211a_1 _07320_ (.A1(net862),
    .A2(_02347_),
    .B1(_02346_),
    .C1(net791),
    .X(_02348_));
 sky130_fd_sc_hd__mux4_1 _07321_ (.A0(\reg_module.gprf[115] ),
    .A1(\reg_module.gprf[83] ),
    .A2(\reg_module.gprf[51] ),
    .A3(\reg_module.gprf[19] ),
    .S0(net920),
    .S1(net884),
    .X(_02349_));
 sky130_fd_sc_hd__mux4_1 _07322_ (.A0(\reg_module.gprf[243] ),
    .A1(\reg_module.gprf[211] ),
    .A2(\reg_module.gprf[179] ),
    .A3(\reg_module.gprf[147] ),
    .S0(net921),
    .S1(net885),
    .X(_02350_));
 sky130_fd_sc_hd__mux2_1 _07323_ (.A0(_02349_),
    .A1(_02350_),
    .S(net804),
    .X(_02351_));
 sky130_fd_sc_hd__a21o_1 _07324_ (.A1(net853),
    .A2(_02351_),
    .B1(net785),
    .X(_02352_));
 sky130_fd_sc_hd__o211ai_1 _07325_ (.A1(_02348_),
    .A2(_02352_),
    .B1(net585),
    .C1(_02344_),
    .Y(_02353_));
 sky130_fd_sc_hd__a21oi_1 _07326_ (.A1(\rWrDataWB[19] ),
    .A2(net579),
    .B1(net613),
    .Y(_02354_));
 sky130_fd_sc_hd__o2bb2a_1 _07327_ (.A1_N(_02354_),
    .A2_N(_02353_),
    .B1(net605),
    .B2(\rWrData[19] ),
    .X(net113));
 sky130_fd_sc_hd__mux4_1 _07328_ (.A0(\reg_module.gprf[884] ),
    .A1(\reg_module.gprf[852] ),
    .A2(\reg_module.gprf[820] ),
    .A3(\reg_module.gprf[788] ),
    .S0(net911),
    .S1(net874),
    .X(_02355_));
 sky130_fd_sc_hd__or2_1 _07329_ (.A(net800),
    .B(_02355_),
    .X(_02356_));
 sky130_fd_sc_hd__mux4_1 _07330_ (.A0(\reg_module.gprf[1012] ),
    .A1(\reg_module.gprf[980] ),
    .A2(\reg_module.gprf[948] ),
    .A3(\reg_module.gprf[916] ),
    .S0(net911),
    .S1(net874),
    .X(_02357_));
 sky130_fd_sc_hd__o21a_1 _07331_ (.A1(net859),
    .A2(_02357_),
    .B1(net789),
    .X(_02358_));
 sky130_fd_sc_hd__mux4_1 _07332_ (.A0(\reg_module.gprf[628] ),
    .A1(\reg_module.gprf[596] ),
    .A2(\reg_module.gprf[564] ),
    .A3(\reg_module.gprf[532] ),
    .S0(net911),
    .S1(net874),
    .X(_02359_));
 sky130_fd_sc_hd__mux4_1 _07333_ (.A0(\reg_module.gprf[756] ),
    .A1(\reg_module.gprf[724] ),
    .A2(\reg_module.gprf[692] ),
    .A3(\reg_module.gprf[660] ),
    .S0(net913),
    .S1(net876),
    .X(_02360_));
 sky130_fd_sc_hd__mux2_1 _07334_ (.A0(_02359_),
    .A1(_02360_),
    .S(net800),
    .X(_02361_));
 sky130_fd_sc_hd__a221o_1 _07335_ (.A1(_02356_),
    .A2(_02358_),
    .B1(_02361_),
    .B2(net849),
    .C1(net939),
    .X(_02362_));
 sky130_fd_sc_hd__mux4_1 _07336_ (.A0(\reg_module.gprf[372] ),
    .A1(\reg_module.gprf[340] ),
    .A2(\reg_module.gprf[308] ),
    .A3(\reg_module.gprf[276] ),
    .S0(net911),
    .S1(net874),
    .X(_02363_));
 sky130_fd_sc_hd__mux4_1 _07337_ (.A0(\reg_module.gprf[500] ),
    .A1(\reg_module.gprf[468] ),
    .A2(\reg_module.gprf[436] ),
    .A3(\reg_module.gprf[404] ),
    .S0(net923),
    .S1(net887),
    .X(_02364_));
 sky130_fd_sc_hd__mux2_1 _07338_ (.A0(_02363_),
    .A1(_02364_),
    .S(net800),
    .X(_02365_));
 sky130_fd_sc_hd__mux4_1 _07339_ (.A0(\reg_module.gprf[116] ),
    .A1(\reg_module.gprf[84] ),
    .A2(\reg_module.gprf[52] ),
    .A3(\reg_module.gprf[20] ),
    .S0(net911),
    .S1(net874),
    .X(_02366_));
 sky130_fd_sc_hd__or2_1 _07340_ (.A(net800),
    .B(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__mux4_1 _07341_ (.A0(\reg_module.gprf[244] ),
    .A1(\reg_module.gprf[212] ),
    .A2(\reg_module.gprf[180] ),
    .A3(\reg_module.gprf[148] ),
    .S0(net911),
    .S1(net874),
    .X(_02368_));
 sky130_fd_sc_hd__o211a_1 _07342_ (.A1(net859),
    .A2(_02368_),
    .B1(_02367_),
    .C1(net850),
    .X(_02369_));
 sky130_fd_sc_hd__a21o_1 _07343_ (.A1(net789),
    .A2(_02365_),
    .B1(net783),
    .X(_02370_));
 sky130_fd_sc_hd__o211a_1 _07344_ (.A1(_02369_),
    .A2(_02370_),
    .B1(net583),
    .C1(_02362_),
    .X(_02371_));
 sky130_fd_sc_hd__a21o_1 _07345_ (.A1(\rWrDataWB[20] ),
    .A2(net579),
    .B1(net613),
    .X(_02372_));
 sky130_fd_sc_hd__o22a_1 _07346_ (.A1(\rWrData[20] ),
    .A2(net605),
    .B1(_02371_),
    .B2(_02372_),
    .X(net115));
 sky130_fd_sc_hd__mux4_1 _07347_ (.A0(\reg_module.gprf[885] ),
    .A1(\reg_module.gprf[853] ),
    .A2(\reg_module.gprf[821] ),
    .A3(\reg_module.gprf[789] ),
    .S0(net933),
    .S1(net898),
    .X(_02373_));
 sky130_fd_sc_hd__or2_1 _07348_ (.A(net809),
    .B(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__mux4_1 _07349_ (.A0(\reg_module.gprf[1013] ),
    .A1(\reg_module.gprf[981] ),
    .A2(\reg_module.gprf[949] ),
    .A3(\reg_module.gprf[917] ),
    .S0(net933),
    .S1(net898),
    .X(_02375_));
 sky130_fd_sc_hd__o21a_1 _07350_ (.A1(net864),
    .A2(_02375_),
    .B1(net793),
    .X(_02376_));
 sky130_fd_sc_hd__mux4_1 _07351_ (.A0(\reg_module.gprf[629] ),
    .A1(\reg_module.gprf[597] ),
    .A2(\reg_module.gprf[565] ),
    .A3(\reg_module.gprf[533] ),
    .S0(net933),
    .S1(net898),
    .X(_02377_));
 sky130_fd_sc_hd__mux4_1 _07352_ (.A0(\reg_module.gprf[757] ),
    .A1(\reg_module.gprf[725] ),
    .A2(\reg_module.gprf[693] ),
    .A3(\reg_module.gprf[661] ),
    .S0(net934),
    .S1(net897),
    .X(_02378_));
 sky130_fd_sc_hd__mux2_1 _07353_ (.A0(_02377_),
    .A1(_02378_),
    .S(net809),
    .X(_02379_));
 sky130_fd_sc_hd__a221o_1 _07354_ (.A1(_02374_),
    .A2(_02376_),
    .B1(_02379_),
    .B2(net855),
    .C1(net942),
    .X(_02380_));
 sky130_fd_sc_hd__mux4_1 _07355_ (.A0(\reg_module.gprf[373] ),
    .A1(\reg_module.gprf[341] ),
    .A2(\reg_module.gprf[309] ),
    .A3(\reg_module.gprf[277] ),
    .S0(net934),
    .S1(net897),
    .X(_02381_));
 sky130_fd_sc_hd__or2_1 _07356_ (.A(net809),
    .B(_02381_),
    .X(_02382_));
 sky130_fd_sc_hd__mux4_1 _07357_ (.A0(\reg_module.gprf[501] ),
    .A1(\reg_module.gprf[469] ),
    .A2(\reg_module.gprf[437] ),
    .A3(\reg_module.gprf[405] ),
    .S0(net934),
    .S1(net898),
    .X(_02383_));
 sky130_fd_sc_hd__o211a_1 _07358_ (.A1(net864),
    .A2(_02383_),
    .B1(_02382_),
    .C1(net793),
    .X(_02384_));
 sky130_fd_sc_hd__mux4_1 _07359_ (.A0(\reg_module.gprf[117] ),
    .A1(\reg_module.gprf[85] ),
    .A2(\reg_module.gprf[53] ),
    .A3(\reg_module.gprf[21] ),
    .S0(net934),
    .S1(net898),
    .X(_02385_));
 sky130_fd_sc_hd__mux4_1 _07360_ (.A0(\reg_module.gprf[245] ),
    .A1(\reg_module.gprf[213] ),
    .A2(\reg_module.gprf[181] ),
    .A3(\reg_module.gprf[149] ),
    .S0(net933),
    .S1(net897),
    .X(_02386_));
 sky130_fd_sc_hd__mux2_1 _07361_ (.A0(_02385_),
    .A1(_02386_),
    .S(net809),
    .X(_02387_));
 sky130_fd_sc_hd__a21o_1 _07362_ (.A1(net855),
    .A2(_02387_),
    .B1(net786),
    .X(_02388_));
 sky130_fd_sc_hd__o211ai_2 _07363_ (.A1(_02384_),
    .A2(_02388_),
    .B1(net586),
    .C1(_02380_),
    .Y(_02389_));
 sky130_fd_sc_hd__a21oi_1 _07364_ (.A1(\rWrDataWB[21] ),
    .A2(net580),
    .B1(net615),
    .Y(_02390_));
 sky130_fd_sc_hd__o2bb2a_1 _07365_ (.A1_N(_02390_),
    .A2_N(_02389_),
    .B1(net607),
    .B2(\rWrData[21] ),
    .X(net116));
 sky130_fd_sc_hd__mux4_1 _07366_ (.A0(\reg_module.gprf[886] ),
    .A1(\reg_module.gprf[854] ),
    .A2(\reg_module.gprf[822] ),
    .A3(\reg_module.gprf[790] ),
    .S0(net932),
    .S1(net895),
    .X(_02391_));
 sky130_fd_sc_hd__mux4_1 _07367_ (.A0(\reg_module.gprf[1014] ),
    .A1(\reg_module.gprf[982] ),
    .A2(\reg_module.gprf[950] ),
    .A3(\reg_module.gprf[918] ),
    .S0(net931),
    .S1(net895),
    .X(_02392_));
 sky130_fd_sc_hd__or2_1 _07368_ (.A(\brancher.imm21_j[2] ),
    .B(_02392_),
    .X(_02393_));
 sky130_fd_sc_hd__o21a_1 _07369_ (.A1(net810),
    .A2(_02391_),
    .B1(net794),
    .X(_02394_));
 sky130_fd_sc_hd__mux4_1 _07370_ (.A0(\reg_module.gprf[630] ),
    .A1(\reg_module.gprf[598] ),
    .A2(\reg_module.gprf[566] ),
    .A3(\reg_module.gprf[534] ),
    .S0(net931),
    .S1(net896),
    .X(_02395_));
 sky130_fd_sc_hd__mux4_1 _07371_ (.A0(\reg_module.gprf[758] ),
    .A1(\reg_module.gprf[726] ),
    .A2(\reg_module.gprf[694] ),
    .A3(\reg_module.gprf[662] ),
    .S0(net932),
    .S1(net895),
    .X(_02396_));
 sky130_fd_sc_hd__mux2_1 _07372_ (.A0(_02395_),
    .A1(_02396_),
    .S(net810),
    .X(_02397_));
 sky130_fd_sc_hd__a221o_1 _07373_ (.A1(_02393_),
    .A2(_02394_),
    .B1(_02397_),
    .B2(net856),
    .C1(net942),
    .X(_02398_));
 sky130_fd_sc_hd__mux4_1 _07374_ (.A0(\reg_module.gprf[374] ),
    .A1(\reg_module.gprf[342] ),
    .A2(\reg_module.gprf[310] ),
    .A3(\reg_module.gprf[278] ),
    .S0(net932),
    .S1(net896),
    .X(_02399_));
 sky130_fd_sc_hd__mux4_1 _07375_ (.A0(\reg_module.gprf[502] ),
    .A1(\reg_module.gprf[470] ),
    .A2(\reg_module.gprf[438] ),
    .A3(\reg_module.gprf[406] ),
    .S0(net931),
    .S1(net896),
    .X(_02400_));
 sky130_fd_sc_hd__mux2_1 _07376_ (.A0(_02399_),
    .A1(_02400_),
    .S(net810),
    .X(_02401_));
 sky130_fd_sc_hd__mux4_1 _07377_ (.A0(\reg_module.gprf[118] ),
    .A1(\reg_module.gprf[86] ),
    .A2(\reg_module.gprf[54] ),
    .A3(\reg_module.gprf[22] ),
    .S0(net932),
    .S1(net896),
    .X(_02402_));
 sky130_fd_sc_hd__mux4_1 _07378_ (.A0(\reg_module.gprf[246] ),
    .A1(\reg_module.gprf[214] ),
    .A2(\reg_module.gprf[182] ),
    .A3(\reg_module.gprf[150] ),
    .S0(net932),
    .S1(net895),
    .X(_02403_));
 sky130_fd_sc_hd__or2_1 _07379_ (.A(net864),
    .B(_02403_),
    .X(_02404_));
 sky130_fd_sc_hd__o211a_1 _07380_ (.A1(net810),
    .A2(_02402_),
    .B1(_02404_),
    .C1(net855),
    .X(_02405_));
 sky130_fd_sc_hd__a21o_1 _07381_ (.A1(net793),
    .A2(_02401_),
    .B1(net786),
    .X(_02406_));
 sky130_fd_sc_hd__o211a_1 _07382_ (.A1(_02405_),
    .A2(_02406_),
    .B1(net586),
    .C1(_02398_),
    .X(_02407_));
 sky130_fd_sc_hd__a21o_1 _07383_ (.A1(\rWrDataWB[22] ),
    .A2(net580),
    .B1(net614),
    .X(_02408_));
 sky130_fd_sc_hd__o22a_1 _07384_ (.A1(\rWrData[22] ),
    .A2(net607),
    .B1(_02407_),
    .B2(_02408_),
    .X(net117));
 sky130_fd_sc_hd__mux4_1 _07385_ (.A0(\reg_module.gprf[887] ),
    .A1(\reg_module.gprf[855] ),
    .A2(\reg_module.gprf[823] ),
    .A3(\reg_module.gprf[791] ),
    .S0(net925),
    .S1(net889),
    .X(_02409_));
 sky130_fd_sc_hd__or2_1 _07386_ (.A(net807),
    .B(_02409_),
    .X(_02410_));
 sky130_fd_sc_hd__mux4_1 _07387_ (.A0(\reg_module.gprf[1015] ),
    .A1(\reg_module.gprf[983] ),
    .A2(\reg_module.gprf[951] ),
    .A3(\reg_module.gprf[919] ),
    .S0(net925),
    .S1(net889),
    .X(_02411_));
 sky130_fd_sc_hd__o21a_1 _07388_ (.A1(net863),
    .A2(_02411_),
    .B1(net792),
    .X(_02412_));
 sky130_fd_sc_hd__mux4_1 _07389_ (.A0(\reg_module.gprf[631] ),
    .A1(\reg_module.gprf[599] ),
    .A2(\reg_module.gprf[567] ),
    .A3(\reg_module.gprf[535] ),
    .S0(net925),
    .S1(net889),
    .X(_02413_));
 sky130_fd_sc_hd__mux4_1 _07390_ (.A0(\reg_module.gprf[759] ),
    .A1(\reg_module.gprf[727] ),
    .A2(\reg_module.gprf[695] ),
    .A3(\reg_module.gprf[663] ),
    .S0(net925),
    .S1(net889),
    .X(_02414_));
 sky130_fd_sc_hd__mux2_1 _07391_ (.A0(_02413_),
    .A1(_02414_),
    .S(net807),
    .X(_02415_));
 sky130_fd_sc_hd__a221o_1 _07392_ (.A1(_02410_),
    .A2(_02412_),
    .B1(_02415_),
    .B2(net854),
    .C1(net941),
    .X(_02416_));
 sky130_fd_sc_hd__mux4_1 _07393_ (.A0(\reg_module.gprf[375] ),
    .A1(\reg_module.gprf[343] ),
    .A2(\reg_module.gprf[311] ),
    .A3(\reg_module.gprf[279] ),
    .S0(net924),
    .S1(net888),
    .X(_02417_));
 sky130_fd_sc_hd__mux4_1 _07394_ (.A0(\reg_module.gprf[503] ),
    .A1(\reg_module.gprf[471] ),
    .A2(\reg_module.gprf[439] ),
    .A3(\reg_module.gprf[407] ),
    .S0(net925),
    .S1(net889),
    .X(_02418_));
 sky130_fd_sc_hd__mux2_1 _07395_ (.A0(_02417_),
    .A1(_02418_),
    .S(net807),
    .X(_02419_));
 sky130_fd_sc_hd__mux4_1 _07396_ (.A0(\reg_module.gprf[119] ),
    .A1(\reg_module.gprf[87] ),
    .A2(\reg_module.gprf[55] ),
    .A3(\reg_module.gprf[23] ),
    .S0(net925),
    .S1(net889),
    .X(_02420_));
 sky130_fd_sc_hd__mux4_1 _07397_ (.A0(\reg_module.gprf[247] ),
    .A1(\reg_module.gprf[215] ),
    .A2(\reg_module.gprf[183] ),
    .A3(\reg_module.gprf[151] ),
    .S0(net925),
    .S1(net889),
    .X(_02421_));
 sky130_fd_sc_hd__or2_1 _07398_ (.A(net863),
    .B(_02421_),
    .X(_02422_));
 sky130_fd_sc_hd__o211a_1 _07399_ (.A1(net807),
    .A2(_02420_),
    .B1(_02422_),
    .C1(net854),
    .X(_02423_));
 sky130_fd_sc_hd__a21o_1 _07400_ (.A1(net792),
    .A2(_02419_),
    .B1(net785),
    .X(_02424_));
 sky130_fd_sc_hd__o211a_1 _07401_ (.A1(_02423_),
    .A2(_02424_),
    .B1(net585),
    .C1(_02416_),
    .X(_02425_));
 sky130_fd_sc_hd__a21o_1 _07402_ (.A1(\rWrDataWB[23] ),
    .A2(net578),
    .B1(net612),
    .X(_02426_));
 sky130_fd_sc_hd__o22a_1 _07403_ (.A1(\rWrData[23] ),
    .A2(net606),
    .B1(_02425_),
    .B2(_02426_),
    .X(net118));
 sky130_fd_sc_hd__or2_1 _07404_ (.A(\rWrData[24] ),
    .B(net606),
    .X(_02427_));
 sky130_fd_sc_hd__mux4_1 _07405_ (.A0(\reg_module.gprf[760] ),
    .A1(\reg_module.gprf[728] ),
    .A2(\reg_module.gprf[696] ),
    .A3(\reg_module.gprf[664] ),
    .S0(net926),
    .S1(net890),
    .X(_02428_));
 sky130_fd_sc_hd__mux4_1 _07406_ (.A0(\reg_module.gprf[632] ),
    .A1(\reg_module.gprf[600] ),
    .A2(\reg_module.gprf[568] ),
    .A3(\reg_module.gprf[536] ),
    .S0(net926),
    .S1(net890),
    .X(_02429_));
 sky130_fd_sc_hd__mux2_1 _07407_ (.A0(_02428_),
    .A1(_02429_),
    .S(net863),
    .X(_02430_));
 sky130_fd_sc_hd__mux4_1 _07408_ (.A0(\reg_module.gprf[888] ),
    .A1(\reg_module.gprf[856] ),
    .A2(\reg_module.gprf[824] ),
    .A3(\reg_module.gprf[792] ),
    .S0(net928),
    .S1(net892),
    .X(_02431_));
 sky130_fd_sc_hd__mux4_1 _07409_ (.A0(\reg_module.gprf[1016] ),
    .A1(\reg_module.gprf[984] ),
    .A2(\reg_module.gprf[952] ),
    .A3(\reg_module.gprf[920] ),
    .S0(net928),
    .S1(net892),
    .X(_02432_));
 sky130_fd_sc_hd__mux2_1 _07410_ (.A0(_02431_),
    .A1(_02432_),
    .S(net808),
    .X(_02433_));
 sky130_fd_sc_hd__a21o_1 _07411_ (.A1(net792),
    .A2(_02433_),
    .B1(net941),
    .X(_02434_));
 sky130_fd_sc_hd__a21o_1 _07412_ (.A1(net854),
    .A2(_02430_),
    .B1(_02434_),
    .X(_02435_));
 sky130_fd_sc_hd__mux4_1 _07413_ (.A0(\reg_module.gprf[376] ),
    .A1(\reg_module.gprf[344] ),
    .A2(\reg_module.gprf[312] ),
    .A3(\reg_module.gprf[280] ),
    .S0(net926),
    .S1(net890),
    .X(_02436_));
 sky130_fd_sc_hd__mux4_1 _07414_ (.A0(\reg_module.gprf[504] ),
    .A1(\reg_module.gprf[472] ),
    .A2(\reg_module.gprf[440] ),
    .A3(\reg_module.gprf[408] ),
    .S0(net928),
    .S1(net892),
    .X(_02437_));
 sky130_fd_sc_hd__mux2_1 _07415_ (.A0(_02436_),
    .A1(_02437_),
    .S(net808),
    .X(_02438_));
 sky130_fd_sc_hd__mux4_1 _07416_ (.A0(\reg_module.gprf[120] ),
    .A1(\reg_module.gprf[88] ),
    .A2(\reg_module.gprf[56] ),
    .A3(\reg_module.gprf[24] ),
    .S0(net928),
    .S1(net892),
    .X(_02439_));
 sky130_fd_sc_hd__mux4_1 _07417_ (.A0(\reg_module.gprf[248] ),
    .A1(\reg_module.gprf[216] ),
    .A2(\reg_module.gprf[184] ),
    .A3(\reg_module.gprf[152] ),
    .S0(net926),
    .S1(net890),
    .X(_02440_));
 sky130_fd_sc_hd__mux2_1 _07418_ (.A0(_02439_),
    .A1(_02440_),
    .S(net808),
    .X(_02441_));
 sky130_fd_sc_hd__a21o_1 _07419_ (.A1(net854),
    .A2(_02441_),
    .B1(net785),
    .X(_02442_));
 sky130_fd_sc_hd__a21o_1 _07420_ (.A1(net792),
    .A2(_02438_),
    .B1(_02442_),
    .X(_02443_));
 sky130_fd_sc_hd__and2_1 _07421_ (.A(\rWrDataWB[24] ),
    .B(net578),
    .X(_02444_));
 sky130_fd_sc_hd__a31o_1 _07422_ (.A1(net585),
    .A2(_02435_),
    .A3(_02443_),
    .B1(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__o21a_1 _07423_ (.A1(net612),
    .A2(_02445_),
    .B1(_02427_),
    .X(net119));
 sky130_fd_sc_hd__mux4_1 _07424_ (.A0(\reg_module.gprf[889] ),
    .A1(\reg_module.gprf[857] ),
    .A2(\reg_module.gprf[825] ),
    .A3(\reg_module.gprf[793] ),
    .S0(net924),
    .S1(net888),
    .X(_02446_));
 sky130_fd_sc_hd__or2_1 _07425_ (.A(net807),
    .B(_02446_),
    .X(_02447_));
 sky130_fd_sc_hd__mux4_1 _07426_ (.A0(\reg_module.gprf[1017] ),
    .A1(\reg_module.gprf[985] ),
    .A2(\reg_module.gprf[953] ),
    .A3(\reg_module.gprf[921] ),
    .S0(net926),
    .S1(net890),
    .X(_02448_));
 sky130_fd_sc_hd__o21a_1 _07427_ (.A1(net863),
    .A2(_02448_),
    .B1(net792),
    .X(_02449_));
 sky130_fd_sc_hd__mux4_1 _07428_ (.A0(\reg_module.gprf[633] ),
    .A1(\reg_module.gprf[601] ),
    .A2(\reg_module.gprf[569] ),
    .A3(\reg_module.gprf[537] ),
    .S0(net926),
    .S1(net890),
    .X(_02450_));
 sky130_fd_sc_hd__mux4_1 _07429_ (.A0(\reg_module.gprf[761] ),
    .A1(\reg_module.gprf[729] ),
    .A2(\reg_module.gprf[697] ),
    .A3(\reg_module.gprf[665] ),
    .S0(net929),
    .S1(net893),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _07430_ (.A0(_02450_),
    .A1(_02451_),
    .S(net808),
    .X(_02452_));
 sky130_fd_sc_hd__a221o_1 _07431_ (.A1(_02447_),
    .A2(_02449_),
    .B1(_02452_),
    .B2(net854),
    .C1(net942),
    .X(_02453_));
 sky130_fd_sc_hd__mux4_1 _07432_ (.A0(\reg_module.gprf[377] ),
    .A1(\reg_module.gprf[345] ),
    .A2(\reg_module.gprf[313] ),
    .A3(\reg_module.gprf[281] ),
    .S0(net924),
    .S1(net888),
    .X(_02454_));
 sky130_fd_sc_hd__mux4_1 _07433_ (.A0(\reg_module.gprf[505] ),
    .A1(\reg_module.gprf[473] ),
    .A2(\reg_module.gprf[441] ),
    .A3(\reg_module.gprf[409] ),
    .S0(net926),
    .S1(net890),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _07434_ (.A0(_02454_),
    .A1(_02455_),
    .S(net807),
    .X(_02456_));
 sky130_fd_sc_hd__mux4_1 _07435_ (.A0(\reg_module.gprf[121] ),
    .A1(\reg_module.gprf[89] ),
    .A2(\reg_module.gprf[57] ),
    .A3(\reg_module.gprf[25] ),
    .S0(net929),
    .S1(net888),
    .X(_02457_));
 sky130_fd_sc_hd__or2_1 _07436_ (.A(net808),
    .B(_02457_),
    .X(_02458_));
 sky130_fd_sc_hd__mux4_1 _07437_ (.A0(\reg_module.gprf[249] ),
    .A1(\reg_module.gprf[217] ),
    .A2(\reg_module.gprf[185] ),
    .A3(\reg_module.gprf[153] ),
    .S0(net926),
    .S1(net890),
    .X(_02459_));
 sky130_fd_sc_hd__o211a_1 _07438_ (.A1(net863),
    .A2(_02459_),
    .B1(_02458_),
    .C1(net854),
    .X(_02460_));
 sky130_fd_sc_hd__a21o_1 _07439_ (.A1(net792),
    .A2(_02456_),
    .B1(net785),
    .X(_02461_));
 sky130_fd_sc_hd__o211a_1 _07440_ (.A1(_02460_),
    .A2(_02461_),
    .B1(net585),
    .C1(_02453_),
    .X(_02462_));
 sky130_fd_sc_hd__a21o_1 _07441_ (.A1(\rWrDataWB[25] ),
    .A2(net580),
    .B1(net614),
    .X(_02463_));
 sky130_fd_sc_hd__o22a_1 _07442_ (.A1(\rWrData[25] ),
    .A2(net607),
    .B1(_02462_),
    .B2(_02463_),
    .X(net120));
 sky130_fd_sc_hd__mux4_1 _07443_ (.A0(\reg_module.gprf[762] ),
    .A1(\reg_module.gprf[730] ),
    .A2(\reg_module.gprf[698] ),
    .A3(\reg_module.gprf[666] ),
    .S0(net922),
    .S1(net886),
    .X(_02464_));
 sky130_fd_sc_hd__mux4_1 _07444_ (.A0(\reg_module.gprf[634] ),
    .A1(\reg_module.gprf[602] ),
    .A2(\reg_module.gprf[570] ),
    .A3(\reg_module.gprf[538] ),
    .S0(net922),
    .S1(net894),
    .X(_02465_));
 sky130_fd_sc_hd__or2_1 _07445_ (.A(net806),
    .B(_02465_),
    .X(_02466_));
 sky130_fd_sc_hd__o21a_1 _07446_ (.A1(net862),
    .A2(_02464_),
    .B1(net853),
    .X(_02467_));
 sky130_fd_sc_hd__mux4_1 _07447_ (.A0(\reg_module.gprf[890] ),
    .A1(\reg_module.gprf[858] ),
    .A2(\reg_module.gprf[826] ),
    .A3(\reg_module.gprf[794] ),
    .S0(net927),
    .S1(net891),
    .X(_02468_));
 sky130_fd_sc_hd__mux4_1 _07448_ (.A0(\reg_module.gprf[1018] ),
    .A1(\reg_module.gprf[986] ),
    .A2(\reg_module.gprf[954] ),
    .A3(\reg_module.gprf[922] ),
    .S0(net927),
    .S1(net891),
    .X(_02469_));
 sky130_fd_sc_hd__mux2_1 _07449_ (.A0(_02468_),
    .A1(_02469_),
    .S(net811),
    .X(_02470_));
 sky130_fd_sc_hd__a221o_1 _07450_ (.A1(_02466_),
    .A2(_02467_),
    .B1(_02470_),
    .B2(net793),
    .C1(net941),
    .X(_02471_));
 sky130_fd_sc_hd__mux4_1 _07451_ (.A0(\reg_module.gprf[378] ),
    .A1(\reg_module.gprf[346] ),
    .A2(\reg_module.gprf[314] ),
    .A3(\reg_module.gprf[282] ),
    .S0(net930),
    .S1(net894),
    .X(_02472_));
 sky130_fd_sc_hd__mux4_1 _07452_ (.A0(\reg_module.gprf[506] ),
    .A1(\reg_module.gprf[474] ),
    .A2(\reg_module.gprf[442] ),
    .A3(\reg_module.gprf[410] ),
    .S0(net930),
    .S1(net886),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _07453_ (.A0(_02472_),
    .A1(_02473_),
    .S(net806),
    .X(_02474_));
 sky130_fd_sc_hd__mux4_1 _07454_ (.A0(\reg_module.gprf[122] ),
    .A1(\reg_module.gprf[90] ),
    .A2(\reg_module.gprf[58] ),
    .A3(\reg_module.gprf[26] ),
    .S0(net922),
    .S1(net886),
    .X(_02475_));
 sky130_fd_sc_hd__or2_1 _07455_ (.A(net806),
    .B(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__mux4_1 _07456_ (.A0(\reg_module.gprf[250] ),
    .A1(\reg_module.gprf[218] ),
    .A2(\reg_module.gprf[186] ),
    .A3(\reg_module.gprf[154] ),
    .S0(net922),
    .S1(net886),
    .X(_02477_));
 sky130_fd_sc_hd__o211a_1 _07457_ (.A1(net863),
    .A2(_02477_),
    .B1(_02476_),
    .C1(net856),
    .X(_02478_));
 sky130_fd_sc_hd__a21o_1 _07458_ (.A1(net791),
    .A2(_02474_),
    .B1(net785),
    .X(_02479_));
 sky130_fd_sc_hd__o211a_1 _07459_ (.A1(_02478_),
    .A2(_02479_),
    .B1(net585),
    .C1(_02471_),
    .X(_02480_));
 sky130_fd_sc_hd__a21o_1 _07460_ (.A1(\rWrDataWB[26] ),
    .A2(net580),
    .B1(net614),
    .X(_02481_));
 sky130_fd_sc_hd__o22a_2 _07461_ (.A1(\rWrData[26] ),
    .A2(net607),
    .B1(_02480_),
    .B2(_02481_),
    .X(net121));
 sky130_fd_sc_hd__mux4_1 _07462_ (.A0(\reg_module.gprf[891] ),
    .A1(\reg_module.gprf[859] ),
    .A2(\reg_module.gprf[827] ),
    .A3(\reg_module.gprf[795] ),
    .S0(net920),
    .S1(net884),
    .X(_02482_));
 sky130_fd_sc_hd__or2_1 _07463_ (.A(net805),
    .B(_02482_),
    .X(_02483_));
 sky130_fd_sc_hd__mux4_1 _07464_ (.A0(\reg_module.gprf[1019] ),
    .A1(\reg_module.gprf[987] ),
    .A2(\reg_module.gprf[955] ),
    .A3(\reg_module.gprf[923] ),
    .S0(net920),
    .S1(net884),
    .X(_02484_));
 sky130_fd_sc_hd__o21a_1 _07465_ (.A1(net862),
    .A2(_02484_),
    .B1(net791),
    .X(_02485_));
 sky130_fd_sc_hd__mux4_1 _07466_ (.A0(\reg_module.gprf[635] ),
    .A1(\reg_module.gprf[603] ),
    .A2(\reg_module.gprf[571] ),
    .A3(\reg_module.gprf[539] ),
    .S0(net925),
    .S1(net889),
    .X(_02486_));
 sky130_fd_sc_hd__mux4_1 _07467_ (.A0(\reg_module.gprf[763] ),
    .A1(\reg_module.gprf[731] ),
    .A2(\reg_module.gprf[699] ),
    .A3(\reg_module.gprf[667] ),
    .S0(net921),
    .S1(net885),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _07468_ (.A0(_02486_),
    .A1(_02487_),
    .S(net805),
    .X(_02488_));
 sky130_fd_sc_hd__a221o_1 _07469_ (.A1(_02483_),
    .A2(_02485_),
    .B1(_02488_),
    .B2(net853),
    .C1(net941),
    .X(_02489_));
 sky130_fd_sc_hd__mux4_1 _07470_ (.A0(\reg_module.gprf[379] ),
    .A1(\reg_module.gprf[347] ),
    .A2(\reg_module.gprf[315] ),
    .A3(\reg_module.gprf[283] ),
    .S0(net925),
    .S1(net889),
    .X(_02490_));
 sky130_fd_sc_hd__mux4_1 _07471_ (.A0(\reg_module.gprf[507] ),
    .A1(\reg_module.gprf[475] ),
    .A2(\reg_module.gprf[443] ),
    .A3(\reg_module.gprf[411] ),
    .S0(net920),
    .S1(net884),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _07472_ (.A0(_02490_),
    .A1(_02491_),
    .S(net805),
    .X(_02492_));
 sky130_fd_sc_hd__mux4_1 _07473_ (.A0(\reg_module.gprf[123] ),
    .A1(\reg_module.gprf[91] ),
    .A2(\reg_module.gprf[59] ),
    .A3(\reg_module.gprf[27] ),
    .S0(net925),
    .S1(net889),
    .X(_02493_));
 sky130_fd_sc_hd__or2_1 _07474_ (.A(net805),
    .B(_02493_),
    .X(_02494_));
 sky130_fd_sc_hd__mux4_1 _07475_ (.A0(\reg_module.gprf[251] ),
    .A1(\reg_module.gprf[219] ),
    .A2(\reg_module.gprf[187] ),
    .A3(\reg_module.gprf[155] ),
    .S0(net920),
    .S1(net884),
    .X(_02495_));
 sky130_fd_sc_hd__o211a_1 _07476_ (.A1(net862),
    .A2(_02495_),
    .B1(_02494_),
    .C1(net854),
    .X(_02496_));
 sky130_fd_sc_hd__a21o_1 _07477_ (.A1(net792),
    .A2(_02492_),
    .B1(net785),
    .X(_02497_));
 sky130_fd_sc_hd__o211a_1 _07478_ (.A1(_02496_),
    .A2(_02497_),
    .B1(net585),
    .C1(_02489_),
    .X(_02498_));
 sky130_fd_sc_hd__a21o_1 _07479_ (.A1(\rWrDataWB[27] ),
    .A2(net578),
    .B1(net612),
    .X(_02499_));
 sky130_fd_sc_hd__o22a_1 _07480_ (.A1(\rWrData[27] ),
    .A2(net606),
    .B1(_02498_),
    .B2(_02499_),
    .X(net122));
 sky130_fd_sc_hd__or2_1 _07481_ (.A(\rWrData[28] ),
    .B(net606),
    .X(_02500_));
 sky130_fd_sc_hd__mux4_1 _07482_ (.A0(\reg_module.gprf[892] ),
    .A1(\reg_module.gprf[860] ),
    .A2(\reg_module.gprf[828] ),
    .A3(\reg_module.gprf[796] ),
    .S0(net924),
    .S1(net888),
    .X(_02501_));
 sky130_fd_sc_hd__mux4_1 _07483_ (.A0(\reg_module.gprf[1020] ),
    .A1(\reg_module.gprf[988] ),
    .A2(\reg_module.gprf[956] ),
    .A3(\reg_module.gprf[924] ),
    .S0(net924),
    .S1(net888),
    .X(_02502_));
 sky130_fd_sc_hd__mux2_1 _07484_ (.A0(_02501_),
    .A1(_02502_),
    .S(net807),
    .X(_02503_));
 sky130_fd_sc_hd__mux4_1 _07485_ (.A0(\reg_module.gprf[636] ),
    .A1(\reg_module.gprf[604] ),
    .A2(\reg_module.gprf[572] ),
    .A3(\reg_module.gprf[540] ),
    .S0(net924),
    .S1(net893),
    .X(_02504_));
 sky130_fd_sc_hd__mux4_1 _07486_ (.A0(\reg_module.gprf[764] ),
    .A1(\reg_module.gprf[732] ),
    .A2(\reg_module.gprf[700] ),
    .A3(\reg_module.gprf[668] ),
    .S0(net924),
    .S1(net888),
    .X(_02505_));
 sky130_fd_sc_hd__or2_1 _07487_ (.A(net863),
    .B(_02505_),
    .X(_02506_));
 sky130_fd_sc_hd__o211a_1 _07488_ (.A1(net807),
    .A2(_02504_),
    .B1(_02506_),
    .C1(net854),
    .X(_02507_));
 sky130_fd_sc_hd__a211o_1 _07489_ (.A1(net792),
    .A2(_02503_),
    .B1(_02507_),
    .C1(net941),
    .X(_02508_));
 sky130_fd_sc_hd__mux4_1 _07490_ (.A0(\reg_module.gprf[380] ),
    .A1(\reg_module.gprf[348] ),
    .A2(\reg_module.gprf[316] ),
    .A3(\reg_module.gprf[284] ),
    .S0(net924),
    .S1(net888),
    .X(_02509_));
 sky130_fd_sc_hd__mux4_1 _07491_ (.A0(\reg_module.gprf[508] ),
    .A1(\reg_module.gprf[476] ),
    .A2(\reg_module.gprf[444] ),
    .A3(\reg_module.gprf[412] ),
    .S0(net929),
    .S1(net893),
    .X(_02510_));
 sky130_fd_sc_hd__mux2_1 _07492_ (.A0(_02509_),
    .A1(_02510_),
    .S(net807),
    .X(_02511_));
 sky130_fd_sc_hd__mux4_1 _07493_ (.A0(\reg_module.gprf[124] ),
    .A1(\reg_module.gprf[92] ),
    .A2(\reg_module.gprf[60] ),
    .A3(\reg_module.gprf[28] ),
    .S0(net924),
    .S1(net888),
    .X(_02512_));
 sky130_fd_sc_hd__mux4_1 _07494_ (.A0(\reg_module.gprf[252] ),
    .A1(\reg_module.gprf[220] ),
    .A2(\reg_module.gprf[188] ),
    .A3(\reg_module.gprf[156] ),
    .S0(net924),
    .S1(net888),
    .X(_02513_));
 sky130_fd_sc_hd__mux2_1 _07495_ (.A0(_02512_),
    .A1(_02513_),
    .S(net807),
    .X(_02514_));
 sky130_fd_sc_hd__a21o_1 _07496_ (.A1(net854),
    .A2(_02514_),
    .B1(net785),
    .X(_02515_));
 sky130_fd_sc_hd__a21o_1 _07497_ (.A1(net792),
    .A2(_02511_),
    .B1(_02515_),
    .X(_02516_));
 sky130_fd_sc_hd__a21o_1 _07498_ (.A1(\rWrDataWB[28] ),
    .A2(net578),
    .B1(net612),
    .X(_02517_));
 sky130_fd_sc_hd__a31o_1 _07499_ (.A1(net585),
    .A2(_02508_),
    .A3(_02516_),
    .B1(_02517_),
    .X(_02518_));
 sky130_fd_sc_hd__and2_1 _07500_ (.A(_02500_),
    .B(_02518_),
    .X(net123));
 sky130_fd_sc_hd__mux4_1 _07501_ (.A0(\reg_module.gprf[893] ),
    .A1(\reg_module.gprf[861] ),
    .A2(\reg_module.gprf[829] ),
    .A3(\reg_module.gprf[797] ),
    .S0(net927),
    .S1(net891),
    .X(_02519_));
 sky130_fd_sc_hd__or2_1 _07502_ (.A(net808),
    .B(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__mux4_1 _07503_ (.A0(\reg_module.gprf[1021] ),
    .A1(\reg_module.gprf[989] ),
    .A2(\reg_module.gprf[957] ),
    .A3(\reg_module.gprf[925] ),
    .S0(net927),
    .S1(net891),
    .X(_02521_));
 sky130_fd_sc_hd__o21a_1 _07504_ (.A1(net863),
    .A2(_02521_),
    .B1(net793),
    .X(_02522_));
 sky130_fd_sc_hd__mux4_1 _07505_ (.A0(\reg_module.gprf[637] ),
    .A1(\reg_module.gprf[605] ),
    .A2(\reg_module.gprf[573] ),
    .A3(\reg_module.gprf[541] ),
    .S0(net927),
    .S1(net891),
    .X(_02523_));
 sky130_fd_sc_hd__mux4_1 _07506_ (.A0(\reg_module.gprf[765] ),
    .A1(\reg_module.gprf[733] ),
    .A2(\reg_module.gprf[701] ),
    .A3(\reg_module.gprf[669] ),
    .S0(net927),
    .S1(net891),
    .X(_02524_));
 sky130_fd_sc_hd__mux2_1 _07507_ (.A0(_02523_),
    .A1(_02524_),
    .S(net808),
    .X(_02525_));
 sky130_fd_sc_hd__a221o_1 _07508_ (.A1(_02520_),
    .A2(_02522_),
    .B1(_02525_),
    .B2(net854),
    .C1(net941),
    .X(_02526_));
 sky130_fd_sc_hd__mux4_1 _07509_ (.A0(\reg_module.gprf[381] ),
    .A1(\reg_module.gprf[349] ),
    .A2(\reg_module.gprf[317] ),
    .A3(\reg_module.gprf[285] ),
    .S0(net927),
    .S1(net891),
    .X(_02527_));
 sky130_fd_sc_hd__mux4_1 _07510_ (.A0(\reg_module.gprf[509] ),
    .A1(\reg_module.gprf[477] ),
    .A2(\reg_module.gprf[445] ),
    .A3(\reg_module.gprf[413] ),
    .S0(net927),
    .S1(net891),
    .X(_02528_));
 sky130_fd_sc_hd__mux2_1 _07511_ (.A0(_02527_),
    .A1(_02528_),
    .S(net808),
    .X(_02529_));
 sky130_fd_sc_hd__mux4_1 _07512_ (.A0(\reg_module.gprf[125] ),
    .A1(\reg_module.gprf[93] ),
    .A2(\reg_module.gprf[61] ),
    .A3(\reg_module.gprf[29] ),
    .S0(net927),
    .S1(net891),
    .X(_02530_));
 sky130_fd_sc_hd__or2_1 _07513_ (.A(net808),
    .B(_02530_),
    .X(_02531_));
 sky130_fd_sc_hd__mux4_1 _07514_ (.A0(\reg_module.gprf[253] ),
    .A1(\reg_module.gprf[221] ),
    .A2(\reg_module.gprf[189] ),
    .A3(\reg_module.gprf[157] ),
    .S0(net927),
    .S1(net891),
    .X(_02532_));
 sky130_fd_sc_hd__o211a_1 _07515_ (.A1(net863),
    .A2(_02532_),
    .B1(_02531_),
    .C1(net856),
    .X(_02533_));
 sky130_fd_sc_hd__a21o_1 _07516_ (.A1(net792),
    .A2(_02529_),
    .B1(net786),
    .X(_02534_));
 sky130_fd_sc_hd__o211a_1 _07517_ (.A1(_02533_),
    .A2(_02534_),
    .B1(net586),
    .C1(_02526_),
    .X(_02535_));
 sky130_fd_sc_hd__a21o_1 _07518_ (.A1(\rWrDataWB[29] ),
    .A2(net582),
    .B1(net612),
    .X(_02536_));
 sky130_fd_sc_hd__o22a_1 _07519_ (.A1(\rWrData[29] ),
    .A2(net606),
    .B1(_02535_),
    .B2(_02536_),
    .X(net124));
 sky130_fd_sc_hd__mux4_1 _07520_ (.A0(\reg_module.gprf[894] ),
    .A1(\reg_module.gprf[862] ),
    .A2(\reg_module.gprf[830] ),
    .A3(\reg_module.gprf[798] ),
    .S0(net931),
    .S1(net895),
    .X(_02537_));
 sky130_fd_sc_hd__mux4_1 _07521_ (.A0(\reg_module.gprf[1022] ),
    .A1(\reg_module.gprf[990] ),
    .A2(\reg_module.gprf[958] ),
    .A3(\reg_module.gprf[926] ),
    .S0(net931),
    .S1(net895),
    .X(_02538_));
 sky130_fd_sc_hd__or2_1 _07522_ (.A(\brancher.imm21_j[2] ),
    .B(_02538_),
    .X(_02539_));
 sky130_fd_sc_hd__o21a_1 _07523_ (.A1(net811),
    .A2(_02537_),
    .B1(net793),
    .X(_02540_));
 sky130_fd_sc_hd__mux4_1 _07524_ (.A0(\reg_module.gprf[638] ),
    .A1(\reg_module.gprf[606] ),
    .A2(\reg_module.gprf[574] ),
    .A3(\reg_module.gprf[542] ),
    .S0(net931),
    .S1(net895),
    .X(_02541_));
 sky130_fd_sc_hd__mux4_1 _07525_ (.A0(\reg_module.gprf[766] ),
    .A1(\reg_module.gprf[734] ),
    .A2(\reg_module.gprf[702] ),
    .A3(\reg_module.gprf[670] ),
    .S0(net926),
    .S1(net890),
    .X(_02542_));
 sky130_fd_sc_hd__mux2_1 _07526_ (.A0(_02541_),
    .A1(_02542_),
    .S(net810),
    .X(_02543_));
 sky130_fd_sc_hd__a221o_1 _07527_ (.A1(_02539_),
    .A2(_02540_),
    .B1(_02543_),
    .B2(net856),
    .C1(net942),
    .X(_02544_));
 sky130_fd_sc_hd__mux4_1 _07528_ (.A0(\reg_module.gprf[382] ),
    .A1(\reg_module.gprf[350] ),
    .A2(\reg_module.gprf[318] ),
    .A3(\reg_module.gprf[286] ),
    .S0(net931),
    .S1(net895),
    .X(_02545_));
 sky130_fd_sc_hd__mux4_1 _07529_ (.A0(\reg_module.gprf[510] ),
    .A1(\reg_module.gprf[478] ),
    .A2(\reg_module.gprf[446] ),
    .A3(\reg_module.gprf[414] ),
    .S0(net931),
    .S1(net895),
    .X(_02546_));
 sky130_fd_sc_hd__mux2_1 _07530_ (.A0(_02545_),
    .A1(_02546_),
    .S(net810),
    .X(_02547_));
 sky130_fd_sc_hd__mux4_1 _07531_ (.A0(\reg_module.gprf[126] ),
    .A1(\reg_module.gprf[94] ),
    .A2(\reg_module.gprf[62] ),
    .A3(\reg_module.gprf[30] ),
    .S0(net931),
    .S1(net895),
    .X(_02548_));
 sky130_fd_sc_hd__mux4_1 _07532_ (.A0(\reg_module.gprf[254] ),
    .A1(\reg_module.gprf[222] ),
    .A2(\reg_module.gprf[190] ),
    .A3(\reg_module.gprf[158] ),
    .S0(net926),
    .S1(net890),
    .X(_02549_));
 sky130_fd_sc_hd__or2_1 _07533_ (.A(net864),
    .B(_02549_),
    .X(_02550_));
 sky130_fd_sc_hd__o211a_1 _07534_ (.A1(net810),
    .A2(_02548_),
    .B1(_02550_),
    .C1(net855),
    .X(_02551_));
 sky130_fd_sc_hd__a21o_1 _07535_ (.A1(net794),
    .A2(_02547_),
    .B1(net786),
    .X(_02552_));
 sky130_fd_sc_hd__o211a_1 _07536_ (.A1(_02551_),
    .A2(_02552_),
    .B1(net586),
    .C1(_02544_),
    .X(_02553_));
 sky130_fd_sc_hd__a21o_1 _07537_ (.A1(\rWrDataWB[30] ),
    .A2(net578),
    .B1(net612),
    .X(_02554_));
 sky130_fd_sc_hd__o22a_1 _07538_ (.A1(\rWrData[30] ),
    .A2(net606),
    .B1(_02553_),
    .B2(_02554_),
    .X(net126));
 sky130_fd_sc_hd__mux4_1 _07539_ (.A0(\reg_module.gprf[895] ),
    .A1(\reg_module.gprf[863] ),
    .A2(\reg_module.gprf[831] ),
    .A3(\reg_module.gprf[799] ),
    .S0(net933),
    .S1(net897),
    .X(_02555_));
 sky130_fd_sc_hd__mux4_1 _07540_ (.A0(\reg_module.gprf[1023] ),
    .A1(\reg_module.gprf[991] ),
    .A2(\reg_module.gprf[959] ),
    .A3(\reg_module.gprf[927] ),
    .S0(net934),
    .S1(net897),
    .X(_02556_));
 sky130_fd_sc_hd__or2_1 _07541_ (.A(net864),
    .B(_02556_),
    .X(_02557_));
 sky130_fd_sc_hd__o21a_1 _07542_ (.A1(net809),
    .A2(_02555_),
    .B1(net793),
    .X(_02558_));
 sky130_fd_sc_hd__mux4_1 _07543_ (.A0(\reg_module.gprf[639] ),
    .A1(\reg_module.gprf[607] ),
    .A2(\reg_module.gprf[575] ),
    .A3(\reg_module.gprf[543] ),
    .S0(net933),
    .S1(net897),
    .X(_02559_));
 sky130_fd_sc_hd__mux4_1 _07544_ (.A0(\reg_module.gprf[767] ),
    .A1(\reg_module.gprf[735] ),
    .A2(\reg_module.gprf[703] ),
    .A3(\reg_module.gprf[671] ),
    .S0(net931),
    .S1(net896),
    .X(_02560_));
 sky130_fd_sc_hd__mux2_1 _07545_ (.A0(_02559_),
    .A1(_02560_),
    .S(net810),
    .X(_02561_));
 sky130_fd_sc_hd__a221o_1 _07546_ (.A1(_02557_),
    .A2(_02558_),
    .B1(_02561_),
    .B2(net855),
    .C1(net942),
    .X(_02562_));
 sky130_fd_sc_hd__mux4_1 _07547_ (.A0(\reg_module.gprf[383] ),
    .A1(\reg_module.gprf[351] ),
    .A2(\reg_module.gprf[319] ),
    .A3(\reg_module.gprf[287] ),
    .S0(net933),
    .S1(net897),
    .X(_02563_));
 sky130_fd_sc_hd__mux4_1 _07548_ (.A0(\reg_module.gprf[511] ),
    .A1(\reg_module.gprf[479] ),
    .A2(\reg_module.gprf[447] ),
    .A3(\reg_module.gprf[415] ),
    .S0(net933),
    .S1(net897),
    .X(_02564_));
 sky130_fd_sc_hd__mux2_1 _07549_ (.A0(_02563_),
    .A1(_02564_),
    .S(net809),
    .X(_02565_));
 sky130_fd_sc_hd__mux4_1 _07550_ (.A0(\reg_module.gprf[127] ),
    .A1(\reg_module.gprf[95] ),
    .A2(\reg_module.gprf[63] ),
    .A3(\reg_module.gprf[31] ),
    .S0(net933),
    .S1(net897),
    .X(_02566_));
 sky130_fd_sc_hd__or2_1 _07551_ (.A(net810),
    .B(_02566_),
    .X(_02567_));
 sky130_fd_sc_hd__mux4_1 _07552_ (.A0(\reg_module.gprf[255] ),
    .A1(\reg_module.gprf[223] ),
    .A2(\reg_module.gprf[191] ),
    .A3(\reg_module.gprf[159] ),
    .S0(net933),
    .S1(net897),
    .X(_02568_));
 sky130_fd_sc_hd__o211a_1 _07553_ (.A1(net864),
    .A2(_02568_),
    .B1(_02567_),
    .C1(net855),
    .X(_02569_));
 sky130_fd_sc_hd__a21o_1 _07554_ (.A1(net793),
    .A2(_02565_),
    .B1(net786),
    .X(_02570_));
 sky130_fd_sc_hd__o211a_1 _07555_ (.A1(_02569_),
    .A2(_02570_),
    .B1(net586),
    .C1(_02562_),
    .X(_02571_));
 sky130_fd_sc_hd__a21o_1 _07556_ (.A1(\rWrDataWB[31] ),
    .A2(net580),
    .B1(net615),
    .X(_02572_));
 sky130_fd_sc_hd__o22a_1 _07557_ (.A1(\rWrData[31] ),
    .A2(net608),
    .B1(_02571_),
    .B2(_02572_),
    .X(net127));
 sky130_fd_sc_hd__nor2_1 _07558_ (.A(\alu.op_consShf ),
    .B(\dec.op_intRegImm ),
    .Y(_02573_));
 sky130_fd_sc_hd__or2_1 _07559_ (.A(\alu.op_consShf ),
    .B(\dec.op_intRegImm ),
    .X(_02574_));
 sky130_fd_sc_hd__nor3_1 _07560_ (.A(net948),
    .B(\alu.r_type ),
    .C(net764),
    .Y(_02575_));
 sky130_fd_sc_hd__or3_1 _07561_ (.A(net948),
    .B(\alu.r_type ),
    .C(net765),
    .X(_02576_));
 sky130_fd_sc_hd__nor2_2 _07562_ (.A(\alu.b_type ),
    .B(\alu.r_type ),
    .Y(_02577_));
 sky130_fd_sc_hd__or2_2 _07563_ (.A(\alu.b_type ),
    .B(\alu.r_type ),
    .X(_02578_));
 sky130_fd_sc_hd__nor2_4 _07564_ (.A(net764),
    .B(net759),
    .Y(_02579_));
 sky130_fd_sc_hd__nand2_1 _07565_ (.A(net767),
    .B(net763),
    .Y(_02580_));
 sky130_fd_sc_hd__and3_2 _07566_ (.A(net948),
    .B(net770),
    .C(net760),
    .X(_02581_));
 sky130_fd_sc_hd__nand2_2 _07567_ (.A(net949),
    .B(_02579_),
    .Y(_02582_));
 sky130_fd_sc_hd__nand2_1 _07568_ (.A(net159),
    .B(net733),
    .Y(_02583_));
 sky130_fd_sc_hd__nor2_1 _07569_ (.A(_01215_),
    .B(net980),
    .Y(_02584_));
 sky130_fd_sc_hd__a21oi_2 _07570_ (.A1(net26),
    .A2(net980),
    .B1(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__a21o_1 _07571_ (.A1(net26),
    .A2(net980),
    .B1(_02584_),
    .X(_02586_));
 sky130_fd_sc_hd__mux2_1 _07572_ (.A0(_01969_),
    .A1(net574),
    .S(net594),
    .X(_02587_));
 sky130_fd_sc_hd__a211o_1 _07573_ (.A1(net620),
    .A2(_02587_),
    .B1(_02579_),
    .C1(_01953_),
    .X(_02588_));
 sky130_fd_sc_hd__and2_1 _07574_ (.A(_02583_),
    .B(_02588_),
    .X(_02589_));
 sky130_fd_sc_hd__a21o_1 _07575_ (.A1(net944),
    .A2(net764),
    .B1(net759),
    .X(_02590_));
 sky130_fd_sc_hd__a31o_1 _07576_ (.A1(net949),
    .A2(net842),
    .A3(net769),
    .B1(net726),
    .X(_02591_));
 sky130_fd_sc_hd__a21o_1 _07577_ (.A1(net580),
    .A2(_02586_),
    .B1(net614),
    .X(_02592_));
 sky130_fd_sc_hd__o22a_1 _07578_ (.A1(\rWrData[31] ),
    .A2(net608),
    .B1(_02571_),
    .B2(_02592_),
    .X(_02593_));
 sky130_fd_sc_hd__o21a_1 _07579_ (.A1(net762),
    .A2(_02593_),
    .B1(_02591_),
    .X(_02594_));
 sky130_fd_sc_hd__o21ai_1 _07580_ (.A1(net762),
    .A2(_02593_),
    .B1(_02591_),
    .Y(_02595_));
 sky130_fd_sc_hd__nand2_1 _07581_ (.A(net199),
    .B(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__nor2_1 _07582_ (.A(net199),
    .B(_02595_),
    .Y(_02597_));
 sky130_fd_sc_hd__and3_2 _07583_ (.A(_02583_),
    .B(_02588_),
    .C(_02594_),
    .X(_02598_));
 sky130_fd_sc_hd__nand2_1 _07584_ (.A(net199),
    .B(_02594_),
    .Y(_02599_));
 sky130_fd_sc_hd__a21oi_2 _07585_ (.A1(_02583_),
    .A2(_02588_),
    .B1(_02594_),
    .Y(_02600_));
 sky130_fd_sc_hd__nor2_2 _07586_ (.A(_02598_),
    .B(_02600_),
    .Y(_02601_));
 sky130_fd_sc_hd__inv_2 _07587_ (.A(_02601_),
    .Y(_02602_));
 sky130_fd_sc_hd__and2b_1 _07588_ (.A_N(net971),
    .B(\rWrDataWB[6] ),
    .X(_02603_));
 sky130_fd_sc_hd__a21oi_1 _07589_ (.A1(net971),
    .A2(net30),
    .B1(_02603_),
    .Y(_02604_));
 sky130_fd_sc_hd__a21o_1 _07590_ (.A1(net971),
    .A2(net30),
    .B1(_02603_),
    .X(_02605_));
 sky130_fd_sc_hd__nand2_1 _07591_ (.A(net587),
    .B(_02605_),
    .Y(_02606_));
 sky130_fd_sc_hd__o211a_1 _07592_ (.A1(net587),
    .A2(_01412_),
    .B1(_02606_),
    .C1(net616),
    .X(_02607_));
 sky130_fd_sc_hd__o21ai_1 _07593_ (.A1(\rWrData[6] ),
    .A2(net616),
    .B1(net734),
    .Y(_02608_));
 sky130_fd_sc_hd__o2bb2a_4 _07594_ (.A1_N(net163),
    .A2_N(net728),
    .B1(_02607_),
    .B2(_02608_),
    .X(_02609_));
 sky130_fd_sc_hd__inv_2 _07595_ (.A(_02609_),
    .Y(_02610_));
 sky130_fd_sc_hd__a21o_1 _07596_ (.A1(net575),
    .A2(_02605_),
    .B1(net609),
    .X(_02611_));
 sky130_fd_sc_hd__o22a_1 _07597_ (.A1(\rWrData[6] ),
    .A2(net601),
    .B1(_02117_),
    .B2(_02611_),
    .X(_02612_));
 sky130_fd_sc_hd__a21o_1 _07598_ (.A1(\brancher.imm12_i_s[6] ),
    .A2(net764),
    .B1(net759),
    .X(_02613_));
 sky130_fd_sc_hd__o21a_2 _07599_ (.A1(net761),
    .A2(_02612_),
    .B1(_02613_),
    .X(_02614_));
 sky130_fd_sc_hd__and2_1 _07600_ (.A(_02610_),
    .B(_02614_),
    .X(_02615_));
 sky130_fd_sc_hd__inv_2 _07601_ (.A(_02615_),
    .Y(_02616_));
 sky130_fd_sc_hd__or2_1 _07602_ (.A(_02610_),
    .B(_02614_),
    .X(_02617_));
 sky130_fd_sc_hd__nor2_1 _07603_ (.A(_02609_),
    .B(_02614_),
    .Y(_02618_));
 sky130_fd_sc_hd__or2_1 _07604_ (.A(_02609_),
    .B(_02614_),
    .X(_02619_));
 sky130_fd_sc_hd__xnor2_1 _07605_ (.A(_02609_),
    .B(_02614_),
    .Y(_02620_));
 sky130_fd_sc_hd__nand2_1 _07606_ (.A(_02616_),
    .B(_02617_),
    .Y(_02621_));
 sky130_fd_sc_hd__and2b_1 _07607_ (.A_N(net973),
    .B(\rWrDataWB[7] ),
    .X(_02622_));
 sky130_fd_sc_hd__a21oi_1 _07608_ (.A1(net973),
    .A2(net31),
    .B1(_02622_),
    .Y(_02623_));
 sky130_fd_sc_hd__a21o_1 _07609_ (.A1(net973),
    .A2(net31),
    .B1(_02622_),
    .X(_02624_));
 sky130_fd_sc_hd__a211o_1 _07610_ (.A1(net587),
    .A2(_02624_),
    .B1(_01438_),
    .C1(net622),
    .X(_02625_));
 sky130_fd_sc_hd__o21a_1 _07611_ (.A1(\rWrData[7] ),
    .A2(net616),
    .B1(net734),
    .X(_02626_));
 sky130_fd_sc_hd__a22oi_4 _07612_ (.A1(net164),
    .A2(net728),
    .B1(_02625_),
    .B2(_02626_),
    .Y(_02627_));
 sky130_fd_sc_hd__inv_2 _07613_ (.A(_02627_),
    .Y(_02628_));
 sky130_fd_sc_hd__a21o_1 _07614_ (.A1(net575),
    .A2(_02624_),
    .B1(net609),
    .X(_02629_));
 sky130_fd_sc_hd__o22a_1 _07615_ (.A1(\rWrData[7] ),
    .A2(net601),
    .B1(_02135_),
    .B2(_02629_),
    .X(_02630_));
 sky130_fd_sc_hd__a21o_1 _07616_ (.A1(\brancher.imm12_i_s[7] ),
    .A2(net764),
    .B1(net759),
    .X(_02631_));
 sky130_fd_sc_hd__o21a_2 _07617_ (.A1(net761),
    .A2(_02630_),
    .B1(_02631_),
    .X(_02632_));
 sky130_fd_sc_hd__and2_1 _07618_ (.A(_02628_),
    .B(_02632_),
    .X(_02633_));
 sky130_fd_sc_hd__inv_2 _07619_ (.A(_02633_),
    .Y(_02634_));
 sky130_fd_sc_hd__or2_1 _07620_ (.A(_02628_),
    .B(_02632_),
    .X(_02635_));
 sky130_fd_sc_hd__nand2_1 _07621_ (.A(_02627_),
    .B(_02632_),
    .Y(_02636_));
 sky130_fd_sc_hd__nor2_1 _07622_ (.A(_02627_),
    .B(_02632_),
    .Y(_02637_));
 sky130_fd_sc_hd__xnor2_2 _07623_ (.A(_02627_),
    .B(_02632_),
    .Y(_02638_));
 sky130_fd_sc_hd__or2_1 _07624_ (.A(_02620_),
    .B(_02638_),
    .X(_02639_));
 sky130_fd_sc_hd__nand2b_1 _07625_ (.A_N(net28),
    .B(net974),
    .Y(_02640_));
 sky130_fd_sc_hd__o21a_1 _07626_ (.A1(net974),
    .A2(\rWrDataWB[4] ),
    .B1(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__o21ai_2 _07627_ (.A1(net974),
    .A2(\rWrDataWB[4] ),
    .B1(_02640_),
    .Y(_02642_));
 sky130_fd_sc_hd__nor2_1 _07628_ (.A(net584),
    .B(net723),
    .Y(_02643_));
 sky130_fd_sc_hd__o21ai_2 _07629_ (.A1(_02081_),
    .A2(_02643_),
    .B1(net603),
    .Y(_02644_));
 sky130_fd_sc_hd__a21oi_2 _07630_ (.A1(\brancher.imm12_i_s[4] ),
    .A2(net765),
    .B1(net758),
    .Y(_02645_));
 sky130_fd_sc_hd__a31oi_4 _07631_ (.A1(_02064_),
    .A2(net758),
    .A3(_02644_),
    .B1(_02645_),
    .Y(_02646_));
 sky130_fd_sc_hd__a31o_1 _07632_ (.A1(_02064_),
    .A2(net758),
    .A3(_02644_),
    .B1(_02645_),
    .X(_02647_));
 sky130_fd_sc_hd__a211o_1 _07633_ (.A1(net589),
    .A2(_02641_),
    .B1(_01368_),
    .C1(net624),
    .X(_02648_));
 sky130_fd_sc_hd__o21a_1 _07634_ (.A1(\rWrData[4] ),
    .A2(net617),
    .B1(net736),
    .X(_02649_));
 sky130_fd_sc_hd__a22oi_4 _07635_ (.A1(net161),
    .A2(net730),
    .B1(_02648_),
    .B2(_02649_),
    .Y(_02650_));
 sky130_fd_sc_hd__or2_1 _07636_ (.A(net194),
    .B(_02650_),
    .X(_02651_));
 sky130_fd_sc_hd__xnor2_4 _07637_ (.A(net194),
    .B(_02650_),
    .Y(_02652_));
 sky130_fd_sc_hd__and2b_1 _07638_ (.A_N(net973),
    .B(\rWrDataWB[5] ),
    .X(_02653_));
 sky130_fd_sc_hd__a21oi_1 _07639_ (.A1(net973),
    .A2(net29),
    .B1(_02653_),
    .Y(_02654_));
 sky130_fd_sc_hd__a21o_1 _07640_ (.A1(net973),
    .A2(net29),
    .B1(_02653_),
    .X(_02655_));
 sky130_fd_sc_hd__nor2_1 _07641_ (.A(net595),
    .B(_02654_),
    .Y(_02656_));
 sky130_fd_sc_hd__a211o_1 _07642_ (.A1(net595),
    .A2(_01389_),
    .B1(_02656_),
    .C1(net622),
    .X(_02657_));
 sky130_fd_sc_hd__o21a_1 _07643_ (.A1(\rWrData[5] ),
    .A2(net617),
    .B1(net734),
    .X(_02658_));
 sky130_fd_sc_hd__a22oi_4 _07644_ (.A1(net162),
    .A2(net728),
    .B1(_02657_),
    .B2(_02658_),
    .Y(_02659_));
 sky130_fd_sc_hd__a21o_1 _07645_ (.A1(net577),
    .A2(_02655_),
    .B1(net610),
    .X(_02660_));
 sky130_fd_sc_hd__o22a_1 _07646_ (.A1(\rWrData[5] ),
    .A2(net602),
    .B1(_02099_),
    .B2(_02660_),
    .X(_02661_));
 sky130_fd_sc_hd__a21o_1 _07647_ (.A1(\brancher.imm12_i_s[5] ),
    .A2(net764),
    .B1(net759),
    .X(_02662_));
 sky130_fd_sc_hd__o21a_2 _07648_ (.A1(net761),
    .A2(_02661_),
    .B1(_02662_),
    .X(_02663_));
 sky130_fd_sc_hd__or2_1 _07649_ (.A(_02659_),
    .B(_02663_),
    .X(_02664_));
 sky130_fd_sc_hd__and2_1 _07650_ (.A(_02659_),
    .B(_02663_),
    .X(_02665_));
 sky130_fd_sc_hd__and2b_1 _07651_ (.A_N(_02659_),
    .B(_02663_),
    .X(_02666_));
 sky130_fd_sc_hd__nand2b_1 _07652_ (.A_N(_02659_),
    .B(_02663_),
    .Y(_02667_));
 sky130_fd_sc_hd__nand2b_1 _07653_ (.A_N(_02663_),
    .B(_02659_),
    .Y(_02668_));
 sky130_fd_sc_hd__and2_2 _07654_ (.A(_02667_),
    .B(_02668_),
    .X(_02669_));
 sky130_fd_sc_hd__or3_1 _07655_ (.A(_02639_),
    .B(_02652_),
    .C(_02669_),
    .X(_02670_));
 sky130_fd_sc_hd__nand2b_1 _07656_ (.A_N(net13),
    .B(net974),
    .Y(_02671_));
 sky130_fd_sc_hd__o21a_1 _07657_ (.A1(net974),
    .A2(\rWrDataWB[1] ),
    .B1(_02671_),
    .X(_02672_));
 sky130_fd_sc_hd__o21ai_2 _07658_ (.A1(net974),
    .A2(\rWrDataWB[1] ),
    .B1(_02671_),
    .Y(_02673_));
 sky130_fd_sc_hd__nand2_1 _07659_ (.A(net589),
    .B(_02672_),
    .Y(_02674_));
 sky130_fd_sc_hd__a21oi_1 _07660_ (.A1(_01303_),
    .A2(_02674_),
    .B1(net624),
    .Y(_02675_));
 sky130_fd_sc_hd__o21ai_2 _07661_ (.A1(_01287_),
    .A2(_02675_),
    .B1(net736),
    .Y(_02676_));
 sky130_fd_sc_hd__nand2_1 _07662_ (.A(net146),
    .B(net730),
    .Y(_02677_));
 sky130_fd_sc_hd__and2_1 _07663_ (.A(_02676_),
    .B(_02677_),
    .X(_02678_));
 sky130_fd_sc_hd__nor2_1 _07664_ (.A(net584),
    .B(net721),
    .Y(_02679_));
 sky130_fd_sc_hd__o21a_1 _07665_ (.A1(_02024_),
    .A2(_02679_),
    .B1(net603),
    .X(_02680_));
 sky130_fd_sc_hd__or2_1 _07666_ (.A(\brancher.imm12_i_s[1] ),
    .B(net758),
    .X(_02681_));
 sky130_fd_sc_hd__o311a_2 _07667_ (.A1(_02007_),
    .A2(net760),
    .A3(_02680_),
    .B1(_02681_),
    .C1(net736),
    .X(_02682_));
 sky130_fd_sc_hd__o311ai_2 _07668_ (.A1(_02007_),
    .A2(net760),
    .A3(_02680_),
    .B1(_02681_),
    .C1(net736),
    .Y(_02683_));
 sky130_fd_sc_hd__and2b_1 _07669_ (.A_N(net973),
    .B(\rWrDataWB[0] ),
    .X(_02684_));
 sky130_fd_sc_hd__a21oi_4 _07670_ (.A1(net973),
    .A2(net2),
    .B1(_02684_),
    .Y(_02685_));
 sky130_fd_sc_hd__a21o_2 _07671_ (.A1(net973),
    .A2(net2),
    .B1(_02684_),
    .X(_02686_));
 sky130_fd_sc_hd__nand2_1 _07672_ (.A(net577),
    .B(_02685_),
    .Y(_02687_));
 sky130_fd_sc_hd__a21oi_2 _07673_ (.A1(_02005_),
    .A2(_02687_),
    .B1(net610),
    .Y(_02688_));
 sky130_fd_sc_hd__o21a_1 _07674_ (.A1(_01973_),
    .A2(_02688_),
    .B1(net758),
    .X(_02689_));
 sky130_fd_sc_hd__o21ai_1 _07675_ (.A1(_01973_),
    .A2(_02688_),
    .B1(net758),
    .Y(_02690_));
 sky130_fd_sc_hd__a21oi_1 _07676_ (.A1(\brancher.imm12_i_s[0] ),
    .A2(net765),
    .B1(net758),
    .Y(_02691_));
 sky130_fd_sc_hd__a21o_1 _07677_ (.A1(\brancher.imm12_i_s[0] ),
    .A2(net765),
    .B1(net758),
    .X(_02692_));
 sky130_fd_sc_hd__nor2_2 _07678_ (.A(net233),
    .B(net718),
    .Y(_02693_));
 sky130_fd_sc_hd__nand2_1 _07679_ (.A(net230),
    .B(net715),
    .Y(_02694_));
 sky130_fd_sc_hd__nor2_1 _07680_ (.A(net595),
    .B(_02686_),
    .Y(_02695_));
 sky130_fd_sc_hd__o21ai_2 _07681_ (.A1(_01280_),
    .A2(_02695_),
    .B1(net617),
    .Y(_02696_));
 sky130_fd_sc_hd__a32oi_4 _07682_ (.A1(_01252_),
    .A2(net739),
    .A3(_02696_),
    .B1(net730),
    .B2(net135),
    .Y(_02697_));
 sky130_fd_sc_hd__a21oi_1 _07683_ (.A1(net229),
    .A2(net714),
    .B1(_02697_),
    .Y(_02698_));
 sky130_fd_sc_hd__o21ba_1 _07684_ (.A1(net236),
    .A2(_02698_),
    .B1_N(_02678_),
    .X(_02699_));
 sky130_fd_sc_hd__and2_2 _07685_ (.A(net236),
    .B(_02698_),
    .X(_02700_));
 sky130_fd_sc_hd__nand2b_1 _07686_ (.A_N(net24),
    .B(net975),
    .Y(_02701_));
 sky130_fd_sc_hd__o21a_2 _07687_ (.A1(net975),
    .A2(\rWrDataWB[2] ),
    .B1(_02701_),
    .X(_02702_));
 sky130_fd_sc_hd__o21ai_2 _07688_ (.A1(net975),
    .A2(\rWrDataWB[2] ),
    .B1(_02701_),
    .Y(_02703_));
 sky130_fd_sc_hd__nand2_1 _07689_ (.A(net582),
    .B(_02702_),
    .Y(_02704_));
 sky130_fd_sc_hd__a21o_1 _07690_ (.A1(_02043_),
    .A2(_02704_),
    .B1(net610),
    .X(_02705_));
 sky130_fd_sc_hd__a21oi_2 _07691_ (.A1(\brancher.imm12_i_s[2] ),
    .A2(net765),
    .B1(net758),
    .Y(_02706_));
 sky130_fd_sc_hd__a31oi_4 _07692_ (.A1(_02026_),
    .A2(_02578_),
    .A3(_02705_),
    .B1(_02706_),
    .Y(_02707_));
 sky130_fd_sc_hd__a31o_2 _07693_ (.A1(_02026_),
    .A2(_02578_),
    .A3(_02705_),
    .B1(_02706_),
    .X(_02708_));
 sky130_fd_sc_hd__nor2_1 _07694_ (.A(net597),
    .B(_02703_),
    .Y(_02709_));
 sky130_fd_sc_hd__a211o_1 _07695_ (.A1(net597),
    .A2(_01326_),
    .B1(_02709_),
    .C1(net623),
    .X(_02710_));
 sky130_fd_sc_hd__a32oi_4 _07696_ (.A1(_01310_),
    .A2(net736),
    .A3(_02710_),
    .B1(net730),
    .B2(net157),
    .Y(_02711_));
 sky130_fd_sc_hd__nand2_1 _07697_ (.A(net226),
    .B(_02711_),
    .Y(_02712_));
 sky130_fd_sc_hd__or2_2 _07698_ (.A(net226),
    .B(_02711_),
    .X(_02713_));
 sky130_fd_sc_hd__nand2_2 _07699_ (.A(_02712_),
    .B(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__nand2b_1 _07700_ (.A_N(net27),
    .B(net971),
    .Y(_02715_));
 sky130_fd_sc_hd__o21a_1 _07701_ (.A1(net971),
    .A2(\rWrDataWB[3] ),
    .B1(_02715_),
    .X(_02716_));
 sky130_fd_sc_hd__o21ai_4 _07702_ (.A1(net972),
    .A2(\rWrDataWB[3] ),
    .B1(_02715_),
    .Y(_02717_));
 sky130_fd_sc_hd__nor2_1 _07703_ (.A(net584),
    .B(_02717_),
    .Y(_02718_));
 sky130_fd_sc_hd__o21ai_1 _07704_ (.A1(_02062_),
    .A2(_02718_),
    .B1(net602),
    .Y(_02719_));
 sky130_fd_sc_hd__a21oi_1 _07705_ (.A1(\rWrData[3] ),
    .A2(net610),
    .B1(net760),
    .Y(_02720_));
 sky130_fd_sc_hd__a21oi_1 _07706_ (.A1(\brancher.imm12_i_s[3] ),
    .A2(net764),
    .B1(net758),
    .Y(_02721_));
 sky130_fd_sc_hd__a21oi_1 _07707_ (.A1(_02719_),
    .A2(_02720_),
    .B1(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__a21o_1 _07708_ (.A1(_02719_),
    .A2(_02720_),
    .B1(_02721_),
    .X(_02723_));
 sky130_fd_sc_hd__nor2_1 _07709_ (.A(net597),
    .B(_02717_),
    .Y(_02724_));
 sky130_fd_sc_hd__a211o_1 _07710_ (.A1(net597),
    .A2(_01346_),
    .B1(_02724_),
    .C1(net624),
    .X(_02725_));
 sky130_fd_sc_hd__o21a_1 _07711_ (.A1(\rWrData[3] ),
    .A2(net617),
    .B1(net736),
    .X(_02726_));
 sky130_fd_sc_hd__a22oi_4 _07712_ (.A1(net160),
    .A2(net730),
    .B1(_02725_),
    .B2(_02726_),
    .Y(_02727_));
 sky130_fd_sc_hd__nand2_1 _07713_ (.A(net207),
    .B(_02727_),
    .Y(_02728_));
 sky130_fd_sc_hd__nor2_1 _07714_ (.A(net207),
    .B(_02727_),
    .Y(_02729_));
 sky130_fd_sc_hd__or2_1 _07715_ (.A(net210),
    .B(_02727_),
    .X(_02730_));
 sky130_fd_sc_hd__and2_1 _07716_ (.A(net210),
    .B(_02727_),
    .X(_02731_));
 sky130_fd_sc_hd__nand2_1 _07717_ (.A(net210),
    .B(_02727_),
    .Y(_02732_));
 sky130_fd_sc_hd__nand2_1 _07718_ (.A(_02730_),
    .B(_02732_),
    .Y(_02733_));
 sky130_fd_sc_hd__or4_1 _07719_ (.A(_02699_),
    .B(_02700_),
    .C(_02714_),
    .D(_02733_),
    .X(_02734_));
 sky130_fd_sc_hd__nand2b_1 _07720_ (.A_N(_02712_),
    .B(_02730_),
    .Y(_02735_));
 sky130_fd_sc_hd__a31o_1 _07721_ (.A1(_02732_),
    .A2(_02734_),
    .A3(_02735_),
    .B1(_02670_),
    .X(_02736_));
 sky130_fd_sc_hd__a21o_1 _07722_ (.A1(net194),
    .A2(_02650_),
    .B1(_02665_),
    .X(_02737_));
 sky130_fd_sc_hd__nand2_1 _07723_ (.A(_02664_),
    .B(_02737_),
    .Y(_02738_));
 sky130_fd_sc_hd__a21boi_1 _07724_ (.A1(_02609_),
    .A2(_02614_),
    .B1_N(_02636_),
    .Y(_02739_));
 sky130_fd_sc_hd__o22a_1 _07725_ (.A1(_02639_),
    .A2(_02738_),
    .B1(_02739_),
    .B2(_02637_),
    .X(_02740_));
 sky130_fd_sc_hd__and2b_1 _07726_ (.A_N(net981),
    .B(\rWrDataWB[30] ),
    .X(_02741_));
 sky130_fd_sc_hd__a21oi_1 _07727_ (.A1(net981),
    .A2(net25),
    .B1(_02741_),
    .Y(_02742_));
 sky130_fd_sc_hd__a21o_1 _07728_ (.A1(net981),
    .A2(net25),
    .B1(_02741_),
    .X(_02743_));
 sky130_fd_sc_hd__a211o_1 _07729_ (.A1(net590),
    .A2(_02743_),
    .B1(_01948_),
    .C1(net625),
    .X(_02744_));
 sky130_fd_sc_hd__o21a_1 _07730_ (.A1(\rWrData[30] ),
    .A2(net620),
    .B1(net739),
    .X(_02745_));
 sky130_fd_sc_hd__a22oi_4 _07731_ (.A1(net158),
    .A2(net733),
    .B1(_02744_),
    .B2(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__a31o_1 _07732_ (.A1(net950),
    .A2(\brancher.imm13_b[10] ),
    .A3(net768),
    .B1(net726),
    .X(_02747_));
 sky130_fd_sc_hd__a21o_1 _07733_ (.A1(net580),
    .A2(_02743_),
    .B1(net614),
    .X(_02748_));
 sky130_fd_sc_hd__o22a_1 _07734_ (.A1(\rWrData[30] ),
    .A2(net607),
    .B1(_02553_),
    .B2(_02748_),
    .X(_02749_));
 sky130_fd_sc_hd__o21a_1 _07735_ (.A1(net762),
    .A2(_02749_),
    .B1(_02747_),
    .X(_02750_));
 sky130_fd_sc_hd__nor2_1 _07736_ (.A(_02746_),
    .B(_02750_),
    .Y(_02751_));
 sky130_fd_sc_hd__xnor2_2 _07737_ (.A(_02746_),
    .B(_02750_),
    .Y(_02752_));
 sky130_fd_sc_hd__nor3_1 _07738_ (.A(_02598_),
    .B(_02600_),
    .C(_02752_),
    .Y(_02753_));
 sky130_fd_sc_hd__or2_1 _07739_ (.A(_02602_),
    .B(_02752_),
    .X(_02754_));
 sky130_fd_sc_hd__and2b_1 _07740_ (.A_N(net978),
    .B(\rWrDataWB[28] ),
    .X(_02755_));
 sky130_fd_sc_hd__a21oi_1 _07741_ (.A1(net977),
    .A2(net22),
    .B1(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__a21o_2 _07742_ (.A1(net977),
    .A2(net22),
    .B1(_02755_),
    .X(_02757_));
 sky130_fd_sc_hd__a21oi_1 _07743_ (.A1(net591),
    .A2(_02757_),
    .B1(net625),
    .Y(_02758_));
 sky130_fd_sc_hd__o21ai_2 _07744_ (.A1(net591),
    .A2(_01906_),
    .B1(_02758_),
    .Y(_02759_));
 sky130_fd_sc_hd__a32oi_4 _07745_ (.A1(_01890_),
    .A2(net738),
    .A3(_02759_),
    .B1(net732),
    .B2(net155),
    .Y(_02760_));
 sky130_fd_sc_hd__a32o_2 _07746_ (.A1(_01890_),
    .A2(net738),
    .A3(_02759_),
    .B1(net732),
    .B2(net155),
    .X(_02761_));
 sky130_fd_sc_hd__a31o_1 _07747_ (.A1(net949),
    .A2(\brancher.imm13_b[8] ),
    .A3(net769),
    .B1(net726),
    .X(_02762_));
 sky130_fd_sc_hd__a21o_1 _07748_ (.A1(net578),
    .A2(_02757_),
    .B1(net612),
    .X(_02763_));
 sky130_fd_sc_hd__a31o_1 _07749_ (.A1(net586),
    .A2(_02508_),
    .A3(_02516_),
    .B1(_02763_),
    .X(_02764_));
 sky130_fd_sc_hd__a21o_1 _07750_ (.A1(_02500_),
    .A2(_02764_),
    .B1(net763),
    .X(_02765_));
 sky130_fd_sc_hd__and3_1 _07751_ (.A(_02760_),
    .B(_02762_),
    .C(_02765_),
    .X(_02766_));
 sky130_fd_sc_hd__a21o_1 _07752_ (.A1(_02762_),
    .A2(_02765_),
    .B1(_02760_),
    .X(_02767_));
 sky130_fd_sc_hd__nand2b_2 _07753_ (.A_N(_02766_),
    .B(_02767_),
    .Y(_02768_));
 sky130_fd_sc_hd__and2b_1 _07754_ (.A_N(net977),
    .B(\rWrDataWB[29] ),
    .X(_02769_));
 sky130_fd_sc_hd__a21oi_1 _07755_ (.A1(net978),
    .A2(net23),
    .B1(_02769_),
    .Y(_02770_));
 sky130_fd_sc_hd__a21o_1 _07756_ (.A1(net978),
    .A2(net23),
    .B1(_02769_),
    .X(_02771_));
 sky130_fd_sc_hd__o211a_1 _07757_ (.A1(net598),
    .A2(_02770_),
    .B1(_01929_),
    .C1(net619),
    .X(_02772_));
 sky130_fd_sc_hd__o32a_2 _07758_ (.A1(_01912_),
    .A2(_02579_),
    .A3(_02772_),
    .B1(_02582_),
    .B2(_01203_),
    .X(_02773_));
 sky130_fd_sc_hd__a31o_1 _07759_ (.A1(net949),
    .A2(\brancher.imm13_b[9] ),
    .A3(net767),
    .B1(_02590_),
    .X(_02774_));
 sky130_fd_sc_hd__a21o_1 _07760_ (.A1(net578),
    .A2(_02771_),
    .B1(net612),
    .X(_02775_));
 sky130_fd_sc_hd__o22a_1 _07761_ (.A1(\rWrData[29] ),
    .A2(net606),
    .B1(_02535_),
    .B2(_02775_),
    .X(_02776_));
 sky130_fd_sc_hd__o21a_1 _07762_ (.A1(net763),
    .A2(_02776_),
    .B1(_02774_),
    .X(_02777_));
 sky130_fd_sc_hd__and2b_1 _07763_ (.A_N(_02773_),
    .B(_02777_),
    .X(_02778_));
 sky130_fd_sc_hd__nand2b_1 _07764_ (.A_N(_02777_),
    .B(_02773_),
    .Y(_02779_));
 sky130_fd_sc_hd__and2_1 _07765_ (.A(_02773_),
    .B(_02777_),
    .X(_02780_));
 sky130_fd_sc_hd__nand2_1 _07766_ (.A(_02773_),
    .B(_02777_),
    .Y(_02781_));
 sky130_fd_sc_hd__or2_2 _07767_ (.A(_02773_),
    .B(_02777_),
    .X(_02782_));
 sky130_fd_sc_hd__nand2_2 _07768_ (.A(_02781_),
    .B(_02782_),
    .Y(_02783_));
 sky130_fd_sc_hd__and4b_1 _07769_ (.A_N(_02766_),
    .B(_02767_),
    .C(_02781_),
    .D(_02782_),
    .X(_02784_));
 sky130_fd_sc_hd__and2b_1 _07770_ (.A_N(net981),
    .B(\rWrDataWB[26] ),
    .X(_02785_));
 sky130_fd_sc_hd__a21oi_1 _07771_ (.A1(net981),
    .A2(net20),
    .B1(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__a21o_1 _07772_ (.A1(net981),
    .A2(net20),
    .B1(_02785_),
    .X(_02787_));
 sky130_fd_sc_hd__o211ai_4 _07773_ (.A1(net598),
    .A2(net708),
    .B1(_01864_),
    .C1(net619),
    .Y(_02788_));
 sky130_fd_sc_hd__a32oi_4 _07774_ (.A1(_01848_),
    .A2(net737),
    .A3(_02788_),
    .B1(net731),
    .B2(net153),
    .Y(_02789_));
 sky130_fd_sc_hd__a32o_2 _07775_ (.A1(_01848_),
    .A2(net737),
    .A3(_02788_),
    .B1(net731),
    .B2(net153),
    .X(_02790_));
 sky130_fd_sc_hd__a31o_1 _07776_ (.A1(net949),
    .A2(\brancher.imm13_b[6] ),
    .A3(net767),
    .B1(net726),
    .X(_02791_));
 sky130_fd_sc_hd__a21o_1 _07777_ (.A1(net578),
    .A2(_02787_),
    .B1(net615),
    .X(_02792_));
 sky130_fd_sc_hd__o22a_1 _07778_ (.A1(\rWrData[26] ),
    .A2(net607),
    .B1(_02480_),
    .B2(_02792_),
    .X(_02793_));
 sky130_fd_sc_hd__o21a_2 _07779_ (.A1(net762),
    .A2(_02793_),
    .B1(_02791_),
    .X(_02794_));
 sky130_fd_sc_hd__nand2_1 _07780_ (.A(_02789_),
    .B(_02794_),
    .Y(_02795_));
 sky130_fd_sc_hd__nor2_1 _07781_ (.A(_02789_),
    .B(_02794_),
    .Y(_02796_));
 sky130_fd_sc_hd__and2_1 _07782_ (.A(_02790_),
    .B(_02794_),
    .X(_02797_));
 sky130_fd_sc_hd__xnor2_4 _07783_ (.A(_02789_),
    .B(_02794_),
    .Y(_02798_));
 sky130_fd_sc_hd__and2b_1 _07784_ (.A_N(net977),
    .B(\rWrDataWB[27] ),
    .X(_02799_));
 sky130_fd_sc_hd__a21oi_1 _07785_ (.A1(net977),
    .A2(net21),
    .B1(_02799_),
    .Y(_02800_));
 sky130_fd_sc_hd__a21o_1 _07786_ (.A1(net977),
    .A2(net21),
    .B1(_02799_),
    .X(_02801_));
 sky130_fd_sc_hd__a21o_1 _07787_ (.A1(net590),
    .A2(_02801_),
    .B1(net625),
    .X(_02802_));
 sky130_fd_sc_hd__a21oi_1 _07788_ (.A1(net598),
    .A2(_01884_),
    .B1(_02802_),
    .Y(_02803_));
 sky130_fd_sc_hd__o32a_4 _07789_ (.A1(_01868_),
    .A2(_02579_),
    .A3(_02803_),
    .B1(_02582_),
    .B2(_01205_),
    .X(_02804_));
 sky130_fd_sc_hd__a31o_1 _07790_ (.A1(net949),
    .A2(\brancher.imm13_b[7] ),
    .A3(net767),
    .B1(net726),
    .X(_02805_));
 sky130_fd_sc_hd__a21o_1 _07791_ (.A1(net578),
    .A2(_02801_),
    .B1(net612),
    .X(_02806_));
 sky130_fd_sc_hd__o22a_1 _07792_ (.A1(\rWrData[27] ),
    .A2(net606),
    .B1(_02498_),
    .B2(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__o21a_2 _07793_ (.A1(net762),
    .A2(_02807_),
    .B1(_02805_),
    .X(_02808_));
 sky130_fd_sc_hd__nand2b_1 _07794_ (.A_N(_02804_),
    .B(_02808_),
    .Y(_02809_));
 sky130_fd_sc_hd__nand2b_1 _07795_ (.A_N(_02808_),
    .B(_02804_),
    .Y(_02810_));
 sky130_fd_sc_hd__nor2_1 _07796_ (.A(_02804_),
    .B(_02808_),
    .Y(_02811_));
 sky130_fd_sc_hd__nand2_1 _07797_ (.A(_02804_),
    .B(_02808_),
    .Y(_02812_));
 sky130_fd_sc_hd__xnor2_2 _07798_ (.A(_02804_),
    .B(_02808_),
    .Y(_02813_));
 sky130_fd_sc_hd__nor2_1 _07799_ (.A(_02798_),
    .B(_02813_),
    .Y(_02814_));
 sky130_fd_sc_hd__and2b_1 _07800_ (.A_N(net981),
    .B(\rWrDataWB[25] ),
    .X(_02815_));
 sky130_fd_sc_hd__a21oi_1 _07801_ (.A1(net977),
    .A2(net19),
    .B1(_02815_),
    .Y(_02816_));
 sky130_fd_sc_hd__a21o_1 _07802_ (.A1(net978),
    .A2(net19),
    .B1(_02815_),
    .X(_02817_));
 sky130_fd_sc_hd__a21oi_1 _07803_ (.A1(net592),
    .A2(_02817_),
    .B1(net627),
    .Y(_02818_));
 sky130_fd_sc_hd__o21ai_2 _07804_ (.A1(net592),
    .A2(_01842_),
    .B1(_02818_),
    .Y(_02819_));
 sky130_fd_sc_hd__a32oi_4 _07805_ (.A1(_01826_),
    .A2(net737),
    .A3(_02819_),
    .B1(net731),
    .B2(net152),
    .Y(_02820_));
 sky130_fd_sc_hd__a32o_2 _07806_ (.A1(_01826_),
    .A2(net737),
    .A3(_02819_),
    .B1(net731),
    .B2(net152),
    .X(_02821_));
 sky130_fd_sc_hd__a31o_1 _07807_ (.A1(net949),
    .A2(\brancher.imm13_b[5] ),
    .A3(net768),
    .B1(_02590_),
    .X(_02822_));
 sky130_fd_sc_hd__a21o_1 _07808_ (.A1(net580),
    .A2(_02817_),
    .B1(net614),
    .X(_02823_));
 sky130_fd_sc_hd__o22a_1 _07809_ (.A1(\rWrData[25] ),
    .A2(net607),
    .B1(_02462_),
    .B2(_02823_),
    .X(_02824_));
 sky130_fd_sc_hd__o21a_2 _07810_ (.A1(net763),
    .A2(_02824_),
    .B1(_02822_),
    .X(_02825_));
 sky130_fd_sc_hd__or2_1 _07811_ (.A(_02821_),
    .B(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__and2_1 _07812_ (.A(_02821_),
    .B(_02825_),
    .X(_02827_));
 sky130_fd_sc_hd__nor2_1 _07813_ (.A(_02820_),
    .B(_02825_),
    .Y(_02828_));
 sky130_fd_sc_hd__xnor2_2 _07814_ (.A(_02820_),
    .B(_02825_),
    .Y(_02829_));
 sky130_fd_sc_hd__inv_2 _07815_ (.A(_02829_),
    .Y(_02830_));
 sky130_fd_sc_hd__and2b_1 _07816_ (.A_N(net978),
    .B(\rWrDataWB[24] ),
    .X(_02831_));
 sky130_fd_sc_hd__a21oi_2 _07817_ (.A1(net978),
    .A2(net18),
    .B1(_02831_),
    .Y(_02832_));
 sky130_fd_sc_hd__a21o_1 _07818_ (.A1(net978),
    .A2(net18),
    .B1(_02831_),
    .X(_02833_));
 sky130_fd_sc_hd__nor2_1 _07819_ (.A(net598),
    .B(net705),
    .Y(_02834_));
 sky130_fd_sc_hd__a211o_1 _07820_ (.A1(net598),
    .A2(_01820_),
    .B1(_02834_),
    .C1(net625),
    .X(_02835_));
 sky130_fd_sc_hd__a32oi_4 _07821_ (.A1(_01804_),
    .A2(net737),
    .A3(_02835_),
    .B1(net731),
    .B2(net151),
    .Y(_02836_));
 sky130_fd_sc_hd__a32o_2 _07822_ (.A1(_01804_),
    .A2(net737),
    .A3(_02835_),
    .B1(net731),
    .B2(net151),
    .X(_02837_));
 sky130_fd_sc_hd__a31o_1 _07823_ (.A1(net950),
    .A2(net942),
    .A3(net768),
    .B1(net726),
    .X(_02838_));
 sky130_fd_sc_hd__a21o_1 _07824_ (.A1(net582),
    .A2(_02833_),
    .B1(net615),
    .X(_02839_));
 sky130_fd_sc_hd__a31o_1 _07825_ (.A1(net586),
    .A2(_02435_),
    .A3(_02443_),
    .B1(_02839_),
    .X(_02840_));
 sky130_fd_sc_hd__a21o_2 _07826_ (.A1(_02427_),
    .A2(_02840_),
    .B1(net763),
    .X(_02841_));
 sky130_fd_sc_hd__nand3_2 _07827_ (.A(_02837_),
    .B(_02838_),
    .C(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__a21o_1 _07828_ (.A1(_02838_),
    .A2(_02841_),
    .B1(_02837_),
    .X(_02843_));
 sky130_fd_sc_hd__a21o_1 _07829_ (.A1(_02838_),
    .A2(_02841_),
    .B1(_02836_),
    .X(_02844_));
 sky130_fd_sc_hd__nand2_2 _07830_ (.A(_02842_),
    .B(_02843_),
    .Y(_02845_));
 sky130_fd_sc_hd__a21oi_1 _07831_ (.A1(_02842_),
    .A2(_02843_),
    .B1(_02829_),
    .Y(_02846_));
 sky130_fd_sc_hd__nand2_1 _07832_ (.A(_02814_),
    .B(_02846_),
    .Y(_02847_));
 sky130_fd_sc_hd__and4_1 _07833_ (.A(net183),
    .B(_02784_),
    .C(_02814_),
    .D(_02846_),
    .X(_02848_));
 sky130_fd_sc_hd__and2b_1 _07834_ (.A_N(net980),
    .B(\rWrDataWB[22] ),
    .X(_02849_));
 sky130_fd_sc_hd__a21oi_1 _07835_ (.A1(net980),
    .A2(net16),
    .B1(_02849_),
    .Y(_02850_));
 sky130_fd_sc_hd__a21o_1 _07836_ (.A1(net980),
    .A2(net16),
    .B1(_02849_),
    .X(_02851_));
 sky130_fd_sc_hd__o211ai_2 _07837_ (.A1(net600),
    .A2(net704),
    .B1(_01777_),
    .C1(net621),
    .Y(_02852_));
 sky130_fd_sc_hd__a32oi_4 _07838_ (.A1(_01761_),
    .A2(net737),
    .A3(_02852_),
    .B1(net731),
    .B2(net149),
    .Y(_02853_));
 sky130_fd_sc_hd__a32o_2 _07839_ (.A1(_01761_),
    .A2(net737),
    .A3(_02852_),
    .B1(net731),
    .B2(net149),
    .X(_02854_));
 sky130_fd_sc_hd__a31o_1 _07840_ (.A1(net949),
    .A2(net864),
    .A3(net767),
    .B1(net726),
    .X(_02855_));
 sky130_fd_sc_hd__a21o_1 _07841_ (.A1(net580),
    .A2(_02851_),
    .B1(net614),
    .X(_02856_));
 sky130_fd_sc_hd__o22a_1 _07842_ (.A1(\rWrData[22] ),
    .A2(net607),
    .B1(_02407_),
    .B2(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__o21a_2 _07843_ (.A1(net762),
    .A2(_02857_),
    .B1(_02855_),
    .X(_02858_));
 sky130_fd_sc_hd__and2_1 _07844_ (.A(_02854_),
    .B(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__nand2_1 _07845_ (.A(_02853_),
    .B(_02858_),
    .Y(_02860_));
 sky130_fd_sc_hd__nor2_1 _07846_ (.A(_02853_),
    .B(_02858_),
    .Y(_02861_));
 sky130_fd_sc_hd__xnor2_4 _07847_ (.A(_02853_),
    .B(_02858_),
    .Y(_02862_));
 sky130_fd_sc_hd__and2b_1 _07848_ (.A_N(net977),
    .B(\rWrDataWB[23] ),
    .X(_02863_));
 sky130_fd_sc_hd__a21oi_1 _07849_ (.A1(net977),
    .A2(net17),
    .B1(_02863_),
    .Y(_02864_));
 sky130_fd_sc_hd__a21o_2 _07850_ (.A1(net977),
    .A2(net17),
    .B1(_02863_),
    .X(_02865_));
 sky130_fd_sc_hd__a21oi_1 _07851_ (.A1(net590),
    .A2(_02865_),
    .B1(net625),
    .Y(_02866_));
 sky130_fd_sc_hd__o21ai_2 _07852_ (.A1(net590),
    .A2(_01798_),
    .B1(_02866_),
    .Y(_02867_));
 sky130_fd_sc_hd__a32oi_4 _07853_ (.A1(_01782_),
    .A2(net737),
    .A3(_02867_),
    .B1(net731),
    .B2(net150),
    .Y(_02868_));
 sky130_fd_sc_hd__a32o_2 _07854_ (.A1(_01782_),
    .A2(net737),
    .A3(_02867_),
    .B1(net731),
    .B2(net150),
    .X(_02869_));
 sky130_fd_sc_hd__a31o_1 _07855_ (.A1(net949),
    .A2(net855),
    .A3(net768),
    .B1(net726),
    .X(_02870_));
 sky130_fd_sc_hd__a21o_1 _07856_ (.A1(net578),
    .A2(_02865_),
    .B1(net612),
    .X(_02871_));
 sky130_fd_sc_hd__o22a_1 _07857_ (.A1(\rWrData[23] ),
    .A2(net606),
    .B1(_02425_),
    .B2(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__o21a_2 _07858_ (.A1(net762),
    .A2(_02872_),
    .B1(_02870_),
    .X(_02873_));
 sky130_fd_sc_hd__and2_1 _07859_ (.A(_02869_),
    .B(_02873_),
    .X(_02874_));
 sky130_fd_sc_hd__nor2_1 _07860_ (.A(_02869_),
    .B(_02873_),
    .Y(_02875_));
 sky130_fd_sc_hd__nand2_1 _07861_ (.A(_02868_),
    .B(_02873_),
    .Y(_02876_));
 sky130_fd_sc_hd__nor2_1 _07862_ (.A(_02868_),
    .B(_02873_),
    .Y(_02877_));
 sky130_fd_sc_hd__xnor2_4 _07863_ (.A(_02868_),
    .B(_02873_),
    .Y(_02878_));
 sky130_fd_sc_hd__or2_1 _07864_ (.A(_02862_),
    .B(_02878_),
    .X(_02879_));
 sky130_fd_sc_hd__and2b_1 _07865_ (.A_N(net979),
    .B(\rWrDataWB[20] ),
    .X(_02880_));
 sky130_fd_sc_hd__a21oi_1 _07866_ (.A1(net976),
    .A2(net14),
    .B1(_02880_),
    .Y(_02881_));
 sky130_fd_sc_hd__a21o_1 _07867_ (.A1(net979),
    .A2(net14),
    .B1(_02880_),
    .X(_02882_));
 sky130_fd_sc_hd__a211o_2 _07868_ (.A1(net593),
    .A2(_02882_),
    .B1(_01733_),
    .C1(net626),
    .X(_02883_));
 sky130_fd_sc_hd__a32oi_4 _07869_ (.A1(_01715_),
    .A2(net738),
    .A3(_02883_),
    .B1(net732),
    .B2(net147),
    .Y(_02884_));
 sky130_fd_sc_hd__a32o_2 _07870_ (.A1(_01715_),
    .A2(net738),
    .A3(_02883_),
    .B1(net732),
    .B2(net147),
    .X(_02885_));
 sky130_fd_sc_hd__a31o_1 _07871_ (.A1(net948),
    .A2(net936),
    .A3(net766),
    .B1(net727),
    .X(_02886_));
 sky130_fd_sc_hd__a21o_1 _07872_ (.A1(net579),
    .A2(_02882_),
    .B1(net613),
    .X(_02887_));
 sky130_fd_sc_hd__o22a_1 _07873_ (.A1(\rWrData[20] ),
    .A2(net605),
    .B1(_02371_),
    .B2(_02887_),
    .X(_02888_));
 sky130_fd_sc_hd__o21a_2 _07874_ (.A1(net761),
    .A2(_02888_),
    .B1(_02886_),
    .X(_02889_));
 sky130_fd_sc_hd__and2_1 _07875_ (.A(_02885_),
    .B(_02889_),
    .X(_02890_));
 sky130_fd_sc_hd__nor2_1 _07876_ (.A(_02884_),
    .B(_02889_),
    .Y(_02891_));
 sky130_fd_sc_hd__xnor2_4 _07877_ (.A(_02884_),
    .B(_02889_),
    .Y(_02892_));
 sky130_fd_sc_hd__and2b_1 _07878_ (.A_N(net980),
    .B(\rWrDataWB[21] ),
    .X(_02893_));
 sky130_fd_sc_hd__a21oi_2 _07879_ (.A1(net981),
    .A2(net15),
    .B1(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__a21o_1 _07880_ (.A1(net981),
    .A2(net15),
    .B1(_02893_),
    .X(_02895_));
 sky130_fd_sc_hd__o211ai_2 _07881_ (.A1(net600),
    .A2(net701),
    .B1(_01755_),
    .C1(net620),
    .Y(_02896_));
 sky130_fd_sc_hd__a32oi_4 _07882_ (.A1(_01738_),
    .A2(net739),
    .A3(_02896_),
    .B1(net733),
    .B2(net148),
    .Y(_02897_));
 sky130_fd_sc_hd__a32o_2 _07883_ (.A1(_01738_),
    .A2(net739),
    .A3(_02896_),
    .B1(net733),
    .B2(net148),
    .X(_02898_));
 sky130_fd_sc_hd__a31o_1 _07884_ (.A1(net949),
    .A2(net900),
    .A3(net769),
    .B1(net726),
    .X(_02899_));
 sky130_fd_sc_hd__a21oi_1 _07885_ (.A1(net581),
    .A2(_02895_),
    .B1(net614),
    .Y(_02900_));
 sky130_fd_sc_hd__o2bb2a_1 _07886_ (.A1_N(_02900_),
    .A2_N(_02389_),
    .B1(net607),
    .B2(\rWrData[21] ),
    .X(_02901_));
 sky130_fd_sc_hd__o21a_2 _07887_ (.A1(net762),
    .A2(_02901_),
    .B1(_02899_),
    .X(_02902_));
 sky130_fd_sc_hd__nor2_1 _07888_ (.A(_02897_),
    .B(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__xnor2_4 _07889_ (.A(_02897_),
    .B(_02902_),
    .Y(_02904_));
 sky130_fd_sc_hd__inv_2 _07890_ (.A(_02904_),
    .Y(_02905_));
 sky130_fd_sc_hd__nor4_1 _07891_ (.A(_02862_),
    .B(_02878_),
    .C(_02892_),
    .D(_02904_),
    .Y(_02906_));
 sky130_fd_sc_hd__or4_1 _07892_ (.A(_02862_),
    .B(_02878_),
    .C(_02892_),
    .D(_02904_),
    .X(_02907_));
 sky130_fd_sc_hd__and2b_1 _07893_ (.A_N(net976),
    .B(\rWrDataWB[18] ),
    .X(_02908_));
 sky130_fd_sc_hd__a21oi_2 _07894_ (.A1(net976),
    .A2(net11),
    .B1(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__a21o_1 _07895_ (.A1(net976),
    .A2(net11),
    .B1(_02908_),
    .X(_02910_));
 sky130_fd_sc_hd__nor2_1 _07896_ (.A(net599),
    .B(_02909_),
    .Y(_02911_));
 sky130_fd_sc_hd__a211o_1 _07897_ (.A1(net599),
    .A2(_01689_),
    .B1(_02911_),
    .C1(net626),
    .X(_02912_));
 sky130_fd_sc_hd__a32oi_2 _07898_ (.A1(_01673_),
    .A2(net738),
    .A3(_02912_),
    .B1(net729),
    .B2(net144),
    .Y(_02913_));
 sky130_fd_sc_hd__a32o_2 _07899_ (.A1(_01673_),
    .A2(net738),
    .A3(_02912_),
    .B1(net729),
    .B2(net144),
    .X(_02914_));
 sky130_fd_sc_hd__a31o_1 _07900_ (.A1(net950),
    .A2(net990),
    .A3(net768),
    .B1(net727),
    .X(_02915_));
 sky130_fd_sc_hd__a21oi_1 _07901_ (.A1(net579),
    .A2(_02910_),
    .B1(net613),
    .Y(_02916_));
 sky130_fd_sc_hd__o2bb2a_2 _07902_ (.A1_N(_02916_),
    .A2_N(_02335_),
    .B1(net605),
    .B2(\rWrData[18] ),
    .X(_02917_));
 sky130_fd_sc_hd__o21ai_2 _07903_ (.A1(net760),
    .A2(_02917_),
    .B1(_02915_),
    .Y(_02918_));
 sky130_fd_sc_hd__nor2_1 _07904_ (.A(_02913_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__nand2_1 _07905_ (.A(_02913_),
    .B(_02918_),
    .Y(_02920_));
 sky130_fd_sc_hd__xnor2_2 _07906_ (.A(_02914_),
    .B(_02918_),
    .Y(_02921_));
 sky130_fd_sc_hd__and2b_1 _07907_ (.A_N(net976),
    .B(\rWrDataWB[19] ),
    .X(_02922_));
 sky130_fd_sc_hd__a21oi_2 _07908_ (.A1(net976),
    .A2(net12),
    .B1(_02922_),
    .Y(_02923_));
 sky130_fd_sc_hd__a21o_1 _07909_ (.A1(net976),
    .A2(net12),
    .B1(_02922_),
    .X(_02924_));
 sky130_fd_sc_hd__o211a_1 _07910_ (.A1(net599),
    .A2(_02923_),
    .B1(_01710_),
    .C1(net621),
    .X(_02925_));
 sky130_fd_sc_hd__o32a_4 _07911_ (.A1(_01694_),
    .A2(_02579_),
    .A3(_02925_),
    .B1(_02582_),
    .B2(_01206_),
    .X(_02926_));
 sky130_fd_sc_hd__a31o_1 _07912_ (.A1(net950),
    .A2(net1069),
    .A3(net768),
    .B1(net726),
    .X(_02927_));
 sky130_fd_sc_hd__a21oi_1 _07913_ (.A1(net579),
    .A2(_02924_),
    .B1(net613),
    .Y(_02928_));
 sky130_fd_sc_hd__o2bb2a_1 _07914_ (.A1_N(_02928_),
    .A2_N(_02353_),
    .B1(net605),
    .B2(\rWrData[19] ),
    .X(_02929_));
 sky130_fd_sc_hd__o21a_2 _07915_ (.A1(net762),
    .A2(_02929_),
    .B1(_02927_),
    .X(_02930_));
 sky130_fd_sc_hd__and2b_1 _07916_ (.A_N(_02926_),
    .B(_02930_),
    .X(_02931_));
 sky130_fd_sc_hd__and2b_1 _07917_ (.A_N(_02930_),
    .B(_02926_),
    .X(_02932_));
 sky130_fd_sc_hd__nand2_1 _07918_ (.A(_02926_),
    .B(_02930_),
    .Y(_02933_));
 sky130_fd_sc_hd__nor2_1 _07919_ (.A(_02926_),
    .B(_02930_),
    .Y(_02934_));
 sky130_fd_sc_hd__xnor2_2 _07920_ (.A(_02926_),
    .B(_02930_),
    .Y(_02935_));
 sky130_fd_sc_hd__nor2_1 _07921_ (.A(_02921_),
    .B(_02935_),
    .Y(_02936_));
 sky130_fd_sc_hd__and2b_1 _07922_ (.A_N(net980),
    .B(\rWrDataWB[16] ),
    .X(_02937_));
 sky130_fd_sc_hd__a21oi_2 _07923_ (.A1(net980),
    .A2(net9),
    .B1(_02937_),
    .Y(_02938_));
 sky130_fd_sc_hd__a21o_1 _07924_ (.A1(net980),
    .A2(net9),
    .B1(_02937_),
    .X(_02939_));
 sky130_fd_sc_hd__o211ai_4 _07925_ (.A1(net600),
    .A2(net698),
    .B1(_01645_),
    .C1(net620),
    .Y(_02940_));
 sky130_fd_sc_hd__a32oi_4 _07926_ (.A1(_01629_),
    .A2(net736),
    .A3(_02940_),
    .B1(net730),
    .B2(net142),
    .Y(_02941_));
 sky130_fd_sc_hd__a32o_1 _07927_ (.A1(_01629_),
    .A2(net736),
    .A3(_02940_),
    .B1(net730),
    .B2(net142),
    .X(_02942_));
 sky130_fd_sc_hd__a31o_1 _07928_ (.A1(net948),
    .A2(net1030),
    .A3(net770),
    .B1(net727),
    .X(_02943_));
 sky130_fd_sc_hd__a21o_1 _07929_ (.A1(net581),
    .A2(_02939_),
    .B1(net614),
    .X(_02944_));
 sky130_fd_sc_hd__a31o_1 _07930_ (.A1(net586),
    .A2(_02290_),
    .A3(_02298_),
    .B1(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__a21o_1 _07931_ (.A1(_02282_),
    .A2(_02945_),
    .B1(net763),
    .X(_02946_));
 sky130_fd_sc_hd__and3_1 _07932_ (.A(_02941_),
    .B(_02943_),
    .C(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__a21oi_1 _07933_ (.A1(_02943_),
    .A2(_02946_),
    .B1(_02941_),
    .Y(_02948_));
 sky130_fd_sc_hd__nor2_1 _07934_ (.A(_02947_),
    .B(_02948_),
    .Y(_02949_));
 sky130_fd_sc_hd__and2b_1 _07935_ (.A_N(net976),
    .B(\rWrDataWB[17] ),
    .X(_02950_));
 sky130_fd_sc_hd__a21oi_1 _07936_ (.A1(net976),
    .A2(net10),
    .B1(_02950_),
    .Y(_02951_));
 sky130_fd_sc_hd__a21o_2 _07937_ (.A1(net976),
    .A2(net10),
    .B1(_02950_),
    .X(_02952_));
 sky130_fd_sc_hd__a21oi_1 _07938_ (.A1(net593),
    .A2(_02952_),
    .B1(net626),
    .Y(_02953_));
 sky130_fd_sc_hd__o21ai_2 _07939_ (.A1(net593),
    .A2(_01666_),
    .B1(_02953_),
    .Y(_02954_));
 sky130_fd_sc_hd__a32oi_4 _07940_ (.A1(_01650_),
    .A2(net738),
    .A3(_02954_),
    .B1(net732),
    .B2(net143),
    .Y(_02955_));
 sky130_fd_sc_hd__a32o_4 _07941_ (.A1(_01650_),
    .A2(net738),
    .A3(_02954_),
    .B1(net732),
    .B2(net143),
    .X(_02956_));
 sky130_fd_sc_hd__a31o_1 _07942_ (.A1(net950),
    .A2(net997),
    .A3(net768),
    .B1(net727),
    .X(_02957_));
 sky130_fd_sc_hd__a21o_1 _07943_ (.A1(net579),
    .A2(_02952_),
    .B1(net613),
    .X(_02958_));
 sky130_fd_sc_hd__o22a_1 _07944_ (.A1(\rWrData[17] ),
    .A2(net605),
    .B1(_02317_),
    .B2(_02958_),
    .X(_02959_));
 sky130_fd_sc_hd__o21a_2 _07945_ (.A1(net762),
    .A2(_02959_),
    .B1(_02957_),
    .X(_02960_));
 sky130_fd_sc_hd__and2_1 _07946_ (.A(_02956_),
    .B(_02960_),
    .X(_02961_));
 sky130_fd_sc_hd__or2_1 _07947_ (.A(_02956_),
    .B(_02960_),
    .X(_02962_));
 sky130_fd_sc_hd__nor2_1 _07948_ (.A(_02955_),
    .B(_02960_),
    .Y(_02963_));
 sky130_fd_sc_hd__xnor2_4 _07949_ (.A(_02956_),
    .B(_02960_),
    .Y(_02964_));
 sky130_fd_sc_hd__and3_1 _07950_ (.A(_02936_),
    .B(net181),
    .C(_02964_),
    .X(_02965_));
 sky130_fd_sc_hd__and4_1 _07951_ (.A(_02906_),
    .B(_02936_),
    .C(net181),
    .D(_02964_),
    .X(_02966_));
 sky130_fd_sc_hd__nand2_1 _07952_ (.A(_02848_),
    .B(_02966_),
    .Y(_02967_));
 sky130_fd_sc_hd__and2b_1 _07953_ (.A_N(net982),
    .B(\rWrDataWB[14] ),
    .X(_02968_));
 sky130_fd_sc_hd__a21oi_2 _07954_ (.A1(net982),
    .A2(net7),
    .B1(_02968_),
    .Y(_02969_));
 sky130_fd_sc_hd__a21o_1 _07955_ (.A1(net982),
    .A2(net7),
    .B1(_02968_),
    .X(_02970_));
 sky130_fd_sc_hd__o211ai_2 _07956_ (.A1(net599),
    .A2(net696),
    .B1(_01603_),
    .C1(net618),
    .Y(_02971_));
 sky130_fd_sc_hd__a32oi_4 _07957_ (.A1(_01585_),
    .A2(net735),
    .A3(_02971_),
    .B1(net729),
    .B2(net140),
    .Y(_02972_));
 sky130_fd_sc_hd__a32o_2 _07958_ (.A1(_01585_),
    .A2(net735),
    .A3(_02971_),
    .B1(net729),
    .B2(net140),
    .X(_02973_));
 sky130_fd_sc_hd__a31o_1 _07959_ (.A1(net948),
    .A2(net943),
    .A3(net766),
    .B1(net727),
    .X(_02974_));
 sky130_fd_sc_hd__a21o_1 _07960_ (.A1(net577),
    .A2(_02970_),
    .B1(net611),
    .X(_02975_));
 sky130_fd_sc_hd__o22a_1 _07961_ (.A1(\rWrData[14] ),
    .A2(net603),
    .B1(_02262_),
    .B2(_02975_),
    .X(_02976_));
 sky130_fd_sc_hd__o21a_1 _07962_ (.A1(net760),
    .A2(_02976_),
    .B1(_02974_),
    .X(_02977_));
 sky130_fd_sc_hd__and2_1 _07963_ (.A(_02972_),
    .B(_02977_),
    .X(_02978_));
 sky130_fd_sc_hd__nand2_1 _07964_ (.A(_02972_),
    .B(_02977_),
    .Y(_02979_));
 sky130_fd_sc_hd__nor2_1 _07965_ (.A(_02972_),
    .B(_02977_),
    .Y(_02980_));
 sky130_fd_sc_hd__nor2_1 _07966_ (.A(_02978_),
    .B(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__xnor2_2 _07967_ (.A(_02972_),
    .B(_02977_),
    .Y(_02982_));
 sky130_fd_sc_hd__and2b_1 _07968_ (.A_N(net982),
    .B(\rWrDataWB[15] ),
    .X(_02983_));
 sky130_fd_sc_hd__a21oi_2 _07969_ (.A1(net982),
    .A2(net8),
    .B1(_02983_),
    .Y(_02984_));
 sky130_fd_sc_hd__a21o_1 _07970_ (.A1(net982),
    .A2(net8),
    .B1(_02983_),
    .X(_02985_));
 sky130_fd_sc_hd__nor2_1 _07971_ (.A(net599),
    .B(_02984_),
    .Y(_02986_));
 sky130_fd_sc_hd__a211o_1 _07972_ (.A1(net599),
    .A2(_01624_),
    .B1(_02986_),
    .C1(net626),
    .X(_02987_));
 sky130_fd_sc_hd__a32oi_4 _07973_ (.A1(_01608_),
    .A2(net735),
    .A3(_02987_),
    .B1(net729),
    .B2(net141),
    .Y(_02988_));
 sky130_fd_sc_hd__a31o_1 _07974_ (.A1(net948),
    .A2(net1064),
    .A3(net766),
    .B1(net727),
    .X(_02989_));
 sky130_fd_sc_hd__a21o_1 _07975_ (.A1(net579),
    .A2(_02985_),
    .B1(net613),
    .X(_02990_));
 sky130_fd_sc_hd__o22a_1 _07976_ (.A1(\rWrData[15] ),
    .A2(net605),
    .B1(_02280_),
    .B2(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__o21a_2 _07977_ (.A1(net760),
    .A2(_02991_),
    .B1(_02989_),
    .X(_02992_));
 sky130_fd_sc_hd__nand2b_1 _07978_ (.A_N(_02992_),
    .B(net205),
    .Y(_02993_));
 sky130_fd_sc_hd__and2b_1 _07979_ (.A_N(net205),
    .B(_02992_),
    .X(_02994_));
 sky130_fd_sc_hd__nand2_1 _07980_ (.A(net205),
    .B(_02992_),
    .Y(_02995_));
 sky130_fd_sc_hd__nor2_1 _07981_ (.A(net205),
    .B(_02992_),
    .Y(_02996_));
 sky130_fd_sc_hd__xnor2_4 _07982_ (.A(_02988_),
    .B(_02992_),
    .Y(_02997_));
 sky130_fd_sc_hd__nor2_1 _07983_ (.A(_02982_),
    .B(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__and2b_1 _07984_ (.A_N(net972),
    .B(\rWrDataWB[13] ),
    .X(_02999_));
 sky130_fd_sc_hd__a21oi_2 _07985_ (.A1(net972),
    .A2(net6),
    .B1(_02999_),
    .Y(_03000_));
 sky130_fd_sc_hd__a21o_1 _07986_ (.A1(net972),
    .A2(net6),
    .B1(_02999_),
    .X(_03001_));
 sky130_fd_sc_hd__nor2_1 _07987_ (.A(net596),
    .B(_03000_),
    .Y(_03002_));
 sky130_fd_sc_hd__a211o_1 _07988_ (.A1(net596),
    .A2(_01580_),
    .B1(_03002_),
    .C1(net622),
    .X(_03003_));
 sky130_fd_sc_hd__a32o_4 _07989_ (.A1(_01564_),
    .A2(net734),
    .A3(_03003_),
    .B1(net728),
    .B2(net139),
    .X(_03004_));
 sky130_fd_sc_hd__inv_2 _07990_ (.A(_03004_),
    .Y(_03005_));
 sky130_fd_sc_hd__a31o_1 _07991_ (.A1(net948),
    .A2(net845),
    .A3(net770),
    .B1(net727),
    .X(_03006_));
 sky130_fd_sc_hd__a21o_1 _07992_ (.A1(net576),
    .A2(_03001_),
    .B1(net609),
    .X(_03007_));
 sky130_fd_sc_hd__o22a_2 _07993_ (.A1(\rWrData[13] ),
    .A2(net604),
    .B1(_02244_),
    .B2(_03007_),
    .X(_03008_));
 sky130_fd_sc_hd__o21ai_4 _07994_ (.A1(net760),
    .A2(_03008_),
    .B1(_03006_),
    .Y(_03009_));
 sky130_fd_sc_hd__and2_1 _07995_ (.A(_03004_),
    .B(_03009_),
    .X(_03010_));
 sky130_fd_sc_hd__or2_1 _07996_ (.A(_03004_),
    .B(_03009_),
    .X(_03011_));
 sky130_fd_sc_hd__xor2_2 _07997_ (.A(_03004_),
    .B(_03009_),
    .X(_03012_));
 sky130_fd_sc_hd__and2b_1 _07998_ (.A_N(net972),
    .B(\rWrDataWB[12] ),
    .X(_03013_));
 sky130_fd_sc_hd__a21oi_2 _07999_ (.A1(net972),
    .A2(net5),
    .B1(_03013_),
    .Y(_03014_));
 sky130_fd_sc_hd__a21o_1 _08000_ (.A1(net972),
    .A2(net5),
    .B1(_03013_),
    .X(_03015_));
 sky130_fd_sc_hd__nor2_1 _08001_ (.A(net596),
    .B(_03014_),
    .Y(_03016_));
 sky130_fd_sc_hd__a211o_1 _08002_ (.A1(net596),
    .A2(_01558_),
    .B1(_03016_),
    .C1(net623),
    .X(_03017_));
 sky130_fd_sc_hd__a32o_4 _08003_ (.A1(_01542_),
    .A2(net735),
    .A3(_03017_),
    .B1(net729),
    .B2(net138),
    .X(_03018_));
 sky130_fd_sc_hd__a31o_1 _08004_ (.A1(net948),
    .A2(net847),
    .A3(net766),
    .B1(net727),
    .X(_03019_));
 sky130_fd_sc_hd__a21o_1 _08005_ (.A1(net576),
    .A2(_03015_),
    .B1(net611),
    .X(_03020_));
 sky130_fd_sc_hd__a31o_1 _08006_ (.A1(net584),
    .A2(_02217_),
    .A3(_02225_),
    .B1(_03020_),
    .X(_03021_));
 sky130_fd_sc_hd__a21o_1 _08007_ (.A1(_02209_),
    .A2(_03021_),
    .B1(net761),
    .X(_03022_));
 sky130_fd_sc_hd__nand2_1 _08008_ (.A(_03019_),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__a21oi_2 _08009_ (.A1(_03019_),
    .A2(_03022_),
    .B1(_03018_),
    .Y(_03024_));
 sky130_fd_sc_hd__and3_1 _08010_ (.A(_03018_),
    .B(_03019_),
    .C(_03022_),
    .X(_03025_));
 sky130_fd_sc_hd__nor2_2 _08011_ (.A(_03024_),
    .B(_03025_),
    .Y(_03026_));
 sky130_fd_sc_hd__o21ai_1 _08012_ (.A1(_03024_),
    .A2(_03025_),
    .B1(_03012_),
    .Y(_03027_));
 sky130_fd_sc_hd__or4b_1 _08013_ (.A(_02982_),
    .B(_02997_),
    .C(_03026_),
    .D_N(_03012_),
    .X(_03028_));
 sky130_fd_sc_hd__and2b_1 _08014_ (.A_N(net971),
    .B(\rWrDataWB[10] ),
    .X(_03029_));
 sky130_fd_sc_hd__a21oi_1 _08015_ (.A1(net971),
    .A2(net3),
    .B1(_03029_),
    .Y(_03030_));
 sky130_fd_sc_hd__a21o_2 _08016_ (.A1(net971),
    .A2(net3),
    .B1(_03029_),
    .X(_03031_));
 sky130_fd_sc_hd__nand2_1 _08017_ (.A(net588),
    .B(_03031_),
    .Y(_03032_));
 sky130_fd_sc_hd__o211a_1 _08018_ (.A1(net588),
    .A2(_01509_),
    .B1(_03032_),
    .C1(net616),
    .X(_03033_));
 sky130_fd_sc_hd__o21ai_1 _08019_ (.A1(\rWrData[10] ),
    .A2(net616),
    .B1(net734),
    .Y(_03034_));
 sky130_fd_sc_hd__a2bb2o_4 _08020_ (.A1_N(_03033_),
    .A2_N(_03034_),
    .B1(net136),
    .B2(net728),
    .X(_03035_));
 sky130_fd_sc_hd__a21o_1 _08021_ (.A1(net575),
    .A2(_03031_),
    .B1(net609),
    .X(_03036_));
 sky130_fd_sc_hd__o22ai_4 _08022_ (.A1(\rWrData[10] ),
    .A2(net601),
    .B1(_02189_),
    .B2(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__and2_1 _08023_ (.A(net759),
    .B(_03037_),
    .X(_03038_));
 sky130_fd_sc_hd__a21oi_2 _08024_ (.A1(\brancher.imm12_i_s[10] ),
    .A2(net764),
    .B1(net759),
    .Y(_03039_));
 sky130_fd_sc_hd__a21oi_4 _08025_ (.A1(net759),
    .A2(_03037_),
    .B1(_03039_),
    .Y(_03040_));
 sky130_fd_sc_hd__and2_1 _08026_ (.A(_03035_),
    .B(_03040_),
    .X(_03041_));
 sky130_fd_sc_hd__xor2_4 _08027_ (.A(_03035_),
    .B(_03040_),
    .X(_03042_));
 sky130_fd_sc_hd__and2b_1 _08028_ (.A_N(net983),
    .B(\rWrDataWB[11] ),
    .X(_03043_));
 sky130_fd_sc_hd__a21oi_2 _08029_ (.A1(net972),
    .A2(net4),
    .B1(_03043_),
    .Y(_03044_));
 sky130_fd_sc_hd__a21o_1 _08030_ (.A1(net983),
    .A2(net4),
    .B1(_03043_),
    .X(_03045_));
 sky130_fd_sc_hd__nor2_1 _08031_ (.A(net596),
    .B(_03044_),
    .Y(_03046_));
 sky130_fd_sc_hd__a211o_1 _08032_ (.A1(net596),
    .A2(_01534_),
    .B1(_03046_),
    .C1(net622),
    .X(_03047_));
 sky130_fd_sc_hd__a32oi_4 _08033_ (.A1(_01518_),
    .A2(net735),
    .A3(_03047_),
    .B1(net728),
    .B2(net137),
    .Y(_03048_));
 sky130_fd_sc_hd__a32o_2 _08034_ (.A1(_01518_),
    .A2(net734),
    .A3(_03047_),
    .B1(net728),
    .B2(net137),
    .X(_03049_));
 sky130_fd_sc_hd__a21o_1 _08035_ (.A1(net576),
    .A2(_03045_),
    .B1(net609),
    .X(_03050_));
 sky130_fd_sc_hd__o22a_1 _08036_ (.A1(\rWrData[11] ),
    .A2(net601),
    .B1(_02207_),
    .B2(_03050_),
    .X(_03051_));
 sky130_fd_sc_hd__o21a_1 _08037_ (.A1(net761),
    .A2(_03051_),
    .B1(net727),
    .X(_03052_));
 sky130_fd_sc_hd__nand2_1 _08038_ (.A(_03049_),
    .B(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__or2_1 _08039_ (.A(_03049_),
    .B(_03052_),
    .X(_03054_));
 sky130_fd_sc_hd__nor2_1 _08040_ (.A(_03048_),
    .B(_03052_),
    .Y(_03055_));
 sky130_fd_sc_hd__nand2_1 _08041_ (.A(_03048_),
    .B(_03052_),
    .Y(_03056_));
 sky130_fd_sc_hd__xnor2_2 _08042_ (.A(_03048_),
    .B(_03052_),
    .Y(_03057_));
 sky130_fd_sc_hd__inv_2 _08043_ (.A(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__or2_1 _08044_ (.A(_03042_),
    .B(_03057_),
    .X(_03059_));
 sky130_fd_sc_hd__and2b_1 _08045_ (.A_N(net971),
    .B(\rWrDataWB[9] ),
    .X(_03060_));
 sky130_fd_sc_hd__a21oi_1 _08046_ (.A1(net971),
    .A2(net33),
    .B1(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__a21o_2 _08047_ (.A1(net972),
    .A2(net33),
    .B1(_03060_),
    .X(_03062_));
 sky130_fd_sc_hd__a21oi_1 _08048_ (.A1(net588),
    .A2(_03062_),
    .B1(net622),
    .Y(_03063_));
 sky130_fd_sc_hd__o21ai_2 _08049_ (.A1(net587),
    .A2(_01485_),
    .B1(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__a32oi_4 _08050_ (.A1(_01469_),
    .A2(net734),
    .A3(_03064_),
    .B1(net728),
    .B2(net166),
    .Y(_03065_));
 sky130_fd_sc_hd__a32o_4 _08051_ (.A1(_01469_),
    .A2(net734),
    .A3(_03064_),
    .B1(net728),
    .B2(net166),
    .X(_03066_));
 sky130_fd_sc_hd__a21o_1 _08052_ (.A1(net575),
    .A2(_03062_),
    .B1(net609),
    .X(_03067_));
 sky130_fd_sc_hd__o22a_1 _08053_ (.A1(\rWrData[9] ),
    .A2(net601),
    .B1(_02171_),
    .B2(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__a21o_1 _08054_ (.A1(\brancher.imm12_i_s[9] ),
    .A2(net764),
    .B1(net759),
    .X(_03069_));
 sky130_fd_sc_hd__o21a_2 _08055_ (.A1(net760),
    .A2(_03068_),
    .B1(_03069_),
    .X(_03070_));
 sky130_fd_sc_hd__nor2_1 _08056_ (.A(_03065_),
    .B(_03070_),
    .Y(_03071_));
 sky130_fd_sc_hd__nand2_1 _08057_ (.A(_03066_),
    .B(_03070_),
    .Y(_03072_));
 sky130_fd_sc_hd__or2_1 _08058_ (.A(_03066_),
    .B(_03070_),
    .X(_03073_));
 sky130_fd_sc_hd__xnor2_2 _08059_ (.A(_03066_),
    .B(_03070_),
    .Y(_03074_));
 sky130_fd_sc_hd__and2_1 _08060_ (.A(_03072_),
    .B(_03073_),
    .X(_03075_));
 sky130_fd_sc_hd__and2b_1 _08061_ (.A_N(net973),
    .B(\rWrDataWB[8] ),
    .X(_03076_));
 sky130_fd_sc_hd__a21oi_1 _08062_ (.A1(net974),
    .A2(net32),
    .B1(_03076_),
    .Y(_03077_));
 sky130_fd_sc_hd__a21o_1 _08063_ (.A1(net974),
    .A2(net32),
    .B1(_03076_),
    .X(_03078_));
 sky130_fd_sc_hd__a211o_1 _08064_ (.A1(net589),
    .A2(_03078_),
    .B1(_01461_),
    .C1(net624),
    .X(_03079_));
 sky130_fd_sc_hd__a32oi_4 _08065_ (.A1(_01446_),
    .A2(net734),
    .A3(_03079_),
    .B1(net728),
    .B2(net165),
    .Y(_03080_));
 sky130_fd_sc_hd__a32o_2 _08066_ (.A1(_01446_),
    .A2(net734),
    .A3(_03079_),
    .B1(net729),
    .B2(net165),
    .X(_03081_));
 sky130_fd_sc_hd__a21o_1 _08067_ (.A1(net577),
    .A2(_03078_),
    .B1(net610),
    .X(_03082_));
 sky130_fd_sc_hd__o22a_1 _08068_ (.A1(\rWrData[8] ),
    .A2(net602),
    .B1(_02153_),
    .B2(_03082_),
    .X(_03083_));
 sky130_fd_sc_hd__a21o_1 _08069_ (.A1(\brancher.imm12_i_s[8] ),
    .A2(net764),
    .B1(net759),
    .X(_03084_));
 sky130_fd_sc_hd__o21a_1 _08070_ (.A1(net760),
    .A2(_03083_),
    .B1(_03084_),
    .X(_03085_));
 sky130_fd_sc_hd__inv_2 _08071_ (.A(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__and2_1 _08072_ (.A(_03081_),
    .B(_03085_),
    .X(_03087_));
 sky130_fd_sc_hd__nor2_1 _08073_ (.A(_03081_),
    .B(_03085_),
    .Y(_03088_));
 sky130_fd_sc_hd__nor2_1 _08074_ (.A(_03080_),
    .B(_03085_),
    .Y(_03089_));
 sky130_fd_sc_hd__inv_2 _08075_ (.A(_03089_),
    .Y(_03090_));
 sky130_fd_sc_hd__nor2_2 _08076_ (.A(_03087_),
    .B(_03088_),
    .Y(_03091_));
 sky130_fd_sc_hd__inv_2 _08077_ (.A(_03091_),
    .Y(_03092_));
 sky130_fd_sc_hd__or3_1 _08078_ (.A(_03059_),
    .B(_03075_),
    .C(_03091_),
    .X(_03093_));
 sky130_fd_sc_hd__or2_1 _08079_ (.A(_03028_),
    .B(_03093_),
    .X(_03094_));
 sky130_fd_sc_hd__inv_2 _08080_ (.A(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__a211o_1 _08081_ (.A1(_02736_),
    .A2(_02740_),
    .B1(_02967_),
    .C1(_03094_),
    .X(_03096_));
 sky130_fd_sc_hd__a32o_1 _08082_ (.A1(_02941_),
    .A2(_02943_),
    .A3(_02946_),
    .B1(_02955_),
    .B2(_02960_),
    .X(_03097_));
 sky130_fd_sc_hd__or4b_1 _08083_ (.A(_02921_),
    .B(_02935_),
    .C(_02963_),
    .D_N(_03097_),
    .X(_03098_));
 sky130_fd_sc_hd__or3_1 _08084_ (.A(_02914_),
    .B(_02918_),
    .C(_02934_),
    .X(_03099_));
 sky130_fd_sc_hd__a31oi_1 _08085_ (.A1(_02933_),
    .A2(_03098_),
    .A3(_03099_),
    .B1(_02907_),
    .Y(_03100_));
 sky130_fd_sc_hd__a22o_1 _08086_ (.A1(_02884_),
    .A2(_02889_),
    .B1(_02897_),
    .B2(_02902_),
    .X(_03101_));
 sky130_fd_sc_hd__nor3b_1 _08087_ (.A(_02879_),
    .B(_02903_),
    .C_N(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__a21oi_1 _08088_ (.A1(_02860_),
    .A2(_02876_),
    .B1(_02877_),
    .Y(_03103_));
 sky130_fd_sc_hd__o31a_1 _08089_ (.A1(_03100_),
    .A2(_03102_),
    .A3(_03103_),
    .B1(_02848_),
    .X(_03104_));
 sky130_fd_sc_hd__a32o_1 _08090_ (.A1(_02836_),
    .A2(_02838_),
    .A3(_02841_),
    .B1(_02825_),
    .B2(_02820_),
    .X(_03105_));
 sky130_fd_sc_hd__or4b_1 _08091_ (.A(_02798_),
    .B(_02813_),
    .C(_02828_),
    .D_N(_03105_),
    .X(_03106_));
 sky130_fd_sc_hd__o211ai_1 _08092_ (.A1(_02795_),
    .A2(_02811_),
    .B1(_02812_),
    .C1(_03106_),
    .Y(_03107_));
 sky130_fd_sc_hd__a21o_1 _08093_ (.A1(_02766_),
    .A2(_02782_),
    .B1(_02780_),
    .X(_03108_));
 sky130_fd_sc_hd__and3b_1 _08094_ (.A_N(_02600_),
    .B(_02746_),
    .C(_02750_),
    .X(_03109_));
 sky130_fd_sc_hd__a211o_1 _08095_ (.A1(_02753_),
    .A2(_03108_),
    .B1(_03109_),
    .C1(_02598_),
    .X(_03110_));
 sky130_fd_sc_hd__a31o_1 _08096_ (.A1(net183),
    .A2(_02784_),
    .A3(_03107_),
    .B1(_03110_),
    .X(_03111_));
 sky130_fd_sc_hd__o21a_1 _08097_ (.A1(_03018_),
    .A2(_03023_),
    .B1(_03011_),
    .X(_03112_));
 sky130_fd_sc_hd__or3b_1 _08098_ (.A(_03010_),
    .B(_03112_),
    .C_N(_02998_),
    .X(_03113_));
 sky130_fd_sc_hd__o21a_1 _08099_ (.A1(_02979_),
    .A2(_02996_),
    .B1(_02995_),
    .X(_03114_));
 sky130_fd_sc_hd__o2bb2a_1 _08100_ (.A1_N(_03065_),
    .A2_N(_03070_),
    .B1(_03081_),
    .B2(_03086_),
    .X(_03115_));
 sky130_fd_sc_hd__o41a_1 _08101_ (.A1(_03035_),
    .A2(_03038_),
    .A3(_03039_),
    .A4(_03055_),
    .B1(_03056_),
    .X(_03116_));
 sky130_fd_sc_hd__o31a_1 _08102_ (.A1(_03059_),
    .A2(_03071_),
    .A3(_03115_),
    .B1(_03116_),
    .X(_03117_));
 sky130_fd_sc_hd__o211ai_2 _08103_ (.A1(_03028_),
    .A2(_03117_),
    .B1(_03114_),
    .C1(_03113_),
    .Y(_03118_));
 sky130_fd_sc_hd__a311oi_2 _08104_ (.A1(_02848_),
    .A2(_02966_),
    .A3(_03118_),
    .B1(_03111_),
    .C1(_03104_),
    .Y(_03119_));
 sky130_fd_sc_hd__nand2_1 _08105_ (.A(_03096_),
    .B(_03119_),
    .Y(_03120_));
 sky130_fd_sc_hd__a21oi_2 _08106_ (.A1(_02676_),
    .A2(_02677_),
    .B1(net236),
    .Y(_03121_));
 sky130_fd_sc_hd__a21o_1 _08107_ (.A1(_02676_),
    .A2(_02677_),
    .B1(net236),
    .X(_03122_));
 sky130_fd_sc_hd__nand3_2 _08108_ (.A(_02676_),
    .B(_02677_),
    .C(net236),
    .Y(_03123_));
 sky130_fd_sc_hd__and3_1 _08109_ (.A(net229),
    .B(net714),
    .C(_02697_),
    .X(_03124_));
 sky130_fd_sc_hd__a21o_1 _08110_ (.A1(_03122_),
    .A2(_03123_),
    .B1(_03124_),
    .X(_03125_));
 sky130_fd_sc_hd__or3_1 _08111_ (.A(_02698_),
    .B(_02714_),
    .C(_02733_),
    .X(_03126_));
 sky130_fd_sc_hd__or3_1 _08112_ (.A(_02670_),
    .B(_03125_),
    .C(_03126_),
    .X(_03127_));
 sky130_fd_sc_hd__o311a_1 _08113_ (.A1(_02967_),
    .A2(_03094_),
    .A3(_03127_),
    .B1(_01218_),
    .C1(net846),
    .X(_03128_));
 sky130_fd_sc_hd__nor2_2 _08114_ (.A(\alu.b_type ),
    .B(net951),
    .Y(_03129_));
 sky130_fd_sc_hd__o21ai_2 _08115_ (.A1(\alu.r_type ),
    .A2(\alu.op_consShf ),
    .B1(\brancher.imm13_b[10] ),
    .Y(_03130_));
 sky130_fd_sc_hd__o21ai_2 _08116_ (.A1(net951),
    .A2(_03130_),
    .B1(_01209_),
    .Y(_03131_));
 sky130_fd_sc_hd__a21o_1 _08117_ (.A1(net847),
    .A2(_03129_),
    .B1(net688),
    .X(_03132_));
 sky130_fd_sc_hd__or4b_1 _08118_ (.A(net948),
    .B(_03132_),
    .C(_02598_),
    .D_N(_03128_),
    .X(_03133_));
 sky130_fd_sc_hd__o21ba_1 _08119_ (.A1(_02602_),
    .A2(_03120_),
    .B1_N(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__nand3_1 _08120_ (.A(net847),
    .B(_03129_),
    .C(_03130_),
    .Y(_03135_));
 sky130_fd_sc_hd__and4_1 _08121_ (.A(net847),
    .B(_03128_),
    .C(_03129_),
    .D(_03130_),
    .X(_03136_));
 sky130_fd_sc_hd__nand2_2 _08122_ (.A(net943),
    .B(_03129_),
    .Y(_03137_));
 sky130_fd_sc_hd__nor2_1 _08123_ (.A(_01227_),
    .B(_03137_),
    .Y(_03138_));
 sky130_fd_sc_hd__or2_2 _08124_ (.A(_01227_),
    .B(_03137_),
    .X(_03139_));
 sky130_fd_sc_hd__and3_1 _08125_ (.A(net231),
    .B(net716),
    .C(_02773_),
    .X(_03140_));
 sky130_fd_sc_hd__a21oi_1 _08126_ (.A1(net189),
    .A2(_02760_),
    .B1(_03140_),
    .Y(_03141_));
 sky130_fd_sc_hd__o21a_1 _08127_ (.A1(net234),
    .A2(net719),
    .B1(_02746_),
    .X(_03142_));
 sky130_fd_sc_hd__a21oi_1 _08128_ (.A1(net199),
    .A2(net190),
    .B1(_03142_),
    .Y(_03143_));
 sky130_fd_sc_hd__mux2_2 _08129_ (.A0(_03141_),
    .A1(_03143_),
    .S(net247),
    .X(_03144_));
 sky130_fd_sc_hd__a21o_1 _08130_ (.A1(net231),
    .A2(net716),
    .B1(_02790_),
    .X(_03145_));
 sky130_fd_sc_hd__or3b_1 _08131_ (.A(net234),
    .B(net719),
    .C_N(_02804_),
    .X(_03146_));
 sky130_fd_sc_hd__a21o_1 _08132_ (.A1(net231),
    .A2(net716),
    .B1(_02837_),
    .X(_03147_));
 sky130_fd_sc_hd__or3_1 _08133_ (.A(net234),
    .B(net719),
    .C(_02821_),
    .X(_03148_));
 sky130_fd_sc_hd__and3_1 _08134_ (.A(net242),
    .B(_03147_),
    .C(_03148_),
    .X(_03149_));
 sky130_fd_sc_hd__a31o_1 _08135_ (.A1(net247),
    .A2(_03145_),
    .A3(_03146_),
    .B1(_03149_),
    .X(_03150_));
 sky130_fd_sc_hd__mux2_2 _08136_ (.A0(_03144_),
    .A1(_03150_),
    .S(net224),
    .X(_03151_));
 sky130_fd_sc_hd__a21o_1 _08137_ (.A1(net231),
    .A2(net716),
    .B1(_02854_),
    .X(_03152_));
 sky130_fd_sc_hd__or3_1 _08138_ (.A(net234),
    .B(net719),
    .C(_02869_),
    .X(_03153_));
 sky130_fd_sc_hd__and3_1 _08139_ (.A(net248),
    .B(_03152_),
    .C(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__or3_1 _08140_ (.A(net234),
    .B(net719),
    .C(_02898_),
    .X(_03155_));
 sky130_fd_sc_hd__a21o_1 _08141_ (.A1(net231),
    .A2(net716),
    .B1(_02885_),
    .X(_03156_));
 sky130_fd_sc_hd__and3_1 _08142_ (.A(net241),
    .B(_03155_),
    .C(_03156_),
    .X(_03157_));
 sky130_fd_sc_hd__or2_1 _08143_ (.A(_03154_),
    .B(_03157_),
    .X(_03158_));
 sky130_fd_sc_hd__a21o_1 _08144_ (.A1(net231),
    .A2(net716),
    .B1(_02914_),
    .X(_03159_));
 sky130_fd_sc_hd__a21boi_1 _08145_ (.A1(net190),
    .A2(_02926_),
    .B1_N(_03159_),
    .Y(_03160_));
 sky130_fd_sc_hd__or3_1 _08146_ (.A(net233),
    .B(net718),
    .C(_02956_),
    .X(_03161_));
 sky130_fd_sc_hd__o21a_1 _08147_ (.A1(net190),
    .A2(_02942_),
    .B1(_03161_),
    .X(_03162_));
 sky130_fd_sc_hd__mux2_1 _08148_ (.A0(_03160_),
    .A1(_03162_),
    .S(net239),
    .X(_03163_));
 sky130_fd_sc_hd__mux2_1 _08149_ (.A0(_03158_),
    .A1(_03163_),
    .S(net220),
    .X(_03164_));
 sky130_fd_sc_hd__mux2_1 _08150_ (.A0(_03151_),
    .A1(_03164_),
    .S(net207),
    .X(_03165_));
 sky130_fd_sc_hd__and3_1 _08151_ (.A(net195),
    .B(net573),
    .C(_03165_),
    .X(_03166_));
 sky130_fd_sc_hd__nor3_2 _08152_ (.A(net233),
    .B(net718),
    .C(_02697_),
    .Y(_03167_));
 sky130_fd_sc_hd__inv_2 _08153_ (.A(_03167_),
    .Y(_03168_));
 sky130_fd_sc_hd__nor3_2 _08154_ (.A(net813),
    .B(_03135_),
    .C(_03137_),
    .Y(_03169_));
 sky130_fd_sc_hd__or3_4 _08155_ (.A(_01217_),
    .B(_03135_),
    .C(_03137_),
    .X(_03170_));
 sky130_fd_sc_hd__or3_2 _08156_ (.A(net846),
    .B(\brancher.funct3[2] ),
    .C(_03135_),
    .X(_03171_));
 sky130_fd_sc_hd__inv_2 _08157_ (.A(_03171_),
    .Y(_03172_));
 sky130_fd_sc_hd__nand2_4 _08158_ (.A(net192),
    .B(net209),
    .Y(_03173_));
 sky130_fd_sc_hd__nor2_4 _08159_ (.A(net227),
    .B(_03173_),
    .Y(_03174_));
 sky130_fd_sc_hd__and2_1 _08160_ (.A(_03172_),
    .B(_03174_),
    .X(_03175_));
 sky130_fd_sc_hd__nor2_4 _08161_ (.A(net194),
    .B(_03171_),
    .Y(_03176_));
 sky130_fd_sc_hd__nand2_1 _08162_ (.A(net192),
    .B(_03172_),
    .Y(_03177_));
 sky130_fd_sc_hd__nor2_1 _08163_ (.A(net210),
    .B(_03171_),
    .Y(_03178_));
 sky130_fd_sc_hd__nand2_1 _08164_ (.A(net208),
    .B(_03172_),
    .Y(_03179_));
 sky130_fd_sc_hd__nor2_2 _08165_ (.A(net194),
    .B(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__nand2_1 _08166_ (.A(net187),
    .B(_02697_),
    .Y(_03181_));
 sky130_fd_sc_hd__nor2_1 _08167_ (.A(_03132_),
    .B(_03137_),
    .Y(_03182_));
 sky130_fd_sc_hd__or2_2 _08168_ (.A(_03132_),
    .B(_03137_),
    .X(_03183_));
 sky130_fd_sc_hd__nor2_1 _08169_ (.A(net813),
    .B(_03183_),
    .Y(_03184_));
 sky130_fd_sc_hd__nand2_4 _08170_ (.A(net845),
    .B(net430),
    .Y(_03185_));
 sky130_fd_sc_hd__nand2_1 _08171_ (.A(_01218_),
    .B(wRamByteEn),
    .Y(_03186_));
 sky130_fd_sc_hd__nand2_2 _08172_ (.A(_03129_),
    .B(_03186_),
    .Y(_03187_));
 sky130_fd_sc_hd__o221a_1 _08173_ (.A1(_03168_),
    .A2(net265),
    .B1(_03187_),
    .B2(net430),
    .C1(_03181_),
    .X(_03188_));
 sky130_fd_sc_hd__a221o_1 _08174_ (.A1(_03167_),
    .A2(net570),
    .B1(_03175_),
    .B2(_02700_),
    .C1(_03188_),
    .X(_03189_));
 sky130_fd_sc_hd__and3_1 _08175_ (.A(net230),
    .B(net715),
    .C(net205),
    .X(_03190_));
 sky130_fd_sc_hd__a21oi_1 _08176_ (.A1(net189),
    .A2(_02972_),
    .B1(_03190_),
    .Y(_03191_));
 sky130_fd_sc_hd__mux2_1 _08177_ (.A0(_03004_),
    .A1(_03018_),
    .S(net188),
    .X(_03192_));
 sky130_fd_sc_hd__mux2_1 _08178_ (.A0(_03191_),
    .A1(_03192_),
    .S(net239),
    .X(_03193_));
 sky130_fd_sc_hd__or3_1 _08179_ (.A(net233),
    .B(net718),
    .C(_03049_),
    .X(_03194_));
 sky130_fd_sc_hd__a21o_1 _08180_ (.A1(net230),
    .A2(net715),
    .B1(_03035_),
    .X(_03195_));
 sky130_fd_sc_hd__or3_1 _08181_ (.A(net233),
    .B(net718),
    .C(_03066_),
    .X(_03196_));
 sky130_fd_sc_hd__a21o_1 _08182_ (.A1(net229),
    .A2(net714),
    .B1(_03081_),
    .X(_03197_));
 sky130_fd_sc_hd__a21o_1 _08183_ (.A1(_03196_),
    .A2(_03197_),
    .B1(net245),
    .X(_03198_));
 sky130_fd_sc_hd__a21o_1 _08184_ (.A1(_03194_),
    .A2(_03195_),
    .B1(net240),
    .X(_03199_));
 sky130_fd_sc_hd__and3_1 _08185_ (.A(net217),
    .B(_03198_),
    .C(_03199_),
    .X(_03200_));
 sky130_fd_sc_hd__a211o_1 _08186_ (.A1(net226),
    .A2(_03193_),
    .B1(_03200_),
    .C1(net206),
    .X(_03201_));
 sky130_fd_sc_hd__nor2_4 _08187_ (.A(net196),
    .B(_03139_),
    .Y(_03202_));
 sky130_fd_sc_hd__nand2_1 _08188_ (.A(_02678_),
    .B(net190),
    .Y(_03203_));
 sky130_fd_sc_hd__o21a_1 _08189_ (.A1(net233),
    .A2(net718),
    .B1(_02711_),
    .X(_03204_));
 sky130_fd_sc_hd__and3_1 _08190_ (.A(net229),
    .B(net714),
    .C(_02727_),
    .X(_03205_));
 sky130_fd_sc_hd__nor2_1 _08191_ (.A(_03204_),
    .B(_03205_),
    .Y(_03206_));
 sky130_fd_sc_hd__mux2_1 _08192_ (.A0(_02610_),
    .A1(_02628_),
    .S(net190),
    .X(_03207_));
 sky130_fd_sc_hd__and3_1 _08193_ (.A(_02659_),
    .B(net229),
    .C(net714),
    .X(_03208_));
 sky130_fd_sc_hd__a21oi_1 _08194_ (.A1(_02650_),
    .A2(net187),
    .B1(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__mux2_1 _08195_ (.A0(_03207_),
    .A1(_03209_),
    .S(net237),
    .X(_03210_));
 sky130_fd_sc_hd__a21o_1 _08196_ (.A1(_03181_),
    .A2(_03203_),
    .B1(net246),
    .X(_03211_));
 sky130_fd_sc_hd__o21a_1 _08197_ (.A1(net237),
    .A2(_03206_),
    .B1(net216),
    .X(_03212_));
 sky130_fd_sc_hd__a221o_1 _08198_ (.A1(net226),
    .A2(_03210_),
    .B1(_03211_),
    .B2(_03212_),
    .C1(net210),
    .X(_03213_));
 sky130_fd_sc_hd__a31o_1 _08199_ (.A1(_03201_),
    .A2(_03202_),
    .A3(_03213_),
    .B1(_03189_),
    .X(_03214_));
 sky130_fd_sc_hd__a211o_1 _08200_ (.A1(_03120_),
    .A2(_03136_),
    .B1(_03166_),
    .C1(_03214_),
    .X(_03215_));
 sky130_fd_sc_hd__nor2_1 _08201_ (.A(_03134_),
    .B(_03215_),
    .Y(_03216_));
 sky130_fd_sc_hd__nor2_4 _08202_ (.A(net952),
    .B(net957),
    .Y(_03217_));
 sky130_fd_sc_hd__or2_4 _08203_ (.A(net952),
    .B(net956),
    .X(_03218_));
 sky130_fd_sc_hd__and3b_1 _08204_ (.A_N(\dec.op_lui ),
    .B(_02575_),
    .C(_03218_),
    .X(_03219_));
 sky130_fd_sc_hd__a2bb2o_1 _08205_ (.A1_N(_02575_),
    .A2_N(_03216_),
    .B1(net566),
    .B2(net1439),
    .X(_00002_));
 sky130_fd_sc_hd__and2_2 _08206_ (.A(_03131_),
    .B(net573),
    .X(_03220_));
 sky130_fd_sc_hd__nand2_2 _08207_ (.A(net688),
    .B(net573),
    .Y(_03221_));
 sky130_fd_sc_hd__or3_1 _08208_ (.A(net234),
    .B(net719),
    .C(_02837_),
    .X(_03222_));
 sky130_fd_sc_hd__a21o_1 _08209_ (.A1(net231),
    .A2(net716),
    .B1(_02869_),
    .X(_03223_));
 sky130_fd_sc_hd__or3_1 _08210_ (.A(net234),
    .B(net719),
    .C(_02854_),
    .X(_03224_));
 sky130_fd_sc_hd__a21o_1 _08211_ (.A1(net231),
    .A2(net716),
    .B1(_02898_),
    .X(_03225_));
 sky130_fd_sc_hd__a21o_1 _08212_ (.A1(_03224_),
    .A2(_03225_),
    .B1(net249),
    .X(_03226_));
 sky130_fd_sc_hd__a21o_1 _08213_ (.A1(_03222_),
    .A2(_03223_),
    .B1(net242),
    .X(_03227_));
 sky130_fd_sc_hd__and3_1 _08214_ (.A(net228),
    .B(_03226_),
    .C(_03227_),
    .X(_03228_));
 sky130_fd_sc_hd__or3_1 _08215_ (.A(net234),
    .B(net719),
    .C(_02885_),
    .X(_03229_));
 sky130_fd_sc_hd__o21ai_1 _08216_ (.A1(net234),
    .A2(net719),
    .B1(_02926_),
    .Y(_03230_));
 sky130_fd_sc_hd__and2_1 _08217_ (.A(_03229_),
    .B(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__or3_1 _08218_ (.A(net234),
    .B(net719),
    .C(_02914_),
    .X(_03232_));
 sky130_fd_sc_hd__a21o_1 _08219_ (.A1(net231),
    .A2(net716),
    .B1(_02956_),
    .X(_03233_));
 sky130_fd_sc_hd__and2_1 _08220_ (.A(_03232_),
    .B(_03233_),
    .X(_03234_));
 sky130_fd_sc_hd__mux2_1 _08221_ (.A0(_03231_),
    .A1(_03234_),
    .S(net241),
    .X(_03235_));
 sky130_fd_sc_hd__a21o_1 _08222_ (.A1(net225),
    .A2(_03235_),
    .B1(_03228_),
    .X(_03236_));
 sky130_fd_sc_hd__and3_1 _08223_ (.A(net232),
    .B(net717),
    .C(_02761_),
    .X(_03237_));
 sky130_fd_sc_hd__a21oi_1 _08224_ (.A1(net232),
    .A2(net717),
    .B1(_02804_),
    .Y(_03238_));
 sky130_fd_sc_hd__or3_1 _08225_ (.A(net235),
    .B(net720),
    .C(_02790_),
    .X(_03239_));
 sky130_fd_sc_hd__a21o_1 _08226_ (.A1(net232),
    .A2(net717),
    .B1(_02821_),
    .X(_03240_));
 sky130_fd_sc_hd__a21o_1 _08227_ (.A1(_03239_),
    .A2(_03240_),
    .B1(net248),
    .X(_03241_));
 sky130_fd_sc_hd__or3_1 _08228_ (.A(net243),
    .B(_03237_),
    .C(_03238_),
    .X(_03242_));
 sky130_fd_sc_hd__a21o_1 _08229_ (.A1(_03241_),
    .A2(_03242_),
    .B1(net228),
    .X(_03243_));
 sky130_fd_sc_hd__or3_1 _08230_ (.A(net235),
    .B(net720),
    .C(_02746_),
    .X(_03244_));
 sky130_fd_sc_hd__a21o_1 _08231_ (.A1(net231),
    .A2(net716),
    .B1(_02773_),
    .X(_03245_));
 sky130_fd_sc_hd__a21oi_1 _08232_ (.A1(_03244_),
    .A2(_03245_),
    .B1(net247),
    .Y(_03246_));
 sky130_fd_sc_hd__a21o_1 _08233_ (.A1(_03244_),
    .A2(_03245_),
    .B1(net247),
    .X(_03247_));
 sky130_fd_sc_hd__nor2_1 _08234_ (.A(net198),
    .B(net243),
    .Y(_03248_));
 sky130_fd_sc_hd__or3_1 _08235_ (.A(net222),
    .B(_03246_),
    .C(_03248_),
    .X(_03249_));
 sky130_fd_sc_hd__and2_1 _08236_ (.A(_03243_),
    .B(_03249_),
    .X(_03250_));
 sky130_fd_sc_hd__mux2_1 _08237_ (.A0(_03236_),
    .A1(_03250_),
    .S(net211),
    .X(_03251_));
 sky130_fd_sc_hd__or3_1 _08238_ (.A(net199),
    .B(net243),
    .C(net190),
    .X(_03252_));
 sky130_fd_sc_hd__or3b_1 _08239_ (.A(net222),
    .B(_03246_),
    .C_N(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__a21o_1 _08240_ (.A1(_03243_),
    .A2(_03253_),
    .B1(net208),
    .X(_03254_));
 sky130_fd_sc_hd__nor2_2 _08241_ (.A(_03131_),
    .B(_03139_),
    .Y(_03255_));
 sky130_fd_sc_hd__or2_1 _08242_ (.A(net688),
    .B(_03139_),
    .X(_03256_));
 sky130_fd_sc_hd__o211a_1 _08243_ (.A1(net211),
    .A2(_03236_),
    .B1(_03254_),
    .C1(_03255_),
    .X(_03257_));
 sky130_fd_sc_hd__a21o_1 _08244_ (.A1(_03220_),
    .A2(_03251_),
    .B1(_03257_),
    .X(_03258_));
 sky130_fd_sc_hd__and2_1 _08245_ (.A(net688),
    .B(_03187_),
    .X(_03259_));
 sky130_fd_sc_hd__nand2_1 _08246_ (.A(net688),
    .B(_03187_),
    .Y(_03260_));
 sky130_fd_sc_hd__nand2_1 _08247_ (.A(_03125_),
    .B(net428),
    .Y(_03261_));
 sky130_fd_sc_hd__a31oi_1 _08248_ (.A1(_03122_),
    .A2(_03123_),
    .A3(_03124_),
    .B1(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__nand2_1 _08249_ (.A(net813),
    .B(_03121_),
    .Y(_03263_));
 sky130_fd_sc_hd__a32o_1 _08250_ (.A1(_03123_),
    .A2(net430),
    .A3(_03263_),
    .B1(net570),
    .B2(_03121_),
    .X(_03264_));
 sky130_fd_sc_hd__or3b_1 _08251_ (.A(_03121_),
    .B(_03168_),
    .C_N(_03123_),
    .X(_03265_));
 sky130_fd_sc_hd__and2b_1 _08252_ (.A_N(net688),
    .B(_03187_),
    .X(_03266_));
 sky130_fd_sc_hd__nand2b_4 _08253_ (.A_N(net688),
    .B(_03187_),
    .Y(_03267_));
 sky130_fd_sc_hd__a21o_1 _08254_ (.A1(_03122_),
    .A2(_03123_),
    .B1(_03167_),
    .X(_03268_));
 sky130_fd_sc_hd__and3_1 _08255_ (.A(_03265_),
    .B(net423),
    .C(_03268_),
    .X(_03269_));
 sky130_fd_sc_hd__a21oi_1 _08256_ (.A1(_02678_),
    .A2(net187),
    .B1(_03124_),
    .Y(_03270_));
 sky130_fd_sc_hd__and2_1 _08257_ (.A(net236),
    .B(_03270_),
    .X(_03271_));
 sky130_fd_sc_hd__a31o_1 _08258_ (.A1(net216),
    .A2(_03180_),
    .A3(_03271_),
    .B1(_03264_),
    .X(_03272_));
 sky130_fd_sc_hd__or3_1 _08259_ (.A(_03262_),
    .B(_03269_),
    .C(_03272_),
    .X(_03273_));
 sky130_fd_sc_hd__and3_1 _08260_ (.A(net229),
    .B(net714),
    .C(_03080_),
    .X(_03274_));
 sky130_fd_sc_hd__a21oi_1 _08261_ (.A1(_02627_),
    .A2(net188),
    .B1(_03274_),
    .Y(_03275_));
 sky130_fd_sc_hd__a211o_1 _08262_ (.A1(_02627_),
    .A2(net188),
    .B1(_03274_),
    .C1(net240),
    .X(_03276_));
 sky130_fd_sc_hd__and3_1 _08263_ (.A(_02609_),
    .B(net229),
    .C(net714),
    .X(_03277_));
 sky130_fd_sc_hd__a21o_1 _08264_ (.A1(_02659_),
    .A2(net187),
    .B1(_03277_),
    .X(_03278_));
 sky130_fd_sc_hd__o21ai_1 _08265_ (.A1(net246),
    .A2(_03278_),
    .B1(_03276_),
    .Y(_03279_));
 sky130_fd_sc_hd__and3_1 _08266_ (.A(net229),
    .B(net714),
    .C(_02711_),
    .X(_03280_));
 sky130_fd_sc_hd__a211o_1 _08267_ (.A1(_02678_),
    .A2(net187),
    .B1(_03280_),
    .C1(net246),
    .X(_03281_));
 sky130_fd_sc_hd__and3_1 _08268_ (.A(_02650_),
    .B(net229),
    .C(net714),
    .X(_03282_));
 sky130_fd_sc_hd__a21o_1 _08269_ (.A1(net187),
    .A2(_02727_),
    .B1(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__o21a_1 _08270_ (.A1(net237),
    .A2(_03283_),
    .B1(net217),
    .X(_03284_));
 sky130_fd_sc_hd__a2bb2o_1 _08271_ (.A1_N(net217),
    .A2_N(_03279_),
    .B1(_03281_),
    .B2(_03284_),
    .X(_03285_));
 sky130_fd_sc_hd__or3_2 _08272_ (.A(net233),
    .B(net718),
    .C(_02942_),
    .X(_03286_));
 sky130_fd_sc_hd__o21ai_1 _08273_ (.A1(net233),
    .A2(net718),
    .B1(net205),
    .Y(_03287_));
 sky130_fd_sc_hd__or3_1 _08274_ (.A(net235),
    .B(net720),
    .C(_02973_),
    .X(_03288_));
 sky130_fd_sc_hd__a21o_1 _08275_ (.A1(net229),
    .A2(net714),
    .B1(_03004_),
    .X(_03289_));
 sky130_fd_sc_hd__and3_1 _08276_ (.A(net240),
    .B(_03288_),
    .C(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__a31o_1 _08277_ (.A1(net246),
    .A2(_03286_),
    .A3(_03287_),
    .B1(_03290_),
    .X(_03291_));
 sky130_fd_sc_hd__or3_1 _08278_ (.A(net233),
    .B(net718),
    .C(_03018_),
    .X(_03292_));
 sky130_fd_sc_hd__a21o_1 _08279_ (.A1(net230),
    .A2(net715),
    .B1(_03049_),
    .X(_03293_));
 sky130_fd_sc_hd__and2_1 _08280_ (.A(_03292_),
    .B(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__or3_1 _08281_ (.A(net233),
    .B(net718),
    .C(_03035_),
    .X(_03295_));
 sky130_fd_sc_hd__a21o_1 _08282_ (.A1(net230),
    .A2(net715),
    .B1(_03066_),
    .X(_03296_));
 sky130_fd_sc_hd__and3_1 _08283_ (.A(net240),
    .B(_03295_),
    .C(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__a21o_1 _08284_ (.A1(net245),
    .A2(_03294_),
    .B1(_03297_),
    .X(_03298_));
 sky130_fd_sc_hd__mux2_1 _08285_ (.A0(_03291_),
    .A1(_03298_),
    .S(net218),
    .X(_03299_));
 sky130_fd_sc_hd__nand2_1 _08286_ (.A(net206),
    .B(_03285_),
    .Y(_03300_));
 sky130_fd_sc_hd__o211a_1 _08287_ (.A1(net207),
    .A2(_03299_),
    .B1(_03300_),
    .C1(_03202_),
    .X(_03301_));
 sky130_fd_sc_hd__a211o_1 _08288_ (.A1(net194),
    .A2(_03258_),
    .B1(_03273_),
    .C1(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__a22o_1 _08289_ (.A1(net1347),
    .A2(net566),
    .B1(_03302_),
    .B2(net740),
    .X(_00013_));
 sky130_fd_sc_hd__a21o_1 _08290_ (.A1(_03152_),
    .A2(_03153_),
    .B1(net248),
    .X(_03303_));
 sky130_fd_sc_hd__a21o_1 _08291_ (.A1(_03147_),
    .A2(_03148_),
    .B1(net242),
    .X(_03304_));
 sky130_fd_sc_hd__and3_1 _08292_ (.A(net249),
    .B(_03155_),
    .C(_03156_),
    .X(_03305_));
 sky130_fd_sc_hd__a211o_1 _08293_ (.A1(net241),
    .A2(_03160_),
    .B1(_03305_),
    .C1(net227),
    .X(_03306_));
 sky130_fd_sc_hd__a21o_1 _08294_ (.A1(_03303_),
    .A2(_03304_),
    .B1(net224),
    .X(_03307_));
 sky130_fd_sc_hd__a21oi_1 _08295_ (.A1(_03306_),
    .A2(_03307_),
    .B1(net213),
    .Y(_03308_));
 sky130_fd_sc_hd__a21o_1 _08296_ (.A1(net243),
    .A2(_03143_),
    .B1(net222),
    .X(_03309_));
 sky130_fd_sc_hd__a21o_1 _08297_ (.A1(_03145_),
    .A2(_03146_),
    .B1(net247),
    .X(_03310_));
 sky130_fd_sc_hd__o21a_1 _08298_ (.A1(net243),
    .A2(_03141_),
    .B1(_03310_),
    .X(_03311_));
 sky130_fd_sc_hd__o21ai_2 _08299_ (.A1(net227),
    .A2(_03311_),
    .B1(_03309_),
    .Y(_03312_));
 sky130_fd_sc_hd__a211o_1 _08300_ (.A1(net212),
    .A2(_03312_),
    .B1(_03308_),
    .C1(_03256_),
    .X(_03313_));
 sky130_fd_sc_hd__o21ai_1 _08301_ (.A1(net227),
    .A2(_03311_),
    .B1(_03248_),
    .Y(_03314_));
 sky130_fd_sc_hd__a31o_1 _08302_ (.A1(net212),
    .A2(_03312_),
    .A3(_03314_),
    .B1(_03308_),
    .X(_03315_));
 sky130_fd_sc_hd__a311o_1 _08303_ (.A1(net212),
    .A2(_03312_),
    .A3(_03314_),
    .B1(_03221_),
    .C1(_03308_),
    .X(_03316_));
 sky130_fd_sc_hd__a21oi_1 _08304_ (.A1(_03313_),
    .A2(_03316_),
    .B1(net191),
    .Y(_03317_));
 sky130_fd_sc_hd__a21o_1 _08305_ (.A1(_03123_),
    .A2(_03167_),
    .B1(_03121_),
    .X(_03318_));
 sky130_fd_sc_hd__nand2_1 _08306_ (.A(_02714_),
    .B(_03318_),
    .Y(_03319_));
 sky130_fd_sc_hd__or2_1 _08307_ (.A(_02714_),
    .B(_03318_),
    .X(_03320_));
 sky130_fd_sc_hd__or2_1 _08308_ (.A(_02678_),
    .B(net246),
    .X(_03321_));
 sky130_fd_sc_hd__a21o_1 _08309_ (.A1(_03125_),
    .A2(_03321_),
    .B1(_02714_),
    .X(_03322_));
 sky130_fd_sc_hd__a31o_1 _08310_ (.A1(_02714_),
    .A2(_03125_),
    .A3(_03321_),
    .B1(net426),
    .X(_03323_));
 sky130_fd_sc_hd__and2b_1 _08311_ (.A_N(_03323_),
    .B(_03322_),
    .X(_03324_));
 sky130_fd_sc_hd__a21oi_1 _08312_ (.A1(_02678_),
    .A2(net190),
    .B1(_03204_),
    .Y(_03325_));
 sky130_fd_sc_hd__mux2_1 _08313_ (.A0(_02698_),
    .A1(_03325_),
    .S(net237),
    .X(_03326_));
 sky130_fd_sc_hd__nor2_1 _08314_ (.A(net216),
    .B(_02711_),
    .Y(_03327_));
 sky130_fd_sc_hd__nor2_1 _08315_ (.A(_02711_),
    .B(_03185_),
    .Y(_03328_));
 sky130_fd_sc_hd__a221o_1 _08316_ (.A1(_02714_),
    .A2(net430),
    .B1(_03327_),
    .B2(net570),
    .C1(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__a211o_1 _08317_ (.A1(_03175_),
    .A2(_03326_),
    .B1(_03329_),
    .C1(_03324_),
    .X(_03330_));
 sky130_fd_sc_hd__a31o_1 _08318_ (.A1(net423),
    .A2(_03319_),
    .A3(_03320_),
    .B1(_03330_),
    .X(_03331_));
 sky130_fd_sc_hd__and3_1 _08319_ (.A(net246),
    .B(_03196_),
    .C(_03197_),
    .X(_03332_));
 sky130_fd_sc_hd__a21o_1 _08320_ (.A1(net236),
    .A2(_03207_),
    .B1(_03332_),
    .X(_03333_));
 sky130_fd_sc_hd__mux2_1 _08321_ (.A0(_03206_),
    .A1(_03209_),
    .S(net246),
    .X(_03334_));
 sky130_fd_sc_hd__mux2_1 _08322_ (.A0(_03333_),
    .A1(_03334_),
    .S(net217),
    .X(_03335_));
 sky130_fd_sc_hd__mux2_1 _08323_ (.A0(_03162_),
    .A1(_03191_),
    .S(net239),
    .X(_03336_));
 sky130_fd_sc_hd__and3_1 _08324_ (.A(net240),
    .B(_03194_),
    .C(_03195_),
    .X(_03337_));
 sky130_fd_sc_hd__a21o_1 _08325_ (.A1(net245),
    .A2(_03192_),
    .B1(_03337_),
    .X(_03338_));
 sky130_fd_sc_hd__mux2_1 _08326_ (.A0(_03336_),
    .A1(_03338_),
    .S(net218),
    .X(_03339_));
 sky130_fd_sc_hd__mux2_1 _08327_ (.A0(_03335_),
    .A1(_03339_),
    .S(net210),
    .X(_03340_));
 sky130_fd_sc_hd__a211o_1 _08328_ (.A1(_03202_),
    .A2(_03340_),
    .B1(_03331_),
    .C1(_03317_),
    .X(_03341_));
 sky130_fd_sc_hd__a22o_1 _08329_ (.A1(net1323),
    .A2(net567),
    .B1(_03341_),
    .B2(net740),
    .X(_00024_));
 sky130_fd_sc_hd__a21o_1 _08330_ (.A1(_03222_),
    .A2(_03223_),
    .B1(net248),
    .X(_03342_));
 sky130_fd_sc_hd__a21o_1 _08331_ (.A1(_03239_),
    .A2(_03240_),
    .B1(net242),
    .X(_03343_));
 sky130_fd_sc_hd__and3_1 _08332_ (.A(net248),
    .B(_03224_),
    .C(_03225_),
    .X(_03344_));
 sky130_fd_sc_hd__a211o_1 _08333_ (.A1(net242),
    .A2(_03231_),
    .B1(_03344_),
    .C1(net227),
    .X(_03345_));
 sky130_fd_sc_hd__a21o_1 _08334_ (.A1(_03342_),
    .A2(_03343_),
    .B1(net224),
    .X(_03346_));
 sky130_fd_sc_hd__a21oi_2 _08335_ (.A1(_03345_),
    .A2(_03346_),
    .B1(net212),
    .Y(_03347_));
 sky130_fd_sc_hd__or3_1 _08336_ (.A(net247),
    .B(_03237_),
    .C(_03238_),
    .X(_03348_));
 sky130_fd_sc_hd__nand3_1 _08337_ (.A(_02682_),
    .B(_03244_),
    .C(_03245_),
    .Y(_03349_));
 sky130_fd_sc_hd__nand3_2 _08338_ (.A(net224),
    .B(_03348_),
    .C(_03349_),
    .Y(_03350_));
 sky130_fd_sc_hd__or2_1 _08339_ (.A(net198),
    .B(net223),
    .X(_03351_));
 sky130_fd_sc_hd__nand2_1 _08340_ (.A(net212),
    .B(_03351_),
    .Y(_03352_));
 sky130_fd_sc_hd__a31o_1 _08341_ (.A1(net212),
    .A2(_03350_),
    .A3(_03351_),
    .B1(_03347_),
    .X(_03353_));
 sky130_fd_sc_hd__and3b_1 _08342_ (.A_N(net199),
    .B(net243),
    .C(net189),
    .X(_03354_));
 sky130_fd_sc_hd__a21bo_1 _08343_ (.A1(net227),
    .A2(_03354_),
    .B1_N(_03350_),
    .X(_03355_));
 sky130_fd_sc_hd__o21ai_1 _08344_ (.A1(net209),
    .A2(_03355_),
    .B1(_03255_),
    .Y(_03356_));
 sky130_fd_sc_hd__nor2_1 _08345_ (.A(_03347_),
    .B(_03356_),
    .Y(_03357_));
 sky130_fd_sc_hd__o22ai_2 _08346_ (.A1(_03221_),
    .A2(_03353_),
    .B1(_03356_),
    .B2(_03347_),
    .Y(_03358_));
 sky130_fd_sc_hd__a21oi_1 _08347_ (.A1(_02713_),
    .A2(_03322_),
    .B1(_02733_),
    .Y(_03359_));
 sky130_fd_sc_hd__a31o_1 _08348_ (.A1(_02713_),
    .A2(_02733_),
    .A3(_03322_),
    .B1(net426),
    .X(_03360_));
 sky130_fd_sc_hd__nor2_1 _08349_ (.A(_03359_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__a21oi_1 _08350_ (.A1(net187),
    .A2(_02727_),
    .B1(_03280_),
    .Y(_03362_));
 sky130_fd_sc_hd__mux2_2 _08351_ (.A0(_03270_),
    .A1(_03362_),
    .S(net236),
    .X(_03363_));
 sky130_fd_sc_hd__nand2_1 _08352_ (.A(net813),
    .B(_02729_),
    .Y(_03364_));
 sky130_fd_sc_hd__a32o_1 _08353_ (.A1(_02728_),
    .A2(net431),
    .A3(_03364_),
    .B1(_02729_),
    .B2(net571),
    .X(_03365_));
 sky130_fd_sc_hd__a211o_1 _08354_ (.A1(_03175_),
    .A2(_03363_),
    .B1(_03365_),
    .C1(_03361_),
    .X(_03366_));
 sky130_fd_sc_hd__and3_1 _08355_ (.A(net245),
    .B(_03295_),
    .C(_03296_),
    .X(_03367_));
 sky130_fd_sc_hd__a21o_1 _08356_ (.A1(net240),
    .A2(_03275_),
    .B1(_03367_),
    .X(_03368_));
 sky130_fd_sc_hd__nor2_1 _08357_ (.A(net217),
    .B(_03368_),
    .Y(_03369_));
 sky130_fd_sc_hd__mux2_1 _08358_ (.A0(_03278_),
    .A1(_03283_),
    .S(net236),
    .X(_03370_));
 sky130_fd_sc_hd__a21o_1 _08359_ (.A1(net217),
    .A2(_03370_),
    .B1(net215),
    .X(_03371_));
 sky130_fd_sc_hd__and3_1 _08360_ (.A(net239),
    .B(_03286_),
    .C(_03287_),
    .X(_03372_));
 sky130_fd_sc_hd__a21oi_1 _08361_ (.A1(net245),
    .A2(_03234_),
    .B1(_03372_),
    .Y(_03373_));
 sky130_fd_sc_hd__and3_1 _08362_ (.A(net245),
    .B(_03288_),
    .C(_03289_),
    .X(_03374_));
 sky130_fd_sc_hd__a21oi_1 _08363_ (.A1(net240),
    .A2(_03294_),
    .B1(_03374_),
    .Y(_03375_));
 sky130_fd_sc_hd__mux2_1 _08364_ (.A0(_03373_),
    .A1(_03375_),
    .S(net218),
    .X(_03376_));
 sky130_fd_sc_hd__o22ai_1 _08365_ (.A1(_03369_),
    .A2(_03371_),
    .B1(_03376_),
    .B2(net206),
    .Y(_03377_));
 sky130_fd_sc_hd__a21oi_1 _08366_ (.A1(_02714_),
    .A2(_03318_),
    .B1(_03327_),
    .Y(_03378_));
 sky130_fd_sc_hd__xnor2_1 _08367_ (.A(_02733_),
    .B(_03378_),
    .Y(_03379_));
 sky130_fd_sc_hd__a22o_1 _08368_ (.A1(_03202_),
    .A2(_03377_),
    .B1(_03379_),
    .B2(net425),
    .X(_03380_));
 sky130_fd_sc_hd__a211o_1 _08369_ (.A1(net194),
    .A2(_03358_),
    .B1(_03366_),
    .C1(_03380_),
    .X(_03381_));
 sky130_fd_sc_hd__a22o_1 _08370_ (.A1(net1343),
    .A2(net566),
    .B1(_03381_),
    .B2(net740),
    .X(_00027_));
 sky130_fd_sc_hd__a211o_1 _08371_ (.A1(_02714_),
    .A2(_03318_),
    .B1(_03327_),
    .C1(_02729_),
    .X(_03382_));
 sky130_fd_sc_hd__a21oi_1 _08372_ (.A1(_02728_),
    .A2(_03382_),
    .B1(_02652_),
    .Y(_03383_));
 sky130_fd_sc_hd__a31o_1 _08373_ (.A1(_02652_),
    .A2(_02728_),
    .A3(_03382_),
    .B1(_03267_),
    .X(_03384_));
 sky130_fd_sc_hd__nor2_1 _08374_ (.A(_03383_),
    .B(_03384_),
    .Y(_03385_));
 sky130_fd_sc_hd__o21a_1 _08375_ (.A1(_03154_),
    .A2(_03157_),
    .B1(net225),
    .X(_03386_));
 sky130_fd_sc_hd__a21o_1 _08376_ (.A1(net227),
    .A2(_03150_),
    .B1(_03386_),
    .X(_03387_));
 sky130_fd_sc_hd__a211o_1 _08377_ (.A1(net228),
    .A2(_03150_),
    .B1(_03386_),
    .C1(net213),
    .X(_03388_));
 sky130_fd_sc_hd__a21o_1 _08378_ (.A1(net222),
    .A2(_03144_),
    .B1(net208),
    .X(_03389_));
 sky130_fd_sc_hd__and3_1 _08379_ (.A(_03255_),
    .B(_03388_),
    .C(_03389_),
    .X(_03390_));
 sky130_fd_sc_hd__a21oi_1 _08380_ (.A1(net225),
    .A2(_03144_),
    .B1(_03352_),
    .Y(_03391_));
 sky130_fd_sc_hd__o21bai_1 _08381_ (.A1(net213),
    .A2(_03387_),
    .B1_N(_03391_),
    .Y(_03392_));
 sky130_fd_sc_hd__and3b_1 _08382_ (.A_N(_03391_),
    .B(_03220_),
    .C(_03388_),
    .X(_03393_));
 sky130_fd_sc_hd__o21ai_1 _08383_ (.A1(_03390_),
    .A2(_03393_),
    .B1(net196),
    .Y(_03394_));
 sky130_fd_sc_hd__a31o_1 _08384_ (.A1(_02713_),
    .A2(_02730_),
    .A3(_03322_),
    .B1(_02731_),
    .X(_03395_));
 sky130_fd_sc_hd__a311o_1 _08385_ (.A1(_02713_),
    .A2(_02730_),
    .A3(_03322_),
    .B1(_02731_),
    .C1(_02652_),
    .X(_03396_));
 sky130_fd_sc_hd__a21oi_1 _08386_ (.A1(_02652_),
    .A2(_03395_),
    .B1(net426),
    .Y(_03397_));
 sky130_fd_sc_hd__mux2_1 _08387_ (.A0(_03163_),
    .A1(_03193_),
    .S(net220),
    .X(_03398_));
 sky130_fd_sc_hd__a31o_1 _08388_ (.A1(net226),
    .A2(_03198_),
    .A3(_03199_),
    .B1(net215),
    .X(_03399_));
 sky130_fd_sc_hd__a21o_1 _08389_ (.A1(net217),
    .A2(_03210_),
    .B1(_03399_),
    .X(_03400_));
 sky130_fd_sc_hd__o211a_1 _08390_ (.A1(net206),
    .A2(_03398_),
    .B1(_03400_),
    .C1(_03202_),
    .X(_03401_));
 sky130_fd_sc_hd__a21oi_1 _08391_ (.A1(_02650_),
    .A2(net188),
    .B1(_03205_),
    .Y(_03402_));
 sky130_fd_sc_hd__mux2_1 _08392_ (.A0(_03325_),
    .A1(_03402_),
    .S(net237),
    .X(_03403_));
 sky130_fd_sc_hd__mux2_2 _08393_ (.A0(_02700_),
    .A1(_03403_),
    .S(net218),
    .X(_03404_));
 sky130_fd_sc_hd__nor2_1 _08394_ (.A(net193),
    .B(_02650_),
    .Y(_03405_));
 sky130_fd_sc_hd__nor2_1 _08395_ (.A(_02650_),
    .B(_03185_),
    .Y(_03406_));
 sky130_fd_sc_hd__a221o_1 _08396_ (.A1(_03180_),
    .A2(_03404_),
    .B1(_03405_),
    .B2(net571),
    .C1(_03406_),
    .X(_03407_));
 sky130_fd_sc_hd__a211oi_1 _08397_ (.A1(_02652_),
    .A2(net431),
    .B1(_03401_),
    .C1(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__a21oi_1 _08398_ (.A1(_03396_),
    .A2(_03397_),
    .B1(_03385_),
    .Y(_03409_));
 sky130_fd_sc_hd__and3_1 _08399_ (.A(_03394_),
    .B(_03408_),
    .C(_03409_),
    .X(_03410_));
 sky130_fd_sc_hd__a2bb2o_1 _08400_ (.A1_N(_02575_),
    .A2_N(_03410_),
    .B1(net566),
    .B2(net1324),
    .X(_00028_));
 sky130_fd_sc_hd__a31o_1 _08401_ (.A1(_02652_),
    .A2(_02728_),
    .A3(_03382_),
    .B1(_03405_),
    .X(_03411_));
 sky130_fd_sc_hd__a21oi_1 _08402_ (.A1(_02669_),
    .A2(_03411_),
    .B1(_03267_),
    .Y(_03412_));
 sky130_fd_sc_hd__o21a_1 _08403_ (.A1(_02669_),
    .A2(_03411_),
    .B1(_03412_),
    .X(_03413_));
 sky130_fd_sc_hd__and3_1 _08404_ (.A(net228),
    .B(_03241_),
    .C(_03242_),
    .X(_03414_));
 sky130_fd_sc_hd__and3_1 _08405_ (.A(net224),
    .B(_03226_),
    .C(_03227_),
    .X(_03415_));
 sky130_fd_sc_hd__or3_1 _08406_ (.A(net212),
    .B(_03414_),
    .C(_03415_),
    .X(_03416_));
 sky130_fd_sc_hd__a21o_1 _08407_ (.A1(_03247_),
    .A2(_03252_),
    .B1(net227),
    .X(_03417_));
 sky130_fd_sc_hd__nand2_1 _08408_ (.A(net211),
    .B(_03417_),
    .Y(_03418_));
 sky130_fd_sc_hd__and3_1 _08409_ (.A(_03255_),
    .B(_03416_),
    .C(_03418_),
    .X(_03419_));
 sky130_fd_sc_hd__o21a_1 _08410_ (.A1(_03246_),
    .A2(_03248_),
    .B1(net222),
    .X(_03420_));
 sky130_fd_sc_hd__o32a_1 _08411_ (.A1(net212),
    .A2(_03414_),
    .A3(_03415_),
    .B1(_03420_),
    .B2(_03352_),
    .X(_03421_));
 sky130_fd_sc_hd__a32o_1 _08412_ (.A1(_03255_),
    .A2(_03416_),
    .A3(_03418_),
    .B1(_03421_),
    .B2(_03220_),
    .X(_03422_));
 sky130_fd_sc_hd__a21oi_1 _08413_ (.A1(_02659_),
    .A2(net187),
    .B1(_03282_),
    .Y(_03423_));
 sky130_fd_sc_hd__mux2_1 _08414_ (.A0(_03362_),
    .A1(_03423_),
    .S(net238),
    .X(_03424_));
 sky130_fd_sc_hd__mux2_2 _08415_ (.A0(_03271_),
    .A1(_03424_),
    .S(net216),
    .X(_03425_));
 sky130_fd_sc_hd__o211a_1 _08416_ (.A1(net846),
    .A2(_02667_),
    .B1(_02668_),
    .C1(net431),
    .X(_03426_));
 sky130_fd_sc_hd__a221o_1 _08417_ (.A1(_02666_),
    .A2(net571),
    .B1(_03180_),
    .B2(_03425_),
    .C1(_03426_),
    .X(_03427_));
 sky130_fd_sc_hd__a211o_1 _08418_ (.A1(net245),
    .A2(_03294_),
    .B1(_03297_),
    .C1(net218),
    .X(_03428_));
 sky130_fd_sc_hd__o211a_1 _08419_ (.A1(net226),
    .A2(_03279_),
    .B1(_03428_),
    .C1(net206),
    .X(_03429_));
 sky130_fd_sc_hd__a311o_1 _08420_ (.A1(net245),
    .A2(_03286_),
    .A3(_03287_),
    .B1(_03290_),
    .C1(net226),
    .X(_03430_));
 sky130_fd_sc_hd__o21a_1 _08421_ (.A1(net220),
    .A2(_03235_),
    .B1(_03430_),
    .X(_03431_));
 sky130_fd_sc_hd__o211a_1 _08422_ (.A1(net219),
    .A2(_03235_),
    .B1(_03430_),
    .C1(net210),
    .X(_03432_));
 sky130_fd_sc_hd__o21a_1 _08423_ (.A1(_03429_),
    .A2(_03432_),
    .B1(_03202_),
    .X(_03433_));
 sky130_fd_sc_hd__a211o_1 _08424_ (.A1(net194),
    .A2(_03422_),
    .B1(_03427_),
    .C1(_03433_),
    .X(_03434_));
 sky130_fd_sc_hd__a21o_1 _08425_ (.A1(_02651_),
    .A2(_03396_),
    .B1(_02669_),
    .X(_03435_));
 sky130_fd_sc_hd__a31oi_1 _08426_ (.A1(_02651_),
    .A2(_02669_),
    .A3(_03396_),
    .B1(net426),
    .Y(_03436_));
 sky130_fd_sc_hd__a211o_1 _08427_ (.A1(_03435_),
    .A2(_03436_),
    .B1(_03413_),
    .C1(_03434_),
    .X(_03437_));
 sky130_fd_sc_hd__a22o_1 _08428_ (.A1(net1326),
    .A2(net566),
    .B1(_03437_),
    .B2(net740),
    .X(_00029_));
 sky130_fd_sc_hd__and2_1 _08429_ (.A(_02651_),
    .B(_02664_),
    .X(_03438_));
 sky130_fd_sc_hd__nor2_1 _08430_ (.A(_02665_),
    .B(_03438_),
    .Y(_03439_));
 sky130_fd_sc_hd__nor2_1 _08431_ (.A(_02669_),
    .B(_03396_),
    .Y(_03440_));
 sky130_fd_sc_hd__a211o_1 _08432_ (.A1(_03396_),
    .A2(_03438_),
    .B1(_02620_),
    .C1(_02665_),
    .X(_03441_));
 sky130_fd_sc_hd__o311a_1 _08433_ (.A1(_02621_),
    .A2(_03439_),
    .A3(_03440_),
    .B1(_03441_),
    .C1(net428),
    .X(_03442_));
 sky130_fd_sc_hd__nand4_2 _08434_ (.A(_02652_),
    .B(_02669_),
    .C(_02728_),
    .D(_03382_),
    .Y(_03443_));
 sky130_fd_sc_hd__a21oi_1 _08435_ (.A1(_02668_),
    .A2(_03405_),
    .B1(_02666_),
    .Y(_03444_));
 sky130_fd_sc_hd__a21oi_1 _08436_ (.A1(_03443_),
    .A2(_03444_),
    .B1(_02621_),
    .Y(_03445_));
 sky130_fd_sc_hd__a31o_1 _08437_ (.A1(_02621_),
    .A2(_03443_),
    .A3(_03444_),
    .B1(_03267_),
    .X(_03446_));
 sky130_fd_sc_hd__nor2_1 _08438_ (.A(_03445_),
    .B(_03446_),
    .Y(_03447_));
 sky130_fd_sc_hd__o211a_1 _08439_ (.A1(net243),
    .A2(_03141_),
    .B1(_03310_),
    .C1(net227),
    .X(_03448_));
 sky130_fd_sc_hd__and3_1 _08440_ (.A(net224),
    .B(_03303_),
    .C(_03304_),
    .X(_03449_));
 sky130_fd_sc_hd__or2_1 _08441_ (.A(_03448_),
    .B(_03449_),
    .X(_03450_));
 sky130_fd_sc_hd__or3_1 _08442_ (.A(net211),
    .B(_03448_),
    .C(_03449_),
    .X(_03451_));
 sky130_fd_sc_hd__a2111o_1 _08443_ (.A1(net199),
    .A2(net190),
    .B1(net227),
    .C1(_03142_),
    .D1(net247),
    .X(_03452_));
 sky130_fd_sc_hd__nand2_1 _08444_ (.A(net214),
    .B(_03452_),
    .Y(_03453_));
 sky130_fd_sc_hd__o31a_1 _08445_ (.A1(net214),
    .A2(_03448_),
    .A3(_03449_),
    .B1(_03453_),
    .X(_03454_));
 sky130_fd_sc_hd__a21oi_1 _08446_ (.A1(net243),
    .A2(net222),
    .B1(net198),
    .Y(_03455_));
 sky130_fd_sc_hd__a31o_1 _08447_ (.A1(net688),
    .A2(_03451_),
    .A3(_03455_),
    .B1(_03454_),
    .X(_03456_));
 sky130_fd_sc_hd__a211o_1 _08448_ (.A1(net239),
    .A2(_03160_),
    .B1(_03305_),
    .C1(net219),
    .X(_03457_));
 sky130_fd_sc_hd__o21a_1 _08449_ (.A1(net226),
    .A2(_03336_),
    .B1(_03457_),
    .X(_03458_));
 sky130_fd_sc_hd__and2_1 _08450_ (.A(net217),
    .B(_03333_),
    .X(_03459_));
 sky130_fd_sc_hd__a21o_1 _08451_ (.A1(_02707_),
    .A2(_03338_),
    .B1(net215),
    .X(_03460_));
 sky130_fd_sc_hd__o221a_1 _08452_ (.A1(net206),
    .A2(_03458_),
    .B1(_03459_),
    .B2(_03460_),
    .C1(_03202_),
    .X(_03461_));
 sky130_fd_sc_hd__a21oi_1 _08453_ (.A1(_02609_),
    .A2(net187),
    .B1(_03208_),
    .Y(_03462_));
 sky130_fd_sc_hd__mux2_1 _08454_ (.A0(_03402_),
    .A1(_03462_),
    .S(net236),
    .X(_03463_));
 sky130_fd_sc_hd__mux2_1 _08455_ (.A0(_03326_),
    .A1(_03463_),
    .S(net219),
    .X(_03464_));
 sky130_fd_sc_hd__o211a_1 _08456_ (.A1(net845),
    .A2(_02616_),
    .B1(_02617_),
    .C1(net431),
    .X(_03465_));
 sky130_fd_sc_hd__a221o_1 _08457_ (.A1(_02615_),
    .A2(net571),
    .B1(_03180_),
    .B2(_03464_),
    .C1(_03465_),
    .X(_03466_));
 sky130_fd_sc_hd__a31o_1 _08458_ (.A1(net194),
    .A2(net573),
    .A3(_03456_),
    .B1(_03466_),
    .X(_03467_));
 sky130_fd_sc_hd__or4_2 _08459_ (.A(_03442_),
    .B(_03447_),
    .C(_03461_),
    .D(_03467_),
    .X(_03468_));
 sky130_fd_sc_hd__a22o_1 _08460_ (.A1(net1309),
    .A2(net566),
    .B1(_03468_),
    .B2(net740),
    .X(_00030_));
 sky130_fd_sc_hd__a21oi_1 _08461_ (.A1(_02619_),
    .A2(_03441_),
    .B1(_02638_),
    .Y(_03469_));
 sky130_fd_sc_hd__a311oi_1 _08462_ (.A1(_02619_),
    .A2(_02638_),
    .A3(_03441_),
    .B1(_03469_),
    .C1(net426),
    .Y(_03470_));
 sky130_fd_sc_hd__or3_1 _08463_ (.A(_02615_),
    .B(_02638_),
    .C(_03445_),
    .X(_03471_));
 sky130_fd_sc_hd__o21ai_1 _08464_ (.A1(_02615_),
    .A2(_03445_),
    .B1(_02638_),
    .Y(_03472_));
 sky130_fd_sc_hd__and3_1 _08465_ (.A(net423),
    .B(_03471_),
    .C(_03472_),
    .X(_03473_));
 sky130_fd_sc_hd__a21o_1 _08466_ (.A1(_03342_),
    .A2(_03343_),
    .B1(net228),
    .X(_03474_));
 sky130_fd_sc_hd__a21o_1 _08467_ (.A1(_03348_),
    .A2(_03349_),
    .B1(net224),
    .X(_03475_));
 sky130_fd_sc_hd__a21oi_1 _08468_ (.A1(_03474_),
    .A2(_03475_),
    .B1(net212),
    .Y(_03476_));
 sky130_fd_sc_hd__nand2_1 _08469_ (.A(net223),
    .B(_03354_),
    .Y(_03477_));
 sky130_fd_sc_hd__a211oi_1 _08470_ (.A1(net211),
    .A2(_03477_),
    .B1(_03476_),
    .C1(_03256_),
    .Y(_03478_));
 sky130_fd_sc_hd__a21oi_1 _08471_ (.A1(net198),
    .A2(net211),
    .B1(_03476_),
    .Y(_03479_));
 sky130_fd_sc_hd__a21o_1 _08472_ (.A1(_03220_),
    .A2(_03479_),
    .B1(_03478_),
    .X(_03480_));
 sky130_fd_sc_hd__a21oi_1 _08473_ (.A1(_02627_),
    .A2(net187),
    .B1(_03277_),
    .Y(_03481_));
 sky130_fd_sc_hd__mux2_1 _08474_ (.A0(_03423_),
    .A1(_03481_),
    .S(net238),
    .X(_03482_));
 sky130_fd_sc_hd__mux2_2 _08475_ (.A0(_03363_),
    .A1(_03482_),
    .S(net221),
    .X(_03483_));
 sky130_fd_sc_hd__o211a_1 _08476_ (.A1(net845),
    .A2(_02634_),
    .B1(_02635_),
    .C1(net430),
    .X(_03484_));
 sky130_fd_sc_hd__a221o_1 _08477_ (.A1(_02633_),
    .A2(net571),
    .B1(_03180_),
    .B2(_03483_),
    .C1(_03484_),
    .X(_03485_));
 sky130_fd_sc_hd__a211o_1 _08478_ (.A1(net242),
    .A2(_03231_),
    .B1(_03344_),
    .C1(net225),
    .X(_03486_));
 sky130_fd_sc_hd__a21boi_2 _08479_ (.A1(net220),
    .A2(_03373_),
    .B1_N(_03486_),
    .Y(_03487_));
 sky130_fd_sc_hd__nor2_1 _08480_ (.A(net218),
    .B(_03375_),
    .Y(_03488_));
 sky130_fd_sc_hd__a211o_1 _08481_ (.A1(net218),
    .A2(_03368_),
    .B1(_03488_),
    .C1(net215),
    .X(_03489_));
 sky130_fd_sc_hd__o211a_1 _08482_ (.A1(net207),
    .A2(_03487_),
    .B1(_03489_),
    .C1(_03202_),
    .X(_03490_));
 sky130_fd_sc_hd__a211o_1 _08483_ (.A1(net195),
    .A2(_03480_),
    .B1(_03485_),
    .C1(_03490_),
    .X(_03491_));
 sky130_fd_sc_hd__or3_2 _08484_ (.A(_03470_),
    .B(_03473_),
    .C(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__a22o_1 _08485_ (.A1(net1349),
    .A2(net566),
    .B1(_03492_),
    .B2(net740),
    .X(_00031_));
 sky130_fd_sc_hd__nand2_1 _08486_ (.A(_02615_),
    .B(_02635_),
    .Y(_03493_));
 sky130_fd_sc_hd__and3_1 _08487_ (.A(_02634_),
    .B(_03444_),
    .C(_03493_),
    .X(_03494_));
 sky130_fd_sc_hd__o21ai_1 _08488_ (.A1(_02617_),
    .A2(_02633_),
    .B1(_02635_),
    .Y(_03495_));
 sky130_fd_sc_hd__a21oi_2 _08489_ (.A1(_03443_),
    .A2(_03494_),
    .B1(_03495_),
    .Y(_03496_));
 sky130_fd_sc_hd__xnor2_1 _08490_ (.A(_03092_),
    .B(_03496_),
    .Y(_03497_));
 sky130_fd_sc_hd__a311o_1 _08491_ (.A1(_02713_),
    .A2(_02730_),
    .A3(_03322_),
    .B1(_02731_),
    .C1(_02670_),
    .X(_03498_));
 sky130_fd_sc_hd__o21ai_1 _08492_ (.A1(_02618_),
    .A2(_02637_),
    .B1(_02636_),
    .Y(_03499_));
 sky130_fd_sc_hd__o31a_1 _08493_ (.A1(_02639_),
    .A2(_02665_),
    .A3(_03438_),
    .B1(_03499_),
    .X(_03500_));
 sky130_fd_sc_hd__nand2_1 _08494_ (.A(_03498_),
    .B(_03500_),
    .Y(_03501_));
 sky130_fd_sc_hd__and2_1 _08495_ (.A(_03092_),
    .B(_03501_),
    .X(_03502_));
 sky130_fd_sc_hd__a31o_1 _08496_ (.A1(_03091_),
    .A2(_03498_),
    .A3(_03500_),
    .B1(net426),
    .X(_03503_));
 sky130_fd_sc_hd__o21a_1 _08497_ (.A1(_02628_),
    .A2(net188),
    .B1(_03197_),
    .X(_03504_));
 sky130_fd_sc_hd__mux2_1 _08498_ (.A0(_03462_),
    .A1(_03504_),
    .S(net237),
    .X(_03505_));
 sky130_fd_sc_hd__mux2_1 _08499_ (.A0(_03403_),
    .A1(_03505_),
    .S(net217),
    .X(_03506_));
 sky130_fd_sc_hd__nor2_1 _08500_ (.A(net207),
    .B(_03171_),
    .Y(_03507_));
 sky130_fd_sc_hd__a32o_1 _08501_ (.A1(_02700_),
    .A2(net216),
    .A3(_03507_),
    .B1(_03506_),
    .B2(_03178_),
    .X(_03508_));
 sky130_fd_sc_hd__a211o_1 _08502_ (.A1(net226),
    .A2(_03193_),
    .B1(_03200_),
    .C1(net210),
    .X(_03509_));
 sky130_fd_sc_hd__o211a_1 _08503_ (.A1(net206),
    .A2(_03164_),
    .B1(_03509_),
    .C1(_03138_),
    .X(_03510_));
 sky130_fd_sc_hd__o21a_1 _08504_ (.A1(_03508_),
    .A2(_03510_),
    .B1(net193),
    .X(_03511_));
 sky130_fd_sc_hd__nor2_4 _08505_ (.A(net846),
    .B(_03183_),
    .Y(_03512_));
 sky130_fd_sc_hd__nand2_2 _08506_ (.A(net813),
    .B(net430),
    .Y(_03513_));
 sky130_fd_sc_hd__nor2_1 _08507_ (.A(_03088_),
    .B(_03185_),
    .Y(_03514_));
 sky130_fd_sc_hd__a221o_1 _08508_ (.A1(_03087_),
    .A2(net570),
    .B1(_03512_),
    .B2(_03091_),
    .C1(_03514_),
    .X(_03515_));
 sky130_fd_sc_hd__nor2_1 _08509_ (.A(net198),
    .B(net208),
    .Y(_03516_));
 sky130_fd_sc_hd__a22o_1 _08510_ (.A1(net207),
    .A2(_03151_),
    .B1(_03516_),
    .B2(net688),
    .X(_03517_));
 sky130_fd_sc_hd__a31o_1 _08511_ (.A1(net195),
    .A2(net573),
    .A3(_03517_),
    .B1(_03515_),
    .X(_03518_));
 sky130_fd_sc_hd__a211o_1 _08512_ (.A1(net423),
    .A2(_03497_),
    .B1(_03511_),
    .C1(_03518_),
    .X(_03519_));
 sky130_fd_sc_hd__o21bai_1 _08513_ (.A1(_03502_),
    .A2(_03503_),
    .B1_N(_03519_),
    .Y(_03520_));
 sky130_fd_sc_hd__a22o_1 _08514_ (.A1(net1328),
    .A2(net566),
    .B1(_03520_),
    .B2(net740),
    .X(_00032_));
 sky130_fd_sc_hd__a21oi_1 _08515_ (.A1(_03091_),
    .A2(_03496_),
    .B1(_03087_),
    .Y(_03521_));
 sky130_fd_sc_hd__a211o_1 _08516_ (.A1(_03091_),
    .A2(_03496_),
    .B1(_03075_),
    .C1(_03087_),
    .X(_03522_));
 sky130_fd_sc_hd__nor2_1 _08517_ (.A(_03074_),
    .B(_03092_),
    .Y(_03523_));
 sky130_fd_sc_hd__o211a_1 _08518_ (.A1(_03074_),
    .A2(_03521_),
    .B1(_03522_),
    .C1(net423),
    .X(_03524_));
 sky130_fd_sc_hd__mux2_1 _08519_ (.A0(_03236_),
    .A1(_03299_),
    .S(net206),
    .X(_03525_));
 sky130_fd_sc_hd__and2b_1 _08520_ (.A_N(_03274_),
    .B(_03296_),
    .X(_03526_));
 sky130_fd_sc_hd__mux2_1 _08521_ (.A0(_03481_),
    .A1(_03526_),
    .S(net238),
    .X(_03527_));
 sky130_fd_sc_hd__mux2_1 _08522_ (.A0(_03424_),
    .A1(_03527_),
    .S(net221),
    .X(_03528_));
 sky130_fd_sc_hd__a32o_1 _08523_ (.A1(net216),
    .A2(_03271_),
    .A3(net185),
    .B1(_03528_),
    .B2(net186),
    .X(_03529_));
 sky130_fd_sc_hd__nand2_2 _08524_ (.A(net208),
    .B(_03255_),
    .Y(_03530_));
 sky130_fd_sc_hd__nand3b_1 _08525_ (.A_N(_03530_),
    .B(_03253_),
    .C(_03243_),
    .Y(_03531_));
 sky130_fd_sc_hd__inv_2 _08526_ (.A(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__a31o_1 _08527_ (.A1(net208),
    .A2(_03243_),
    .A3(_03249_),
    .B1(_03516_),
    .X(_03533_));
 sky130_fd_sc_hd__o211a_1 _08528_ (.A1(net846),
    .A2(_03072_),
    .B1(_03073_),
    .C1(net430),
    .X(_03534_));
 sky130_fd_sc_hd__nor2_1 _08529_ (.A(_03072_),
    .B(_03170_),
    .Y(_03535_));
 sky130_fd_sc_hd__a211o_1 _08530_ (.A1(_03220_),
    .A2(_03533_),
    .B1(_03532_),
    .C1(net191),
    .X(_03536_));
 sky130_fd_sc_hd__a211o_1 _08531_ (.A1(_03138_),
    .A2(_03525_),
    .B1(_03529_),
    .C1(net195),
    .X(_03537_));
 sky130_fd_sc_hd__a211oi_1 _08532_ (.A1(_03536_),
    .A2(_03537_),
    .B1(_03534_),
    .C1(_03535_),
    .Y(_03538_));
 sky130_fd_sc_hd__a211o_1 _08533_ (.A1(_03498_),
    .A2(_03500_),
    .B1(_03075_),
    .C1(_03091_),
    .X(_03539_));
 sky130_fd_sc_hd__o211a_1 _08534_ (.A1(_03075_),
    .A2(_03090_),
    .B1(net428),
    .C1(_03539_),
    .X(_03540_));
 sky130_fd_sc_hd__o31a_1 _08535_ (.A1(_03074_),
    .A2(_03089_),
    .A3(_03502_),
    .B1(_03540_),
    .X(_03541_));
 sky130_fd_sc_hd__or3b_1 _08536_ (.A(_03524_),
    .B(_03541_),
    .C_N(_03538_),
    .X(_03542_));
 sky130_fd_sc_hd__a22o_1 _08537_ (.A1(net1303),
    .A2(net566),
    .B1(_03542_),
    .B2(net740),
    .X(_00033_));
 sky130_fd_sc_hd__o31a_1 _08538_ (.A1(_03074_),
    .A2(_03080_),
    .A3(_03086_),
    .B1(_03072_),
    .X(_03543_));
 sky130_fd_sc_hd__a21bo_1 _08539_ (.A1(_03496_),
    .A2(_03523_),
    .B1_N(_03543_),
    .X(_03544_));
 sky130_fd_sc_hd__a21oi_1 _08540_ (.A1(_03042_),
    .A2(_03544_),
    .B1(_03267_),
    .Y(_03545_));
 sky130_fd_sc_hd__o21a_1 _08541_ (.A1(_03042_),
    .A2(_03544_),
    .B1(_03545_),
    .X(_03546_));
 sky130_fd_sc_hd__a21oi_1 _08542_ (.A1(_03074_),
    .A2(_03089_),
    .B1(_03071_),
    .Y(_03547_));
 sky130_fd_sc_hd__and3_1 _08543_ (.A(_03042_),
    .B(_03539_),
    .C(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__a21oi_1 _08544_ (.A1(_03539_),
    .A2(_03547_),
    .B1(_03042_),
    .Y(_03549_));
 sky130_fd_sc_hd__or3_1 _08545_ (.A(net426),
    .B(_03548_),
    .C(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__a21oi_1 _08546_ (.A1(_03312_),
    .A2(_03314_),
    .B1(net211),
    .Y(_03551_));
 sky130_fd_sc_hd__o21a_1 _08547_ (.A1(_03516_),
    .A2(_03551_),
    .B1(_03220_),
    .X(_03552_));
 sky130_fd_sc_hd__or2_1 _08548_ (.A(_03312_),
    .B(_03530_),
    .X(_03553_));
 sky130_fd_sc_hd__nand2_1 _08549_ (.A(net196),
    .B(_03553_),
    .Y(_03554_));
 sky130_fd_sc_hd__a21o_1 _08550_ (.A1(_03306_),
    .A2(_03307_),
    .B1(net209),
    .X(_03555_));
 sky130_fd_sc_hd__o211a_1 _08551_ (.A1(net213),
    .A2(_03339_),
    .B1(_03555_),
    .C1(net573),
    .X(_03556_));
 sky130_fd_sc_hd__and2_1 _08552_ (.A(_03195_),
    .B(_03196_),
    .X(_03557_));
 sky130_fd_sc_hd__mux2_1 _08553_ (.A0(_03504_),
    .A1(_03557_),
    .S(net240),
    .X(_03558_));
 sky130_fd_sc_hd__mux2_1 _08554_ (.A0(_03463_),
    .A1(_03558_),
    .S(net219),
    .X(_03559_));
 sky130_fd_sc_hd__a32o_1 _08555_ (.A1(net216),
    .A2(_03326_),
    .A3(net185),
    .B1(_03559_),
    .B2(net186),
    .X(_03560_));
 sky130_fd_sc_hd__o32a_1 _08556_ (.A1(net196),
    .A2(_03556_),
    .A3(_03560_),
    .B1(_03552_),
    .B2(_03554_),
    .X(_03561_));
 sky130_fd_sc_hd__nand2_1 _08557_ (.A(net813),
    .B(_03041_),
    .Y(_03562_));
 sky130_fd_sc_hd__o21a_1 _08558_ (.A1(_03035_),
    .A2(_03040_),
    .B1(net430),
    .X(_03563_));
 sky130_fd_sc_hd__a221o_1 _08559_ (.A1(_03041_),
    .A2(net570),
    .B1(_03562_),
    .B2(_03563_),
    .C1(_03561_),
    .X(_03564_));
 sky130_fd_sc_hd__or3b_2 _08560_ (.A(_03546_),
    .B(_03564_),
    .C_N(_03550_),
    .X(_03565_));
 sky130_fd_sc_hd__a22o_1 _08561_ (.A1(net1319),
    .A2(net566),
    .B1(_03565_),
    .B2(net740),
    .X(_00003_));
 sky130_fd_sc_hd__a21oi_1 _08562_ (.A1(_03042_),
    .A2(_03544_),
    .B1(_03041_),
    .Y(_03566_));
 sky130_fd_sc_hd__a211o_1 _08563_ (.A1(_03042_),
    .A2(_03544_),
    .B1(_03057_),
    .C1(_03041_),
    .X(_03567_));
 sky130_fd_sc_hd__o211a_1 _08564_ (.A1(_03058_),
    .A2(_03566_),
    .B1(_03567_),
    .C1(net423),
    .X(_03568_));
 sky130_fd_sc_hd__o21a_1 _08565_ (.A1(_03038_),
    .A2(_03039_),
    .B1(_03035_),
    .X(_03569_));
 sky130_fd_sc_hd__or3_1 _08566_ (.A(_03058_),
    .B(_03549_),
    .C(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__o21ai_1 _08567_ (.A1(_03549_),
    .A2(_03569_),
    .B1(_03058_),
    .Y(_03571_));
 sky130_fd_sc_hd__and3_1 _08568_ (.A(net428),
    .B(_03570_),
    .C(_03571_),
    .X(_03572_));
 sky130_fd_sc_hd__and2_1 _08569_ (.A(_03293_),
    .B(_03295_),
    .X(_03573_));
 sky130_fd_sc_hd__mux2_1 _08570_ (.A0(_03526_),
    .A1(_03573_),
    .S(net239),
    .X(_03574_));
 sky130_fd_sc_hd__mux2_1 _08571_ (.A0(_03482_),
    .A1(_03574_),
    .S(net216),
    .X(_03575_));
 sky130_fd_sc_hd__and3_1 _08572_ (.A(net222),
    .B(_03363_),
    .C(_03507_),
    .X(_03576_));
 sky130_fd_sc_hd__a21oi_1 _08573_ (.A1(_03178_),
    .A2(_03575_),
    .B1(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__a21oi_1 _08574_ (.A1(_03345_),
    .A2(_03346_),
    .B1(net209),
    .Y(_03578_));
 sky130_fd_sc_hd__a211o_1 _08575_ (.A1(net209),
    .A2(_03376_),
    .B1(_03578_),
    .C1(_03139_),
    .X(_03579_));
 sky130_fd_sc_hd__o211a_1 _08576_ (.A1(net845),
    .A2(_03053_),
    .B1(_03054_),
    .C1(net430),
    .X(_03580_));
 sky130_fd_sc_hd__a21oi_1 _08577_ (.A1(net223),
    .A2(net209),
    .B1(net198),
    .Y(_03581_));
 sky130_fd_sc_hd__o21ba_1 _08578_ (.A1(net211),
    .A2(_03350_),
    .B1_N(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__nand2b_1 _08579_ (.A_N(_03530_),
    .B(_03355_),
    .Y(_03583_));
 sky130_fd_sc_hd__o211a_1 _08580_ (.A1(_03221_),
    .A2(_03582_),
    .B1(_03583_),
    .C1(net196),
    .X(_03584_));
 sky130_fd_sc_hd__a31o_1 _08581_ (.A1(net192),
    .A2(_03577_),
    .A3(_03579_),
    .B1(_03584_),
    .X(_03585_));
 sky130_fd_sc_hd__o21ai_1 _08582_ (.A1(_03053_),
    .A2(_03170_),
    .B1(_03585_),
    .Y(_03586_));
 sky130_fd_sc_hd__or4_2 _08583_ (.A(_03568_),
    .B(_03572_),
    .C(_03580_),
    .D(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__a22o_1 _08584_ (.A1(net1314),
    .A2(net567),
    .B1(_03587_),
    .B2(net742),
    .X(_00004_));
 sky130_fd_sc_hd__nand2_1 _08585_ (.A(_03042_),
    .B(_03057_),
    .Y(_03588_));
 sky130_fd_sc_hd__a21boi_1 _08586_ (.A1(_03041_),
    .A2(_03054_),
    .B1_N(_03053_),
    .Y(_03589_));
 sky130_fd_sc_hd__o21ai_1 _08587_ (.A1(_03543_),
    .A2(_03588_),
    .B1(_03589_),
    .Y(_03590_));
 sky130_fd_sc_hd__and3b_1 _08588_ (.A_N(_03588_),
    .B(_03075_),
    .C(_03091_),
    .X(_03591_));
 sky130_fd_sc_hd__a21o_1 _08589_ (.A1(_03496_),
    .A2(_03591_),
    .B1(_03590_),
    .X(_03592_));
 sky130_fd_sc_hd__nor2_1 _08590_ (.A(_03026_),
    .B(_03592_),
    .Y(_03593_));
 sky130_fd_sc_hd__a21o_1 _08591_ (.A1(_03026_),
    .A2(_03592_),
    .B1(_03267_),
    .X(_03594_));
 sky130_fd_sc_hd__a21o_1 _08592_ (.A1(_03498_),
    .A2(_03500_),
    .B1(_03093_),
    .X(_03595_));
 sky130_fd_sc_hd__a21oi_1 _08593_ (.A1(_03056_),
    .A2(_03569_),
    .B1(_03055_),
    .Y(_03596_));
 sky130_fd_sc_hd__o21a_1 _08594_ (.A1(_03059_),
    .A2(_03547_),
    .B1(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__a21oi_1 _08595_ (.A1(_03595_),
    .A2(_03597_),
    .B1(_03026_),
    .Y(_03598_));
 sky130_fd_sc_hd__a311o_1 _08596_ (.A1(_03026_),
    .A2(_03595_),
    .A3(_03597_),
    .B1(_03598_),
    .C1(net426),
    .X(_03599_));
 sky130_fd_sc_hd__o21a_1 _08597_ (.A1(net190),
    .A2(_03018_),
    .B1(_03194_),
    .X(_03600_));
 sky130_fd_sc_hd__mux2_1 _08598_ (.A0(_03557_),
    .A1(_03600_),
    .S(net239),
    .X(_03601_));
 sky130_fd_sc_hd__mux2_1 _08599_ (.A0(_03505_),
    .A1(_03601_),
    .S(net217),
    .X(_03602_));
 sky130_fd_sc_hd__a22o_1 _08600_ (.A1(_03404_),
    .A2(net185),
    .B1(_03602_),
    .B2(net186),
    .X(_03603_));
 sky130_fd_sc_hd__mux2_1 _08601_ (.A0(_03387_),
    .A1(_03398_),
    .S(net206),
    .X(_03604_));
 sky130_fd_sc_hd__a21o_1 _08602_ (.A1(net573),
    .A2(_03604_),
    .B1(_03603_),
    .X(_03605_));
 sky130_fd_sc_hd__nor2_1 _08603_ (.A(_03024_),
    .B(_03185_),
    .Y(_03606_));
 sky130_fd_sc_hd__a221o_1 _08604_ (.A1(_03025_),
    .A2(net570),
    .B1(_03512_),
    .B2(_03026_),
    .C1(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__a32o_1 _08605_ (.A1(net222),
    .A2(net208),
    .A3(_03144_),
    .B1(_03581_),
    .B2(net688),
    .X(_03608_));
 sky130_fd_sc_hd__a31o_1 _08606_ (.A1(net194),
    .A2(net573),
    .A3(_03608_),
    .B1(_03607_),
    .X(_03609_));
 sky130_fd_sc_hd__a21oi_1 _08607_ (.A1(net193),
    .A2(_03605_),
    .B1(_03609_),
    .Y(_03610_));
 sky130_fd_sc_hd__o211ai_2 _08608_ (.A1(_03593_),
    .A2(_03594_),
    .B1(_03599_),
    .C1(_03610_),
    .Y(_03611_));
 sky130_fd_sc_hd__nor3b_4 _08609_ (.A(net951),
    .B(\alu.r_type ),
    .C_N(\dec.op_lui ),
    .Y(_03612_));
 sky130_fd_sc_hd__and3_1 _08610_ (.A(net847),
    .B(net766),
    .C(net757),
    .X(_03613_));
 sky130_fd_sc_hd__a221o_1 _08611_ (.A1(net1311),
    .A2(net567),
    .B1(_03611_),
    .B2(net742),
    .C1(_03613_),
    .X(_00005_));
 sky130_fd_sc_hd__a21oi_1 _08612_ (.A1(_03026_),
    .A2(_03592_),
    .B1(_03025_),
    .Y(_03614_));
 sky130_fd_sc_hd__and2b_1 _08613_ (.A_N(_03012_),
    .B(_03026_),
    .X(_03615_));
 sky130_fd_sc_hd__nand2b_1 _08614_ (.A_N(_03012_),
    .B(_03025_),
    .Y(_03616_));
 sky130_fd_sc_hd__nand2_1 _08615_ (.A(net423),
    .B(_03616_),
    .Y(_03617_));
 sky130_fd_sc_hd__a21o_1 _08616_ (.A1(_03592_),
    .A2(_03615_),
    .B1(_03617_),
    .X(_03618_));
 sky130_fd_sc_hd__a21o_1 _08617_ (.A1(_03012_),
    .A2(_03614_),
    .B1(_03618_),
    .X(_03619_));
 sky130_fd_sc_hd__a21o_1 _08618_ (.A1(_03018_),
    .A2(_03023_),
    .B1(_03598_),
    .X(_03620_));
 sky130_fd_sc_hd__nor2_1 _08619_ (.A(_03012_),
    .B(_03620_),
    .Y(_03621_));
 sky130_fd_sc_hd__a21o_1 _08620_ (.A1(_03012_),
    .A2(_03620_),
    .B1(net426),
    .X(_03622_));
 sky130_fd_sc_hd__and2_1 _08621_ (.A(_03289_),
    .B(_03292_),
    .X(_03623_));
 sky130_fd_sc_hd__mux2_1 _08622_ (.A0(_03573_),
    .A1(_03623_),
    .S(net240),
    .X(_03624_));
 sky130_fd_sc_hd__mux2_1 _08623_ (.A0(_03527_),
    .A1(_03624_),
    .S(net216),
    .X(_03625_));
 sky130_fd_sc_hd__a22o_1 _08624_ (.A1(_03425_),
    .A2(net185),
    .B1(_03625_),
    .B2(net186),
    .X(_03626_));
 sky130_fd_sc_hd__o31a_1 _08625_ (.A1(net209),
    .A2(_03414_),
    .A3(_03415_),
    .B1(net573),
    .X(_03627_));
 sky130_fd_sc_hd__o21a_1 _08626_ (.A1(net210),
    .A2(_03431_),
    .B1(_03627_),
    .X(_03628_));
 sky130_fd_sc_hd__o21ai_1 _08627_ (.A1(_03626_),
    .A2(_03628_),
    .B1(net193),
    .Y(_03629_));
 sky130_fd_sc_hd__a21oi_1 _08628_ (.A1(net209),
    .A2(_03420_),
    .B1(_03581_),
    .Y(_03630_));
 sky130_fd_sc_hd__o22a_1 _08629_ (.A1(_03417_),
    .A2(_03530_),
    .B1(_03630_),
    .B2(_03221_),
    .X(_03631_));
 sky130_fd_sc_hd__or2_1 _08630_ (.A(net193),
    .B(_03631_),
    .X(_03632_));
 sky130_fd_sc_hd__nand2_1 _08631_ (.A(_03004_),
    .B(net265),
    .Y(_03633_));
 sky130_fd_sc_hd__o31a_1 _08632_ (.A1(_03005_),
    .A2(_03009_),
    .A3(_03170_),
    .B1(_03633_),
    .X(_03634_));
 sky130_fd_sc_hd__o2111a_1 _08633_ (.A1(_03012_),
    .A2(_03183_),
    .B1(_03629_),
    .C1(_03632_),
    .D1(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__o211ai_2 _08634_ (.A1(_03621_),
    .A2(_03622_),
    .B1(_03635_),
    .C1(_03619_),
    .Y(_03636_));
 sky130_fd_sc_hd__and3_1 _08635_ (.A(net845),
    .B(net766),
    .C(net757),
    .X(_03637_));
 sky130_fd_sc_hd__a221o_1 _08636_ (.A1(net1296),
    .A2(net567),
    .B1(_03636_),
    .B2(net742),
    .C1(_03637_),
    .X(_00006_));
 sky130_fd_sc_hd__o21ai_1 _08637_ (.A1(_03005_),
    .A2(_03009_),
    .B1(_03616_),
    .Y(_03638_));
 sky130_fd_sc_hd__a21o_1 _08638_ (.A1(_03592_),
    .A2(_03615_),
    .B1(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__xnor2_1 _08639_ (.A(_02981_),
    .B(_03639_),
    .Y(_03640_));
 sky130_fd_sc_hd__a31o_1 _08640_ (.A1(_03011_),
    .A2(_03018_),
    .A3(_03023_),
    .B1(_03010_),
    .X(_03641_));
 sky130_fd_sc_hd__a21oi_1 _08641_ (.A1(_03595_),
    .A2(_03597_),
    .B1(_03027_),
    .Y(_03642_));
 sky130_fd_sc_hd__nor2_1 _08642_ (.A(_03641_),
    .B(_03642_),
    .Y(_03643_));
 sky130_fd_sc_hd__xnor2_1 _08643_ (.A(_02981_),
    .B(_03643_),
    .Y(_03644_));
 sky130_fd_sc_hd__mux2_1 _08644_ (.A0(_02973_),
    .A1(_03004_),
    .S(net190),
    .X(_03645_));
 sky130_fd_sc_hd__mux2_1 _08645_ (.A0(_03600_),
    .A1(_03645_),
    .S(net239),
    .X(_03646_));
 sky130_fd_sc_hd__mux2_1 _08646_ (.A0(_03558_),
    .A1(_03646_),
    .S(net219),
    .X(_03647_));
 sky130_fd_sc_hd__a22o_1 _08647_ (.A1(_03464_),
    .A2(net185),
    .B1(_03647_),
    .B2(net186),
    .X(_03648_));
 sky130_fd_sc_hd__mux2_1 _08648_ (.A0(_03450_),
    .A1(_03458_),
    .S(net206),
    .X(_03649_));
 sky130_fd_sc_hd__a21o_1 _08649_ (.A1(net573),
    .A2(_03649_),
    .B1(_03648_),
    .X(_03650_));
 sky130_fd_sc_hd__nor2_1 _08650_ (.A(net211),
    .B(_03455_),
    .Y(_03651_));
 sky130_fd_sc_hd__a22o_1 _08651_ (.A1(net198),
    .A2(net214),
    .B1(_03452_),
    .B2(_03651_),
    .X(_03652_));
 sky130_fd_sc_hd__o22a_1 _08652_ (.A1(_03452_),
    .A2(_03530_),
    .B1(_03652_),
    .B2(_03221_),
    .X(_03653_));
 sky130_fd_sc_hd__and2_1 _08653_ (.A(_02973_),
    .B(_02977_),
    .X(_03654_));
 sky130_fd_sc_hd__nand2_1 _08654_ (.A(net570),
    .B(_03654_),
    .Y(_03655_));
 sky130_fd_sc_hd__o221a_1 _08655_ (.A1(_02981_),
    .A2(_03183_),
    .B1(_03185_),
    .B2(_02972_),
    .C1(_03655_),
    .X(_03656_));
 sky130_fd_sc_hd__o21ai_1 _08656_ (.A1(net193),
    .A2(_03653_),
    .B1(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__a21o_1 _08657_ (.A1(net193),
    .A2(_03650_),
    .B1(_03657_),
    .X(_03658_));
 sky130_fd_sc_hd__a221o_1 _08658_ (.A1(net423),
    .A2(_03640_),
    .B1(_03644_),
    .B2(net428),
    .C1(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__and3_1 _08659_ (.A(net943),
    .B(net766),
    .C(net757),
    .X(_03660_));
 sky130_fd_sc_hd__a221o_1 _08660_ (.A1(net1294),
    .A2(net567),
    .B1(_03659_),
    .B2(net742),
    .C1(_03660_),
    .X(_00007_));
 sky130_fd_sc_hd__a21oi_1 _08661_ (.A1(_02982_),
    .A2(_03639_),
    .B1(_03654_),
    .Y(_03661_));
 sky130_fd_sc_hd__xnor2_1 _08662_ (.A(_02997_),
    .B(_03661_),
    .Y(_03662_));
 sky130_fd_sc_hd__o21bai_1 _08663_ (.A1(_02982_),
    .A2(_03643_),
    .B1_N(_02980_),
    .Y(_03663_));
 sky130_fd_sc_hd__xnor2_1 _08664_ (.A(_02997_),
    .B(_03663_),
    .Y(_03664_));
 sky130_fd_sc_hd__nand2_4 _08665_ (.A(net192),
    .B(net212),
    .Y(_03665_));
 sky130_fd_sc_hd__inv_2 _08666_ (.A(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__a21o_1 _08667_ (.A1(_03474_),
    .A2(_03475_),
    .B1(_03665_),
    .X(_03667_));
 sky130_fd_sc_hd__nor2_1 _08668_ (.A(_03477_),
    .B(_03530_),
    .Y(_03668_));
 sky130_fd_sc_hd__nor2_1 _08669_ (.A(net198),
    .B(_03221_),
    .Y(_03669_));
 sky130_fd_sc_hd__or2_1 _08670_ (.A(net198),
    .B(_03221_),
    .X(_03670_));
 sky130_fd_sc_hd__nor2_1 _08671_ (.A(_03202_),
    .B(_03669_),
    .Y(_03671_));
 sky130_fd_sc_hd__inv_2 _08672_ (.A(_03671_),
    .Y(_03672_));
 sky130_fd_sc_hd__o22a_1 _08673_ (.A1(_03173_),
    .A2(_03487_),
    .B1(_03668_),
    .B2(_03672_),
    .X(_03673_));
 sky130_fd_sc_hd__and2_1 _08674_ (.A(_03287_),
    .B(_03288_),
    .X(_03674_));
 sky130_fd_sc_hd__mux2_1 _08675_ (.A0(_03623_),
    .A1(_03674_),
    .S(net239),
    .X(_03675_));
 sky130_fd_sc_hd__mux2_1 _08676_ (.A0(_03574_),
    .A1(_03675_),
    .S(net220),
    .X(_03676_));
 sky130_fd_sc_hd__mux2_1 _08677_ (.A0(_03483_),
    .A1(_03676_),
    .S(net208),
    .X(_03677_));
 sky130_fd_sc_hd__a22o_1 _08678_ (.A1(_02994_),
    .A2(net570),
    .B1(net265),
    .B2(_02993_),
    .X(_03678_));
 sky130_fd_sc_hd__a22o_1 _08679_ (.A1(_02997_),
    .A2(_03512_),
    .B1(_03677_),
    .B2(_03176_),
    .X(_03679_));
 sky130_fd_sc_hd__a211o_1 _08680_ (.A1(_03667_),
    .A2(_03673_),
    .B1(_03678_),
    .C1(_03679_),
    .X(_03680_));
 sky130_fd_sc_hd__a221o_1 _08681_ (.A1(net423),
    .A2(_03662_),
    .B1(_03664_),
    .B2(net428),
    .C1(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__a22o_1 _08682_ (.A1(\brancher.pc_return[15] ),
    .A2(net569),
    .B1(_03681_),
    .B2(net741),
    .X(_03682_));
 sky130_fd_sc_hd__a31o_1 _08683_ (.A1(net1064),
    .A2(net766),
    .A3(net757),
    .B1(_03682_),
    .X(_00008_));
 sky130_fd_sc_hd__o21a_1 _08684_ (.A1(_02994_),
    .A2(_03654_),
    .B1(_02993_),
    .X(_03683_));
 sky130_fd_sc_hd__nand4_1 _08685_ (.A(_02982_),
    .B(_02997_),
    .C(_03591_),
    .D(_03615_),
    .Y(_03684_));
 sky130_fd_sc_hd__a211o_1 _08686_ (.A1(_03443_),
    .A2(_03494_),
    .B1(_03495_),
    .C1(_03684_),
    .X(_03685_));
 sky130_fd_sc_hd__a21o_1 _08687_ (.A1(_03590_),
    .A2(_03615_),
    .B1(_03638_),
    .X(_03686_));
 sky130_fd_sc_hd__a31oi_1 _08688_ (.A1(_02982_),
    .A2(_02997_),
    .A3(_03686_),
    .B1(_03683_),
    .Y(_03687_));
 sky130_fd_sc_hd__and2_1 _08689_ (.A(_03685_),
    .B(_03687_),
    .X(_03688_));
 sky130_fd_sc_hd__nand2_1 _08690_ (.A(net181),
    .B(_03688_),
    .Y(_03689_));
 sky130_fd_sc_hd__o21a_1 _08691_ (.A1(net181),
    .A2(_03688_),
    .B1(net423),
    .X(_03690_));
 sky130_fd_sc_hd__nor2_1 _08692_ (.A(_03028_),
    .B(_03597_),
    .Y(_03691_));
 sky130_fd_sc_hd__a221o_1 _08693_ (.A1(_02980_),
    .A2(_02995_),
    .B1(_02998_),
    .B2(_03641_),
    .C1(_02996_),
    .X(_03692_));
 sky130_fd_sc_hd__a211o_2 _08694_ (.A1(_03095_),
    .A2(_03501_),
    .B1(_03691_),
    .C1(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__xnor2_1 _08695_ (.A(net181),
    .B(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__o21ai_1 _08696_ (.A1(net195),
    .A2(_03165_),
    .B1(_03672_),
    .Y(_03695_));
 sky130_fd_sc_hd__nor2_2 _08697_ (.A(net193),
    .B(_03179_),
    .Y(_03696_));
 sky130_fd_sc_hd__nand3_1 _08698_ (.A(_02942_),
    .B(_02943_),
    .C(_02946_),
    .Y(_03697_));
 sky130_fd_sc_hd__o22a_1 _08699_ (.A1(_02941_),
    .A2(_03185_),
    .B1(_03697_),
    .B2(_03170_),
    .X(_03698_));
 sky130_fd_sc_hd__o21ai_1 _08700_ (.A1(net181),
    .A2(_03183_),
    .B1(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__a31o_1 _08701_ (.A1(_02700_),
    .A2(net221),
    .A3(_03696_),
    .B1(_03699_),
    .X(_03700_));
 sky130_fd_sc_hd__a31oi_1 _08702_ (.A1(net210),
    .A2(_03176_),
    .A3(_03506_),
    .B1(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__a21oi_1 _08703_ (.A1(net189),
    .A2(_02941_),
    .B1(_03190_),
    .Y(_03702_));
 sky130_fd_sc_hd__mux2_1 _08704_ (.A0(_03645_),
    .A1(_03702_),
    .S(net239),
    .X(_03703_));
 sky130_fd_sc_hd__or2_1 _08705_ (.A(net226),
    .B(_03703_),
    .X(_03704_));
 sky130_fd_sc_hd__o21ai_1 _08706_ (.A1(net219),
    .A2(_03601_),
    .B1(_03704_),
    .Y(_03705_));
 sky130_fd_sc_hd__o311a_1 _08707_ (.A1(net195),
    .A2(_03179_),
    .A3(_03705_),
    .B1(_03701_),
    .C1(_03695_),
    .X(_03706_));
 sky130_fd_sc_hd__o21ai_1 _08708_ (.A1(net426),
    .A2(_03694_),
    .B1(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__a21oi_1 _08709_ (.A1(_03689_),
    .A2(_03690_),
    .B1(_03707_),
    .Y(_03708_));
 sky130_fd_sc_hd__a2bb2o_1 _08710_ (.A1_N(net743),
    .A2_N(_03708_),
    .B1(net569),
    .B2(\brancher.pc_return[16] ),
    .X(_03709_));
 sky130_fd_sc_hd__a31o_1 _08711_ (.A1(net1030),
    .A2(net766),
    .A3(net757),
    .B1(_03709_),
    .X(_00009_));
 sky130_fd_sc_hd__nor3_1 _08712_ (.A(net181),
    .B(_02964_),
    .C(_03688_),
    .Y(_03710_));
 sky130_fd_sc_hd__nor2_1 _08713_ (.A(_02964_),
    .B(_03697_),
    .Y(_03711_));
 sky130_fd_sc_hd__o211a_1 _08714_ (.A1(net181),
    .A2(_03688_),
    .B1(_03697_),
    .C1(_02964_),
    .X(_03712_));
 sky130_fd_sc_hd__or4_1 _08715_ (.A(_03267_),
    .B(_03710_),
    .C(_03711_),
    .D(_03712_),
    .X(_03713_));
 sky130_fd_sc_hd__a211o_1 _08716_ (.A1(net181),
    .A2(_03693_),
    .B1(_02964_),
    .C1(_02948_),
    .X(_03714_));
 sky130_fd_sc_hd__nand3_1 _08717_ (.A(net181),
    .B(_02964_),
    .C(_03693_),
    .Y(_03715_));
 sky130_fd_sc_hd__and2_1 _08718_ (.A(_02948_),
    .B(_02964_),
    .X(_03716_));
 sky130_fd_sc_hd__inv_2 _08719_ (.A(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__and4_1 _08720_ (.A(net428),
    .B(_03714_),
    .C(_03715_),
    .D(_03717_),
    .X(_03718_));
 sky130_fd_sc_hd__nand2_1 _08721_ (.A(net198),
    .B(net197),
    .Y(_03719_));
 sky130_fd_sc_hd__nand2_2 _08722_ (.A(_03220_),
    .B(_03719_),
    .Y(_03720_));
 sky130_fd_sc_hd__and2_2 _08723_ (.A(_03220_),
    .B(_03719_),
    .X(_03721_));
 sky130_fd_sc_hd__nand2_1 _08724_ (.A(_03233_),
    .B(_03286_),
    .Y(_03722_));
 sky130_fd_sc_hd__nor2_1 _08725_ (.A(net245),
    .B(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__a21oi_1 _08726_ (.A1(net245),
    .A2(_03674_),
    .B1(_03723_),
    .Y(_03724_));
 sky130_fd_sc_hd__inv_2 _08727_ (.A(_03724_),
    .Y(_03725_));
 sky130_fd_sc_hd__mux2_2 _08728_ (.A0(_03624_),
    .A1(_03725_),
    .S(net219),
    .X(_03726_));
 sky130_fd_sc_hd__nor2_1 _08729_ (.A(net191),
    .B(_03670_),
    .Y(_03727_));
 sky130_fd_sc_hd__a221o_1 _08730_ (.A1(_02961_),
    .A2(net570),
    .B1(net265),
    .B2(_02962_),
    .C1(_03727_),
    .X(_03728_));
 sky130_fd_sc_hd__o21bai_1 _08731_ (.A1(_02964_),
    .A2(_03513_),
    .B1_N(_03728_),
    .Y(_03729_));
 sky130_fd_sc_hd__a32o_1 _08732_ (.A1(net221),
    .A2(_03271_),
    .A3(_03696_),
    .B1(_03726_),
    .B2(_03180_),
    .X(_03730_));
 sky130_fd_sc_hd__a21o_1 _08733_ (.A1(net185),
    .A2(_03528_),
    .B1(_03257_),
    .X(_03731_));
 sky130_fd_sc_hd__a221o_1 _08734_ (.A1(_03251_),
    .A2(_03721_),
    .B1(_03731_),
    .B2(net191),
    .C1(_03729_),
    .X(_03732_));
 sky130_fd_sc_hd__or2_1 _08735_ (.A(_03730_),
    .B(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__or3b_1 _08736_ (.A(_03733_),
    .B(_03718_),
    .C_N(_03713_),
    .X(_03734_));
 sky130_fd_sc_hd__and3_1 _08737_ (.A(net997),
    .B(net766),
    .C(net757),
    .X(_03735_));
 sky130_fd_sc_hd__a221o_1 _08738_ (.A1(net1295),
    .A2(net569),
    .B1(_03734_),
    .B2(net741),
    .C1(_03735_),
    .X(_00010_));
 sky130_fd_sc_hd__or2_1 _08739_ (.A(_02961_),
    .B(_03711_),
    .X(_03736_));
 sky130_fd_sc_hd__or3_1 _08740_ (.A(_02921_),
    .B(_03710_),
    .C(_03736_),
    .X(_03737_));
 sky130_fd_sc_hd__o21a_1 _08741_ (.A1(_03710_),
    .A2(_03736_),
    .B1(_02921_),
    .X(_03738_));
 sky130_fd_sc_hd__or3b_1 _08742_ (.A(_03738_),
    .B(_03267_),
    .C_N(_03737_),
    .X(_03739_));
 sky130_fd_sc_hd__nor2_1 _08743_ (.A(_02963_),
    .B(_03716_),
    .Y(_03740_));
 sky130_fd_sc_hd__and3_1 _08744_ (.A(_02921_),
    .B(_03715_),
    .C(_03740_),
    .X(_03741_));
 sky130_fd_sc_hd__a21oi_1 _08745_ (.A1(_03715_),
    .A2(_03740_),
    .B1(_02921_),
    .Y(_03742_));
 sky130_fd_sc_hd__or3_1 _08746_ (.A(net427),
    .B(_03741_),
    .C(_03742_),
    .X(_03743_));
 sky130_fd_sc_hd__a21o_1 _08747_ (.A1(net192),
    .A2(_03315_),
    .B1(_03720_),
    .X(_03744_));
 sky130_fd_sc_hd__and2_1 _08748_ (.A(_03159_),
    .B(_03161_),
    .X(_03745_));
 sky130_fd_sc_hd__mux2_1 _08749_ (.A0(_03702_),
    .A1(_03745_),
    .S(net241),
    .X(_03746_));
 sky130_fd_sc_hd__mux2_1 _08750_ (.A0(_03646_),
    .A1(_03746_),
    .S(net219),
    .X(_03747_));
 sky130_fd_sc_hd__a31o_1 _08751_ (.A1(net216),
    .A2(net186),
    .A3(_03326_),
    .B1(_03176_),
    .X(_03748_));
 sky130_fd_sc_hd__o221a_1 _08752_ (.A1(_03559_),
    .A2(_03665_),
    .B1(_03747_),
    .B2(_03173_),
    .C1(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__nand2_1 _08753_ (.A(net813),
    .B(_02919_),
    .Y(_03750_));
 sky130_fd_sc_hd__a32o_1 _08754_ (.A1(_02920_),
    .A2(net430),
    .A3(_03750_),
    .B1(net570),
    .B2(_02919_),
    .X(_03751_));
 sky130_fd_sc_hd__nor2_1 _08755_ (.A(_03749_),
    .B(_03751_),
    .Y(_03752_));
 sky130_fd_sc_hd__o211a_1 _08756_ (.A1(net196),
    .A2(_03313_),
    .B1(_03744_),
    .C1(_03752_),
    .X(_03753_));
 sky130_fd_sc_hd__and3_1 _08757_ (.A(_03739_),
    .B(_03743_),
    .C(_03753_),
    .X(_03754_));
 sky130_fd_sc_hd__a2bb2o_1 _08758_ (.A1_N(net743),
    .A2_N(_03754_),
    .B1(net569),
    .B2(\brancher.pc_return[18] ),
    .X(_03755_));
 sky130_fd_sc_hd__a31o_1 _08759_ (.A1(net990),
    .A2(net768),
    .A3(net757),
    .B1(_03755_),
    .X(_00011_));
 sky130_fd_sc_hd__or3_1 _08760_ (.A(_02919_),
    .B(_02935_),
    .C(_03738_),
    .X(_03756_));
 sky130_fd_sc_hd__o21ai_1 _08761_ (.A1(_02919_),
    .A2(_03738_),
    .B1(_02935_),
    .Y(_03757_));
 sky130_fd_sc_hd__and3_1 _08762_ (.A(net424),
    .B(_03756_),
    .C(_03757_),
    .X(_03758_));
 sky130_fd_sc_hd__and2_1 _08763_ (.A(_02914_),
    .B(_02918_),
    .X(_03759_));
 sky130_fd_sc_hd__nor2_1 _08764_ (.A(_03742_),
    .B(_03759_),
    .Y(_03760_));
 sky130_fd_sc_hd__or3b_1 _08765_ (.A(_03742_),
    .B(_03759_),
    .C_N(_02935_),
    .X(_03761_));
 sky130_fd_sc_hd__o211a_1 _08766_ (.A1(_02935_),
    .A2(_03760_),
    .B1(_03761_),
    .C1(net428),
    .X(_03762_));
 sky130_fd_sc_hd__nor2_1 _08767_ (.A(net241),
    .B(_03722_),
    .Y(_03763_));
 sky130_fd_sc_hd__and2_1 _08768_ (.A(_03230_),
    .B(_03232_),
    .X(_03764_));
 sky130_fd_sc_hd__a21o_1 _08769_ (.A1(net241),
    .A2(_03764_),
    .B1(_03763_),
    .X(_03765_));
 sky130_fd_sc_hd__mux2_1 _08770_ (.A0(_03675_),
    .A1(_03765_),
    .S(net225),
    .X(_03766_));
 sky130_fd_sc_hd__a221o_1 _08771_ (.A1(net185),
    .A2(_03575_),
    .B1(_03766_),
    .B2(net186),
    .C1(_03357_),
    .X(_03767_));
 sky130_fd_sc_hd__a21oi_1 _08772_ (.A1(net813),
    .A2(_02931_),
    .B1(_02932_),
    .Y(_03768_));
 sky130_fd_sc_hd__a221o_1 _08773_ (.A1(_02931_),
    .A2(_03169_),
    .B1(net431),
    .B2(_03768_),
    .C1(_03727_),
    .X(_03769_));
 sky130_fd_sc_hd__a31o_1 _08774_ (.A1(net222),
    .A2(_03363_),
    .A3(_03696_),
    .B1(_03769_),
    .X(_03770_));
 sky130_fd_sc_hd__a2bb2o_1 _08775_ (.A1_N(_03353_),
    .A2_N(_03720_),
    .B1(_03767_),
    .B2(net192),
    .X(_03771_));
 sky130_fd_sc_hd__or4_1 _08776_ (.A(_03758_),
    .B(_03762_),
    .C(_03770_),
    .D(_03771_),
    .X(_03772_));
 sky130_fd_sc_hd__and3_1 _08777_ (.A(net1069),
    .B(net768),
    .C(net757),
    .X(_03773_));
 sky130_fd_sc_hd__a221o_1 _08778_ (.A1(net1306),
    .A2(net569),
    .B1(_03772_),
    .B2(net741),
    .C1(_03773_),
    .X(_00012_));
 sky130_fd_sc_hd__nand2_1 _08779_ (.A(_02921_),
    .B(_02935_),
    .Y(_03774_));
 sky130_fd_sc_hd__inv_2 _08780_ (.A(_03774_),
    .Y(_03775_));
 sky130_fd_sc_hd__nor2_1 _08781_ (.A(_02919_),
    .B(_02931_),
    .Y(_03776_));
 sky130_fd_sc_hd__o2bb2a_1 _08782_ (.A1_N(_03736_),
    .A2_N(_03775_),
    .B1(_03776_),
    .B2(_02932_),
    .X(_03777_));
 sky130_fd_sc_hd__or3_1 _08783_ (.A(_02949_),
    .B(_02964_),
    .C(_03774_),
    .X(_03778_));
 sky130_fd_sc_hd__o21a_1 _08784_ (.A1(_03688_),
    .A2(_03778_),
    .B1(_03777_),
    .X(_03779_));
 sky130_fd_sc_hd__and2b_1 _08785_ (.A_N(_03779_),
    .B(_02892_),
    .X(_03780_));
 sky130_fd_sc_hd__xnor2_1 _08786_ (.A(_02892_),
    .B(_03779_),
    .Y(_03781_));
 sky130_fd_sc_hd__o21a_1 _08787_ (.A1(_02963_),
    .A2(_03716_),
    .B1(_02936_),
    .X(_03782_));
 sky130_fd_sc_hd__a211o_1 _08788_ (.A1(_02933_),
    .A2(_03759_),
    .B1(_03782_),
    .C1(_02934_),
    .X(_03783_));
 sky130_fd_sc_hd__a21oi_2 _08789_ (.A1(_02965_),
    .A2(_03693_),
    .B1(_03783_),
    .Y(_03784_));
 sky130_fd_sc_hd__nor2_1 _08790_ (.A(_02892_),
    .B(_03784_),
    .Y(_03785_));
 sky130_fd_sc_hd__a21o_1 _08791_ (.A1(_02892_),
    .A2(_03784_),
    .B1(net427),
    .X(_03786_));
 sky130_fd_sc_hd__a21boi_1 _08792_ (.A1(_02693_),
    .A2(_02926_),
    .B1_N(_03156_),
    .Y(_03787_));
 sky130_fd_sc_hd__mux2_1 _08793_ (.A0(_03745_),
    .A1(_03787_),
    .S(net241),
    .X(_03788_));
 sky130_fd_sc_hd__mux2_1 _08794_ (.A0(_03703_),
    .A1(_03788_),
    .S(net225),
    .X(_03789_));
 sky130_fd_sc_hd__a221o_1 _08795_ (.A1(net185),
    .A2(_03602_),
    .B1(_03789_),
    .B2(net186),
    .C1(_03390_),
    .X(_03790_));
 sky130_fd_sc_hd__a21oi_1 _08796_ (.A1(net191),
    .A2(_03392_),
    .B1(_03720_),
    .Y(_03791_));
 sky130_fd_sc_hd__nand2_1 _08797_ (.A(_02890_),
    .B(_03169_),
    .Y(_03792_));
 sky130_fd_sc_hd__o21a_1 _08798_ (.A1(_02885_),
    .A2(_02889_),
    .B1(net265),
    .X(_03793_));
 sky130_fd_sc_hd__a221o_1 _08799_ (.A1(_02892_),
    .A2(_03512_),
    .B1(_03696_),
    .B2(_03404_),
    .C1(_03793_),
    .X(_03794_));
 sky130_fd_sc_hd__a211oi_1 _08800_ (.A1(net191),
    .A2(_03790_),
    .B1(_03791_),
    .C1(_03794_),
    .Y(_03795_));
 sky130_fd_sc_hd__o211ai_1 _08801_ (.A1(_03785_),
    .A2(_03786_),
    .B1(_03792_),
    .C1(_03795_),
    .Y(_03796_));
 sky130_fd_sc_hd__a21o_1 _08802_ (.A1(net424),
    .A2(_03781_),
    .B1(_03796_),
    .X(_03797_));
 sky130_fd_sc_hd__and3_1 _08803_ (.A(net936),
    .B(net768),
    .C(net757),
    .X(_03798_));
 sky130_fd_sc_hd__a221o_1 _08804_ (.A1(net1341),
    .A2(net569),
    .B1(_03797_),
    .B2(net741),
    .C1(_03798_),
    .X(_00014_));
 sky130_fd_sc_hd__nand2_1 _08805_ (.A(_02890_),
    .B(_02904_),
    .Y(_03799_));
 sky130_fd_sc_hd__nand2_1 _08806_ (.A(_02892_),
    .B(_02904_),
    .Y(_03800_));
 sky130_fd_sc_hd__nor2_1 _08807_ (.A(_03779_),
    .B(_03800_),
    .Y(_03801_));
 sky130_fd_sc_hd__o211a_1 _08808_ (.A1(_03779_),
    .A2(_03800_),
    .B1(_03799_),
    .C1(net424),
    .X(_03802_));
 sky130_fd_sc_hd__o31a_1 _08809_ (.A1(_02890_),
    .A2(_02904_),
    .A3(_03780_),
    .B1(_03802_),
    .X(_03803_));
 sky130_fd_sc_hd__nand2_1 _08810_ (.A(_02891_),
    .B(_02905_),
    .Y(_03804_));
 sky130_fd_sc_hd__o311a_1 _08811_ (.A1(_02892_),
    .A2(_02904_),
    .A3(_03784_),
    .B1(_03804_),
    .C1(net428),
    .X(_03805_));
 sky130_fd_sc_hd__o31a_1 _08812_ (.A1(_02891_),
    .A2(_02905_),
    .A3(_03785_),
    .B1(_03805_),
    .X(_03806_));
 sky130_fd_sc_hd__nand2_1 _08813_ (.A(_03225_),
    .B(_03229_),
    .Y(_03807_));
 sky130_fd_sc_hd__nor2_1 _08814_ (.A(net249),
    .B(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__a21oi_1 _08815_ (.A1(net249),
    .A2(_03764_),
    .B1(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__mux2_1 _08816_ (.A0(_03724_),
    .A1(_03809_),
    .S(net219),
    .X(_03810_));
 sky130_fd_sc_hd__a2bb2o_1 _08817_ (.A1_N(_03179_),
    .A2_N(_03810_),
    .B1(net185),
    .B2(_03625_),
    .X(_03811_));
 sky130_fd_sc_hd__o21a_1 _08818_ (.A1(_03419_),
    .A2(_03811_),
    .B1(net192),
    .X(_03812_));
 sky130_fd_sc_hd__nand2_1 _08819_ (.A(_02898_),
    .B(_02902_),
    .Y(_03813_));
 sky130_fd_sc_hd__a2bb2o_1 _08820_ (.A1_N(_03170_),
    .A2_N(_03813_),
    .B1(net431),
    .B2(_02904_),
    .X(_03814_));
 sky130_fd_sc_hd__nor2_1 _08821_ (.A(_02897_),
    .B(_03185_),
    .Y(_03815_));
 sky130_fd_sc_hd__a2111o_1 _08822_ (.A1(_03421_),
    .A2(_03721_),
    .B1(_03727_),
    .C1(_03812_),
    .D1(_03815_),
    .X(_03816_));
 sky130_fd_sc_hd__a211o_1 _08823_ (.A1(_03425_),
    .A2(_03696_),
    .B1(_03814_),
    .C1(_03816_),
    .X(_03817_));
 sky130_fd_sc_hd__or3_1 _08824_ (.A(_03803_),
    .B(_03806_),
    .C(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__and3_1 _08825_ (.A(net900),
    .B(net767),
    .C(_03612_),
    .X(_03819_));
 sky130_fd_sc_hd__a221o_1 _08826_ (.A1(net1345),
    .A2(net568),
    .B1(_03818_),
    .B2(net741),
    .C1(_03819_),
    .X(_00015_));
 sky130_fd_sc_hd__nand2_1 _08827_ (.A(_03799_),
    .B(_03813_),
    .Y(_03820_));
 sky130_fd_sc_hd__or3_1 _08828_ (.A(_02862_),
    .B(_03801_),
    .C(_03820_),
    .X(_03821_));
 sky130_fd_sc_hd__o21a_1 _08829_ (.A1(_03801_),
    .A2(_03820_),
    .B1(_02862_),
    .X(_03822_));
 sky130_fd_sc_hd__and3b_1 _08830_ (.A_N(_03822_),
    .B(net424),
    .C(_03821_),
    .X(_03823_));
 sky130_fd_sc_hd__a21oi_1 _08831_ (.A1(_02891_),
    .A2(_02905_),
    .B1(_02903_),
    .Y(_03824_));
 sky130_fd_sc_hd__o31a_1 _08832_ (.A1(_02892_),
    .A2(_02904_),
    .A3(_03784_),
    .B1(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__o21ai_1 _08833_ (.A1(_02862_),
    .A2(_03825_),
    .B1(net428),
    .Y(_03826_));
 sky130_fd_sc_hd__a21oi_1 _08834_ (.A1(_02862_),
    .A2(_03825_),
    .B1(_03826_),
    .Y(_03827_));
 sky130_fd_sc_hd__o21a_1 _08835_ (.A1(_02854_),
    .A2(_02858_),
    .B1(net265),
    .X(_03828_));
 sky130_fd_sc_hd__a221o_1 _08836_ (.A1(_02859_),
    .A2(net572),
    .B1(_03512_),
    .B2(_02862_),
    .C1(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__a21o_1 _08837_ (.A1(net186),
    .A2(_03464_),
    .B1(_03176_),
    .X(_03830_));
 sky130_fd_sc_hd__and2_1 _08838_ (.A(_03152_),
    .B(_03155_),
    .X(_03831_));
 sky130_fd_sc_hd__mux2_1 _08839_ (.A0(_03787_),
    .A1(_03831_),
    .S(net241),
    .X(_03832_));
 sky130_fd_sc_hd__mux2_1 _08840_ (.A0(_03746_),
    .A1(_03832_),
    .S(net219),
    .X(_03833_));
 sky130_fd_sc_hd__o221a_1 _08841_ (.A1(_03647_),
    .A2(_03665_),
    .B1(_03833_),
    .B2(_03173_),
    .C1(_03830_),
    .X(_03834_));
 sky130_fd_sc_hd__a311o_1 _08842_ (.A1(net191),
    .A2(_03255_),
    .A3(_03454_),
    .B1(_03829_),
    .C1(_03834_),
    .X(_03835_));
 sky130_fd_sc_hd__o22a_1 _08843_ (.A1(net214),
    .A2(_03450_),
    .B1(_03453_),
    .B2(_03455_),
    .X(_03836_));
 sky130_fd_sc_hd__o21a_1 _08844_ (.A1(net196),
    .A2(_03836_),
    .B1(_03721_),
    .X(_03837_));
 sky130_fd_sc_hd__or4_1 _08845_ (.A(_03823_),
    .B(_03827_),
    .C(_03835_),
    .D(_03837_),
    .X(_03838_));
 sky130_fd_sc_hd__and3_1 _08846_ (.A(net864),
    .B(net767),
    .C(net757),
    .X(_03839_));
 sky130_fd_sc_hd__a221o_1 _08847_ (.A1(net1317),
    .A2(net568),
    .B1(_03838_),
    .B2(net741),
    .C1(_03839_),
    .X(_00016_));
 sky130_fd_sc_hd__or3_1 _08848_ (.A(_02859_),
    .B(_02878_),
    .C(_03822_),
    .X(_03840_));
 sky130_fd_sc_hd__o21ai_1 _08849_ (.A1(_02859_),
    .A2(_03822_),
    .B1(_02878_),
    .Y(_03841_));
 sky130_fd_sc_hd__and3_1 _08850_ (.A(net424),
    .B(_03840_),
    .C(_03841_),
    .X(_03842_));
 sky130_fd_sc_hd__o21ba_1 _08851_ (.A1(_02862_),
    .A2(_03825_),
    .B1_N(_02861_),
    .X(_03843_));
 sky130_fd_sc_hd__xor2_1 _08852_ (.A(_02878_),
    .B(_03843_),
    .X(_03844_));
 sky130_fd_sc_hd__o21a_1 _08853_ (.A1(net196),
    .A2(_03479_),
    .B1(_03721_),
    .X(_03845_));
 sky130_fd_sc_hd__nor2_1 _08854_ (.A(_02875_),
    .B(_03185_),
    .Y(_03846_));
 sky130_fd_sc_hd__a221o_1 _08855_ (.A1(_02874_),
    .A2(net572),
    .B1(_03512_),
    .B2(_02878_),
    .C1(_03846_),
    .X(_03847_));
 sky130_fd_sc_hd__a21o_1 _08856_ (.A1(_03483_),
    .A2(_03696_),
    .B1(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__nor2_1 _08857_ (.A(net241),
    .B(_03807_),
    .Y(_03849_));
 sky130_fd_sc_hd__and2_1 _08858_ (.A(_03223_),
    .B(_03224_),
    .X(_03850_));
 sky130_fd_sc_hd__a21o_1 _08859_ (.A1(net241),
    .A2(_03850_),
    .B1(_03849_),
    .X(_03851_));
 sky130_fd_sc_hd__mux2_1 _08860_ (.A0(_03765_),
    .A1(_03851_),
    .S(net225),
    .X(_03852_));
 sky130_fd_sc_hd__a221o_1 _08861_ (.A1(net185),
    .A2(_03676_),
    .B1(_03852_),
    .B2(net186),
    .C1(_03478_),
    .X(_03853_));
 sky130_fd_sc_hd__a211o_1 _08862_ (.A1(net191),
    .A2(_03853_),
    .B1(_03848_),
    .C1(_03845_),
    .X(_03854_));
 sky130_fd_sc_hd__a211o_1 _08863_ (.A1(net429),
    .A2(_03844_),
    .B1(_03854_),
    .C1(_03842_),
    .X(_03855_));
 sky130_fd_sc_hd__and3_1 _08864_ (.A(net855),
    .B(net767),
    .C(_03612_),
    .X(_03856_));
 sky130_fd_sc_hd__a221o_1 _08865_ (.A1(net1308),
    .A2(net568),
    .B1(_03855_),
    .B2(net741),
    .C1(_03856_),
    .X(_00017_));
 sky130_fd_sc_hd__a22oi_2 _08866_ (.A1(_02966_),
    .A2(_03693_),
    .B1(_03783_),
    .B2(net182),
    .Y(_03857_));
 sky130_fd_sc_hd__a21oi_1 _08867_ (.A1(_02861_),
    .A2(_02876_),
    .B1(_02877_),
    .Y(_03858_));
 sky130_fd_sc_hd__o21a_1 _08868_ (.A1(_02879_),
    .A2(_03824_),
    .B1(_03858_),
    .X(_03859_));
 sky130_fd_sc_hd__nand2_1 _08869_ (.A(_03857_),
    .B(_03859_),
    .Y(_03860_));
 sky130_fd_sc_hd__xnor2_1 _08870_ (.A(_02845_),
    .B(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__nand2_1 _08871_ (.A(_02862_),
    .B(_02878_),
    .Y(_03862_));
 sky130_fd_sc_hd__or3_1 _08872_ (.A(_03778_),
    .B(_03800_),
    .C(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__a21o_1 _08873_ (.A1(_03685_),
    .A2(_03687_),
    .B1(_03863_),
    .X(_03864_));
 sky130_fd_sc_hd__o21ba_1 _08874_ (.A1(_03777_),
    .A2(_03800_),
    .B1_N(_03820_),
    .X(_03865_));
 sky130_fd_sc_hd__nor2_1 _08875_ (.A(_02859_),
    .B(_02874_),
    .Y(_03866_));
 sky130_fd_sc_hd__o22a_1 _08876_ (.A1(_03862_),
    .A2(_03865_),
    .B1(_03866_),
    .B2(_02875_),
    .X(_03867_));
 sky130_fd_sc_hd__and2_1 _08877_ (.A(_03864_),
    .B(_03867_),
    .X(_03868_));
 sky130_fd_sc_hd__o21ai_1 _08878_ (.A1(_02845_),
    .A2(_03868_),
    .B1(net424),
    .Y(_03869_));
 sky130_fd_sc_hd__a21o_1 _08879_ (.A1(_02845_),
    .A2(_03868_),
    .B1(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__nand2_1 _08880_ (.A(_03147_),
    .B(_03153_),
    .Y(_03871_));
 sky130_fd_sc_hd__nor2_1 _08881_ (.A(net248),
    .B(_03871_),
    .Y(_03872_));
 sky130_fd_sc_hd__a21oi_1 _08882_ (.A1(net248),
    .A2(_03831_),
    .B1(_03872_),
    .Y(_03873_));
 sky130_fd_sc_hd__nand2_1 _08883_ (.A(_03174_),
    .B(_03873_),
    .Y(_03874_));
 sky130_fd_sc_hd__nor2_1 _08884_ (.A(net224),
    .B(_03173_),
    .Y(_03875_));
 sky130_fd_sc_hd__or2_1 _08885_ (.A(net225),
    .B(_03173_),
    .X(_03876_));
 sky130_fd_sc_hd__o2bb2a_1 _08886_ (.A1_N(_03666_),
    .A2_N(_03705_),
    .B1(_03788_),
    .B2(_03876_),
    .X(_03877_));
 sky130_fd_sc_hd__o211ai_2 _08887_ (.A1(_03176_),
    .A2(_03508_),
    .B1(_03874_),
    .C1(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__nand2_1 _08888_ (.A(_02843_),
    .B(net265),
    .Y(_03879_));
 sky130_fd_sc_hd__and2_1 _08889_ (.A(_03173_),
    .B(_03669_),
    .X(_03880_));
 sky130_fd_sc_hd__a21oi_1 _08890_ (.A1(net208),
    .A2(_03151_),
    .B1(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__o221a_1 _08891_ (.A1(_02845_),
    .A2(_03513_),
    .B1(_03671_),
    .B2(_03881_),
    .C1(_03879_),
    .X(_03882_));
 sky130_fd_sc_hd__o211a_1 _08892_ (.A1(_02842_),
    .A2(_03170_),
    .B1(_03878_),
    .C1(_03882_),
    .X(_03883_));
 sky130_fd_sc_hd__o211a_1 _08893_ (.A1(net427),
    .A2(_03861_),
    .B1(_03870_),
    .C1(_03883_),
    .X(_03884_));
 sky130_fd_sc_hd__a32o_1 _08894_ (.A1(net942),
    .A2(net767),
    .A3(_03612_),
    .B1(net568),
    .B2(\brancher.pc_return[24] ),
    .X(_03885_));
 sky130_fd_sc_hd__o21bai_2 _08895_ (.A1(net743),
    .A2(_03884_),
    .B1_N(_03885_),
    .Y(_00018_));
 sky130_fd_sc_hd__o211ai_1 _08896_ (.A1(_02845_),
    .A2(_03868_),
    .B1(_02830_),
    .C1(_02842_),
    .Y(_03886_));
 sky130_fd_sc_hd__nor2_1 _08897_ (.A(_02830_),
    .B(_02842_),
    .Y(_03887_));
 sky130_fd_sc_hd__a211o_1 _08898_ (.A1(_03864_),
    .A2(_03867_),
    .B1(_02830_),
    .C1(_02845_),
    .X(_03888_));
 sky130_fd_sc_hd__and4b_1 _08899_ (.A_N(_03887_),
    .B(net424),
    .C(_03886_),
    .D(_03888_),
    .X(_03889_));
 sky130_fd_sc_hd__nand2_1 _08900_ (.A(_02829_),
    .B(_02844_),
    .Y(_03890_));
 sky130_fd_sc_hd__a21o_1 _08901_ (.A1(_02845_),
    .A2(_03860_),
    .B1(_03890_),
    .X(_03891_));
 sky130_fd_sc_hd__a21bo_1 _08902_ (.A1(_03857_),
    .A2(_03859_),
    .B1_N(_02846_),
    .X(_03892_));
 sky130_fd_sc_hd__or2_1 _08903_ (.A(_02829_),
    .B(_02844_),
    .X(_03893_));
 sky130_fd_sc_hd__or2_1 _08904_ (.A(_03176_),
    .B(_03529_),
    .X(_03894_));
 sky130_fd_sc_hd__nand2_1 _08905_ (.A(_03222_),
    .B(_03240_),
    .Y(_03895_));
 sky130_fd_sc_hd__nor2_1 _08906_ (.A(net248),
    .B(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__a21oi_1 _08907_ (.A1(net249),
    .A2(_03850_),
    .B1(_03896_),
    .Y(_03897_));
 sky130_fd_sc_hd__a22oi_1 _08908_ (.A1(_03809_),
    .A2(_03875_),
    .B1(_03897_),
    .B2(_03174_),
    .Y(_03898_));
 sky130_fd_sc_hd__o211a_1 _08909_ (.A1(_03665_),
    .A2(_03726_),
    .B1(_03894_),
    .C1(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__and3_1 _08910_ (.A(net208),
    .B(_03250_),
    .C(_03721_),
    .X(_03900_));
 sky130_fd_sc_hd__a221o_1 _08911_ (.A1(_02827_),
    .A2(net572),
    .B1(net265),
    .B2(_02826_),
    .C1(_03880_),
    .X(_03901_));
 sky130_fd_sc_hd__a22o_1 _08912_ (.A1(_02829_),
    .A2(_03512_),
    .B1(_03532_),
    .B2(net191),
    .X(_03902_));
 sky130_fd_sc_hd__or4_1 _08913_ (.A(_03899_),
    .B(_03900_),
    .C(_03901_),
    .D(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__a41o_1 _08914_ (.A1(net429),
    .A2(_03891_),
    .A3(_03892_),
    .A4(_03893_),
    .B1(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__o21a_1 _08915_ (.A1(_03889_),
    .A2(_03904_),
    .B1(net741),
    .X(_03905_));
 sky130_fd_sc_hd__and2_2 _08916_ (.A(net767),
    .B(_03612_),
    .X(_03906_));
 sky130_fd_sc_hd__a221o_1 _08917_ (.A1(net1338),
    .A2(net568),
    .B1(_03906_),
    .B2(\brancher.imm13_b[5] ),
    .C1(_03905_),
    .X(_00019_));
 sky130_fd_sc_hd__and2b_1 _08918_ (.A_N(_02828_),
    .B(_03893_),
    .X(_03907_));
 sky130_fd_sc_hd__and3_1 _08919_ (.A(_02798_),
    .B(_03892_),
    .C(_03907_),
    .X(_03908_));
 sky130_fd_sc_hd__a21oi_1 _08920_ (.A1(_03892_),
    .A2(_03907_),
    .B1(_02798_),
    .Y(_03909_));
 sky130_fd_sc_hd__nor3_1 _08921_ (.A(net427),
    .B(_03908_),
    .C(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__nor2_1 _08922_ (.A(_02827_),
    .B(_03887_),
    .Y(_03911_));
 sky130_fd_sc_hd__and3b_1 _08923_ (.A_N(_02798_),
    .B(_03888_),
    .C(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__a21boi_1 _08924_ (.A1(_03888_),
    .A2(_03911_),
    .B1_N(_02798_),
    .Y(_03913_));
 sky130_fd_sc_hd__or3_1 _08925_ (.A(_03267_),
    .B(_03912_),
    .C(_03913_),
    .X(_03914_));
 sky130_fd_sc_hd__nand2_1 _08926_ (.A(_03145_),
    .B(_03148_),
    .Y(_03915_));
 sky130_fd_sc_hd__mux2_1 _08927_ (.A0(_03871_),
    .A1(_03915_),
    .S(net242),
    .X(_03916_));
 sky130_fd_sc_hd__nand2_1 _08928_ (.A(_03174_),
    .B(_03916_),
    .Y(_03917_));
 sky130_fd_sc_hd__o22a_1 _08929_ (.A1(_03665_),
    .A2(_03747_),
    .B1(_03832_),
    .B2(_03876_),
    .X(_03918_));
 sky130_fd_sc_hd__o211a_1 _08930_ (.A1(_03176_),
    .A2(_03560_),
    .B1(_03917_),
    .C1(_03918_),
    .X(_03919_));
 sky130_fd_sc_hd__o21a_1 _08931_ (.A1(_02790_),
    .A2(_02794_),
    .B1(net265),
    .X(_03920_));
 sky130_fd_sc_hd__a221o_1 _08932_ (.A1(_02797_),
    .A2(net572),
    .B1(_03512_),
    .B2(_02798_),
    .C1(_03920_),
    .X(_03921_));
 sky130_fd_sc_hd__o21bai_1 _08933_ (.A1(net196),
    .A2(_03553_),
    .B1_N(_03921_),
    .Y(_03922_));
 sky130_fd_sc_hd__a211o_1 _08934_ (.A1(_03551_),
    .A2(_03721_),
    .B1(_03919_),
    .C1(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__or4b_1 _08935_ (.A(_03880_),
    .B(_03910_),
    .C(_03923_),
    .D_N(_03914_),
    .X(_03924_));
 sky130_fd_sc_hd__a22o_1 _08936_ (.A1(net1453),
    .A2(net568),
    .B1(_03906_),
    .B2(\brancher.imm13_b[6] ),
    .X(_03925_));
 sky130_fd_sc_hd__a21o_1 _08937_ (.A1(net742),
    .A2(_03924_),
    .B1(_03925_),
    .X(_00020_));
 sky130_fd_sc_hd__o21bai_1 _08938_ (.A1(_02796_),
    .A2(_03909_),
    .B1_N(_02813_),
    .Y(_03926_));
 sky130_fd_sc_hd__or3b_1 _08939_ (.A(_02796_),
    .B(_03909_),
    .C_N(_02813_),
    .X(_03927_));
 sky130_fd_sc_hd__or3_1 _08940_ (.A(_02797_),
    .B(_02813_),
    .C(_03913_),
    .X(_03928_));
 sky130_fd_sc_hd__o21ai_1 _08941_ (.A1(_02797_),
    .A2(_03913_),
    .B1(_02813_),
    .Y(_03929_));
 sky130_fd_sc_hd__nor2_1 _08942_ (.A(_03665_),
    .B(_03766_),
    .Y(_03930_));
 sky130_fd_sc_hd__a21oi_1 _08943_ (.A1(_02693_),
    .A2(_02790_),
    .B1(_03238_),
    .Y(_03931_));
 sky130_fd_sc_hd__mux2_1 _08944_ (.A0(_03895_),
    .A1(_03931_),
    .S(net242),
    .X(_03932_));
 sky130_fd_sc_hd__inv_2 _08945_ (.A(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__a2bb2o_1 _08946_ (.A1_N(_03851_),
    .A2_N(_03876_),
    .B1(_03932_),
    .B2(_03174_),
    .X(_03934_));
 sky130_fd_sc_hd__a211o_1 _08947_ (.A1(_03177_),
    .A2(_03577_),
    .B1(_03930_),
    .C1(_03934_),
    .X(_03935_));
 sky130_fd_sc_hd__or3_1 _08948_ (.A(net211),
    .B(_03350_),
    .C(_03720_),
    .X(_03936_));
 sky130_fd_sc_hd__o211ai_1 _08949_ (.A1(net846),
    .A2(_02809_),
    .B1(_02810_),
    .C1(net431),
    .Y(_03937_));
 sky130_fd_sc_hd__nor2_1 _08950_ (.A(_03174_),
    .B(_03670_),
    .Y(_03938_));
 sky130_fd_sc_hd__o221a_1 _08951_ (.A1(_02809_),
    .A2(_03170_),
    .B1(_03174_),
    .B2(_03670_),
    .C1(_03937_),
    .X(_03939_));
 sky130_fd_sc_hd__o2111ai_2 _08952_ (.A1(net197),
    .A2(_03583_),
    .B1(_03935_),
    .C1(_03936_),
    .D1(_03939_),
    .Y(_03940_));
 sky130_fd_sc_hd__a31o_1 _08953_ (.A1(net424),
    .A2(_03928_),
    .A3(_03929_),
    .B1(_03940_),
    .X(_03941_));
 sky130_fd_sc_hd__a31o_1 _08954_ (.A1(net429),
    .A2(_03926_),
    .A3(_03927_),
    .B1(_03941_),
    .X(_03942_));
 sky130_fd_sc_hd__a22o_1 _08955_ (.A1(net1452),
    .A2(net568),
    .B1(_03906_),
    .B2(\brancher.imm13_b[7] ),
    .X(_03943_));
 sky130_fd_sc_hd__a21o_1 _08956_ (.A1(net741),
    .A2(_03942_),
    .B1(_03943_),
    .X(_00021_));
 sky130_fd_sc_hd__nand2_1 _08957_ (.A(_02798_),
    .B(_02813_),
    .Y(_03944_));
 sky130_fd_sc_hd__nand2_1 _08958_ (.A(_02797_),
    .B(_02810_),
    .Y(_03945_));
 sky130_fd_sc_hd__o211a_1 _08959_ (.A1(_03911_),
    .A2(_03944_),
    .B1(_03945_),
    .C1(_02809_),
    .X(_03946_));
 sky130_fd_sc_hd__o21ai_2 _08960_ (.A1(_03888_),
    .A2(_03944_),
    .B1(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__nand2_1 _08961_ (.A(_02768_),
    .B(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__o211a_1 _08962_ (.A1(_02768_),
    .A2(_03947_),
    .B1(_03948_),
    .C1(net424),
    .X(_03949_));
 sky130_fd_sc_hd__a21o_1 _08963_ (.A1(_03857_),
    .A2(_03859_),
    .B1(_02847_),
    .X(_03950_));
 sky130_fd_sc_hd__o21ai_1 _08964_ (.A1(_02796_),
    .A2(_02811_),
    .B1(_02812_),
    .Y(_03951_));
 sky130_fd_sc_hd__o31a_1 _08965_ (.A1(_02798_),
    .A2(_02813_),
    .A3(_03907_),
    .B1(_03951_),
    .X(_03952_));
 sky130_fd_sc_hd__nand2_1 _08966_ (.A(_03950_),
    .B(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__nand3_1 _08967_ (.A(_02768_),
    .B(_03950_),
    .C(_03952_),
    .Y(_03954_));
 sky130_fd_sc_hd__a21o_1 _08968_ (.A1(_03950_),
    .A2(_03952_),
    .B1(_02768_),
    .X(_03955_));
 sky130_fd_sc_hd__nor2_1 _08969_ (.A(net224),
    .B(_03873_),
    .Y(_03956_));
 sky130_fd_sc_hd__o21a_1 _08970_ (.A1(_02693_),
    .A2(_02761_),
    .B1(_03146_),
    .X(_03957_));
 sky130_fd_sc_hd__nand2_1 _08971_ (.A(net248),
    .B(_03915_),
    .Y(_03958_));
 sky130_fd_sc_hd__o211a_1 _08972_ (.A1(net248),
    .A2(_03957_),
    .B1(_03958_),
    .C1(net224),
    .X(_03959_));
 sky130_fd_sc_hd__or3_1 _08973_ (.A(_03173_),
    .B(_03956_),
    .C(_03959_),
    .X(_03960_));
 sky130_fd_sc_hd__o221a_1 _08974_ (.A1(_03176_),
    .A2(_03603_),
    .B1(_03665_),
    .B2(_03789_),
    .C1(_03960_),
    .X(_03961_));
 sky130_fd_sc_hd__and3_1 _08975_ (.A(_02761_),
    .B(_02762_),
    .C(_02765_),
    .X(_03962_));
 sky130_fd_sc_hd__nor2_1 _08976_ (.A(_02760_),
    .B(_03185_),
    .Y(_03963_));
 sky130_fd_sc_hd__a221o_1 _08977_ (.A1(_02768_),
    .A2(net431),
    .B1(_03962_),
    .B2(net572),
    .C1(_03938_),
    .X(_03964_));
 sky130_fd_sc_hd__a41o_1 _08978_ (.A1(net222),
    .A2(net209),
    .A3(_03144_),
    .A4(_03672_),
    .B1(_03961_),
    .X(_03965_));
 sky130_fd_sc_hd__or3_1 _08979_ (.A(_03963_),
    .B(_03964_),
    .C(_03965_),
    .X(_03966_));
 sky130_fd_sc_hd__a31o_1 _08980_ (.A1(net429),
    .A2(_03954_),
    .A3(_03955_),
    .B1(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__o21a_1 _08981_ (.A1(_03949_),
    .A2(_03967_),
    .B1(net742),
    .X(_03968_));
 sky130_fd_sc_hd__a221o_1 _08982_ (.A1(net1330),
    .A2(net568),
    .B1(_03906_),
    .B2(\brancher.imm13_b[8] ),
    .C1(_03968_),
    .X(_00022_));
 sky130_fd_sc_hd__a211o_1 _08983_ (.A1(_02768_),
    .A2(_03947_),
    .B1(_03962_),
    .C1(_02783_),
    .X(_03969_));
 sky130_fd_sc_hd__and2_1 _08984_ (.A(_02783_),
    .B(_03962_),
    .X(_03970_));
 sky130_fd_sc_hd__a31o_1 _08985_ (.A1(_02768_),
    .A2(_02783_),
    .A3(_03947_),
    .B1(_03970_),
    .X(_03971_));
 sky130_fd_sc_hd__and3b_1 _08986_ (.A_N(_03971_),
    .B(net425),
    .C(_03969_),
    .X(_03972_));
 sky130_fd_sc_hd__a21o_1 _08987_ (.A1(_02767_),
    .A2(_03955_),
    .B1(_02783_),
    .X(_03973_));
 sky130_fd_sc_hd__a31oi_1 _08988_ (.A1(_02767_),
    .A2(_02783_),
    .A3(_03955_),
    .B1(net427),
    .Y(_03974_));
 sky130_fd_sc_hd__and2b_1 _08989_ (.A_N(_03237_),
    .B(_03245_),
    .X(_03975_));
 sky130_fd_sc_hd__mux2_1 _08990_ (.A0(_03931_),
    .A1(_03975_),
    .S(net243),
    .X(_03976_));
 sky130_fd_sc_hd__a22o_1 _08991_ (.A1(_03875_),
    .A2(_03897_),
    .B1(_03976_),
    .B2(_03174_),
    .X(_03977_));
 sky130_fd_sc_hd__a2bb2o_1 _08992_ (.A1_N(_03176_),
    .A2_N(_03626_),
    .B1(_03666_),
    .B2(_03810_),
    .X(_03978_));
 sky130_fd_sc_hd__a21o_1 _08993_ (.A1(net192),
    .A2(_03630_),
    .B1(_03720_),
    .X(_03979_));
 sky130_fd_sc_hd__a22o_1 _08994_ (.A1(_02779_),
    .A2(net265),
    .B1(_03512_),
    .B2(_02783_),
    .X(_03980_));
 sky130_fd_sc_hd__a21oi_1 _08995_ (.A1(_02778_),
    .A2(net572),
    .B1(_03980_),
    .Y(_03981_));
 sky130_fd_sc_hd__o311a_1 _08996_ (.A1(net197),
    .A2(_03417_),
    .A3(_03530_),
    .B1(_03979_),
    .C1(_03981_),
    .X(_03982_));
 sky130_fd_sc_hd__o21ai_1 _08997_ (.A1(_03977_),
    .A2(_03978_),
    .B1(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__a211o_1 _08998_ (.A1(_03973_),
    .A2(_03974_),
    .B1(_03983_),
    .C1(_03972_),
    .X(_03984_));
 sky130_fd_sc_hd__a22o_1 _08999_ (.A1(\brancher.pc_return[29] ),
    .A2(net568),
    .B1(_03906_),
    .B2(\brancher.imm13_b[9] ),
    .X(_03985_));
 sky130_fd_sc_hd__a21o_1 _09000_ (.A1(net741),
    .A2(_03984_),
    .B1(_03985_),
    .X(_00023_));
 sky130_fd_sc_hd__or3_1 _09001_ (.A(_02752_),
    .B(_02778_),
    .C(_03971_),
    .X(_03986_));
 sky130_fd_sc_hd__o21a_1 _09002_ (.A1(_02778_),
    .A2(_03971_),
    .B1(_02752_),
    .X(_03987_));
 sky130_fd_sc_hd__nor2_1 _09003_ (.A(_03267_),
    .B(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__a21oi_1 _09004_ (.A1(_02782_),
    .A2(_03973_),
    .B1(_02752_),
    .Y(_03989_));
 sky130_fd_sc_hd__a311o_1 _09005_ (.A1(_02752_),
    .A2(_02782_),
    .A3(_03973_),
    .B1(_03989_),
    .C1(net427),
    .X(_03990_));
 sky130_fd_sc_hd__a21o_1 _09006_ (.A1(net191),
    .A2(_03652_),
    .B1(_03720_),
    .X(_03991_));
 sky130_fd_sc_hd__and2b_1 _09007_ (.A_N(_02746_),
    .B(_02750_),
    .X(_03992_));
 sky130_fd_sc_hd__a2bb2o_1 _09008_ (.A1_N(_02746_),
    .A2_N(_03185_),
    .B1(_03992_),
    .B2(net572),
    .X(_03993_));
 sky130_fd_sc_hd__a21oi_1 _09009_ (.A1(_02752_),
    .A2(net431),
    .B1(_03993_),
    .Y(_03994_));
 sky130_fd_sc_hd__o311a_1 _09010_ (.A1(net197),
    .A2(_03452_),
    .A3(_03530_),
    .B1(_03991_),
    .C1(_03994_),
    .X(_03995_));
 sky130_fd_sc_hd__nand2_1 _09011_ (.A(net247),
    .B(_03957_),
    .Y(_03996_));
 sky130_fd_sc_hd__or3_1 _09012_ (.A(net247),
    .B(_03140_),
    .C(_03142_),
    .X(_03997_));
 sky130_fd_sc_hd__a32o_1 _09013_ (.A1(_03174_),
    .A2(_03996_),
    .A3(_03997_),
    .B1(_03875_),
    .B2(_03916_),
    .X(_03998_));
 sky130_fd_sc_hd__o22ai_2 _09014_ (.A1(_03176_),
    .A2(_03648_),
    .B1(_03665_),
    .B2(_03833_),
    .Y(_03999_));
 sky130_fd_sc_hd__o2bb2a_1 _09015_ (.A1_N(_03986_),
    .A2_N(_03988_),
    .B1(_03998_),
    .B2(_03999_),
    .X(_04000_));
 sky130_fd_sc_hd__and3_1 _09016_ (.A(_03990_),
    .B(_03995_),
    .C(_04000_),
    .X(_04001_));
 sky130_fd_sc_hd__nor2_1 _09017_ (.A(net743),
    .B(_04001_),
    .Y(_04002_));
 sky130_fd_sc_hd__a221o_1 _09018_ (.A1(net1255),
    .A2(net569),
    .B1(_03906_),
    .B2(\brancher.imm13_b[10] ),
    .C1(_04002_),
    .X(_00025_));
 sky130_fd_sc_hd__o21ai_1 _09019_ (.A1(_03987_),
    .A2(_03992_),
    .B1(_02602_),
    .Y(_04003_));
 sky130_fd_sc_hd__o311a_1 _09020_ (.A1(_02602_),
    .A2(_03987_),
    .A3(_03992_),
    .B1(_04003_),
    .C1(net425),
    .X(_04004_));
 sky130_fd_sc_hd__o21ai_1 _09021_ (.A1(_02751_),
    .A2(_03989_),
    .B1(_02601_),
    .Y(_04005_));
 sky130_fd_sc_hd__o31a_1 _09022_ (.A1(_02601_),
    .A2(_02751_),
    .A3(_03989_),
    .B1(net429),
    .X(_04006_));
 sky130_fd_sc_hd__o21a_1 _09023_ (.A1(net247),
    .A2(_03244_),
    .B1(net223),
    .X(_04007_));
 sky130_fd_sc_hd__o21ai_1 _09024_ (.A1(net243),
    .A2(_03975_),
    .B1(_04007_),
    .Y(_04008_));
 sky130_fd_sc_hd__o221a_1 _09025_ (.A1(net223),
    .A2(_03933_),
    .B1(_04008_),
    .B2(_03354_),
    .C1(_03180_),
    .X(_04009_));
 sky130_fd_sc_hd__a221o_1 _09026_ (.A1(_02597_),
    .A2(net572),
    .B1(_03184_),
    .B2(_02596_),
    .C1(_03669_),
    .X(_04010_));
 sky130_fd_sc_hd__o32a_1 _09027_ (.A1(net197),
    .A2(_03477_),
    .A3(_03530_),
    .B1(_03513_),
    .B2(_02601_),
    .X(_04011_));
 sky130_fd_sc_hd__or3b_1 _09028_ (.A(_04009_),
    .B(_04010_),
    .C_N(_04011_),
    .X(_04012_));
 sky130_fd_sc_hd__a31o_1 _09029_ (.A1(_03172_),
    .A2(_03666_),
    .A3(_03852_),
    .B1(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__a31o_1 _09030_ (.A1(net196),
    .A2(_03172_),
    .A3(_03677_),
    .B1(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__a211oi_2 _09031_ (.A1(_04005_),
    .A2(_04006_),
    .B1(_04014_),
    .C1(_04004_),
    .Y(_04015_));
 sky130_fd_sc_hd__nor2_1 _09032_ (.A(net743),
    .B(_04015_),
    .Y(_04016_));
 sky130_fd_sc_hd__a221o_1 _09033_ (.A1(net1251),
    .A2(net568),
    .B1(_03906_),
    .B2(net842),
    .C1(_04016_),
    .X(_00026_));
 sky130_fd_sc_hd__and2_1 _09034_ (.A(net1133),
    .B(\dec.op_memSt ),
    .X(net168));
 sky130_fd_sc_hd__and2_1 _09035_ (.A(net1133),
    .B(\dec.op_memLd ),
    .X(net167));
 sky130_fd_sc_hd__nand2b_1 _09036_ (.A_N(_02597_),
    .B(_04003_),
    .Y(_04017_));
 sky130_fd_sc_hd__a31o_1 _09037_ (.A1(\alu.b_type ),
    .A2(net846),
    .A3(net943),
    .B1(_02601_),
    .X(_04018_));
 sky130_fd_sc_hd__a211oi_1 _09038_ (.A1(_02767_),
    .A2(_02782_),
    .B1(_02780_),
    .C1(_02754_),
    .Y(_04019_));
 sky130_fd_sc_hd__a31o_1 _09039_ (.A1(net183),
    .A2(_02784_),
    .A3(_03953_),
    .B1(_04019_),
    .X(_04020_));
 sky130_fd_sc_hd__a211oi_1 _09040_ (.A1(_02599_),
    .A2(_02751_),
    .B1(_04020_),
    .C1(_02600_),
    .Y(_04021_));
 sky130_fd_sc_hd__xnor2_1 _09041_ (.A(_04018_),
    .B(_04021_),
    .Y(_04022_));
 sky130_fd_sc_hd__a22oi_1 _09042_ (.A1(net425),
    .A2(_04017_),
    .B1(_04022_),
    .B2(net429),
    .Y(_04023_));
 sky130_fd_sc_hd__a22o_1 _09043_ (.A1(net425),
    .A2(_04017_),
    .B1(_04022_),
    .B2(net429),
    .X(_04024_));
 sky130_fd_sc_hd__a211o_1 _09044_ (.A1(net424),
    .A2(_03781_),
    .B1(_03796_),
    .C1(_03587_),
    .X(_04025_));
 sky130_fd_sc_hd__or4_1 _09045_ (.A(_03681_),
    .B(_03889_),
    .C(_03904_),
    .D(_04025_),
    .X(_04026_));
 sky130_fd_sc_hd__or4b_1 _09046_ (.A(_03302_),
    .B(_03341_),
    .C(_03381_),
    .D_N(_03410_),
    .X(_04027_));
 sky130_fd_sc_hd__or3_1 _09047_ (.A(_03520_),
    .B(_03611_),
    .C(_04027_),
    .X(_04028_));
 sky130_fd_sc_hd__or4_1 _09048_ (.A(_03134_),
    .B(_03215_),
    .C(_03437_),
    .D(_03468_),
    .X(_04029_));
 sky130_fd_sc_hd__or3_1 _09049_ (.A(_03492_),
    .B(_03542_),
    .C(_04029_),
    .X(_04030_));
 sky130_fd_sc_hd__or4_1 _09050_ (.A(_03659_),
    .B(_03734_),
    .C(_04028_),
    .D(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__or3b_1 _09051_ (.A(_03565_),
    .B(_03636_),
    .C_N(_03708_),
    .X(_04032_));
 sky130_fd_sc_hd__or4_1 _09052_ (.A(_03949_),
    .B(_03967_),
    .C(_04031_),
    .D(_04032_),
    .X(_04033_));
 sky130_fd_sc_hd__or4_1 _09053_ (.A(_03924_),
    .B(_03984_),
    .C(_04026_),
    .D(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__nand2_1 _09054_ (.A(_03754_),
    .B(_03884_),
    .Y(_04035_));
 sky130_fd_sc_hd__or4_1 _09055_ (.A(_03772_),
    .B(_03818_),
    .C(_03838_),
    .D(_04035_),
    .X(_04036_));
 sky130_fd_sc_hd__nor4_1 _09056_ (.A(_03855_),
    .B(_03942_),
    .C(_04034_),
    .D(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__nand2_1 _09057_ (.A(wRamByteEn),
    .B(_04024_),
    .Y(_04038_));
 sky130_fd_sc_hd__a41o_1 _09058_ (.A1(_04001_),
    .A2(_04015_),
    .A3(_04023_),
    .A4(net179),
    .B1(_01227_),
    .X(_04039_));
 sky130_fd_sc_hd__mux2_1 _09059_ (.A0(_04038_),
    .A1(_04039_),
    .S(_01218_),
    .X(_04040_));
 sky130_fd_sc_hd__a31o_1 _09060_ (.A1(_04001_),
    .A2(_04015_),
    .A3(net179),
    .B1(_04024_),
    .X(_04041_));
 sky130_fd_sc_hd__o2bb2a_1 _09061_ (.A1_N(net943),
    .A2_N(wRamWordEn),
    .B1(_03186_),
    .B2(_04024_),
    .X(_04042_));
 sky130_fd_sc_hd__nand2_1 _09062_ (.A(net943),
    .B(\brancher.funct3[0] ),
    .Y(_04043_));
 sky130_fd_sc_hd__mux2_1 _09063_ (.A0(_04043_),
    .A1(_04042_),
    .S(_04041_),
    .X(_04044_));
 sky130_fd_sc_hd__a21oi_4 _09064_ (.A1(_04040_),
    .A2(_04044_),
    .B1(_01209_),
    .Y(_04045_));
 sky130_fd_sc_hd__or2_1 _09065_ (.A(_03218_),
    .B(net176),
    .X(_04046_));
 sky130_fd_sc_hd__and2b_1 _09066_ (.A_N(\brancher.rJumping ),
    .B(net1137),
    .X(_04047_));
 sky130_fd_sc_hd__and3b_1 _09067_ (.A_N(net176),
    .B(_04047_),
    .C(_03217_),
    .X(_04048_));
 sky130_fd_sc_hd__and2_1 _09068_ (.A(net266),
    .B(net171),
    .X(_04049_));
 sky130_fd_sc_hd__and2b_1 _09069_ (.A_N(net964),
    .B(net1),
    .X(_04050_));
 sky130_fd_sc_hd__a22o_1 _09070_ (.A1(net961),
    .A2(\dec.rInstrustion[19] ),
    .B1(net753),
    .B2(net44),
    .X(_04051_));
 sky130_fd_sc_hd__a22o_1 _09071_ (.A1(net1070),
    .A2(net256),
    .B1(net169),
    .B2(_04051_),
    .X(_00034_));
 sky130_fd_sc_hd__a22o_1 _09072_ (.A1(net961),
    .A2(\dec.rInstrustion[15] ),
    .B1(net753),
    .B2(net40),
    .X(_04052_));
 sky130_fd_sc_hd__a22o_1 _09073_ (.A1(net1046),
    .A2(net257),
    .B1(net170),
    .B2(_04052_),
    .X(_00035_));
 sky130_fd_sc_hd__a22o_1 _09074_ (.A1(net961),
    .A2(\dec.rInstrustion[16] ),
    .B1(net753),
    .B2(net41),
    .X(_04053_));
 sky130_fd_sc_hd__a22o_1 _09075_ (.A1(net1012),
    .A2(net257),
    .B1(net170),
    .B2(_04053_),
    .X(_00036_));
 sky130_fd_sc_hd__a22o_1 _09076_ (.A1(net961),
    .A2(\dec.rInstrustion[17] ),
    .B1(net753),
    .B2(net42),
    .X(_04054_));
 sky130_fd_sc_hd__a22o_1 _09077_ (.A1(net994),
    .A2(net255),
    .B1(net169),
    .B2(_04054_),
    .X(_00037_));
 sky130_fd_sc_hd__a22o_1 _09078_ (.A1(net961),
    .A2(\dec.rInstrustion[18] ),
    .B1(net753),
    .B2(net43),
    .X(_04055_));
 sky130_fd_sc_hd__a22o_1 _09079_ (.A1(net986),
    .A2(net255),
    .B1(net169),
    .B2(_04055_),
    .X(_00038_));
 sky130_fd_sc_hd__a22o_1 _09080_ (.A1(net961),
    .A2(\dec.rInstrustion[2] ),
    .B1(net755),
    .B2(net56),
    .X(_04056_));
 sky130_fd_sc_hd__a22oi_1 _09081_ (.A1(net962),
    .A2(\dec.rInstrustion[1] ),
    .B1(net754),
    .B2(net45),
    .Y(_04057_));
 sky130_fd_sc_hd__a22oi_1 _09082_ (.A1(net962),
    .A2(\dec.rInstrustion[0] ),
    .B1(net754),
    .B2(net34),
    .Y(_04058_));
 sky130_fd_sc_hd__nor2_1 _09083_ (.A(_04057_),
    .B(_04058_),
    .Y(_04059_));
 sky130_fd_sc_hd__a22o_1 _09084_ (.A1(net962),
    .A2(\dec.rInstrustion[3] ),
    .B1(net754),
    .B2(net59),
    .X(_04060_));
 sky130_fd_sc_hd__inv_2 _09085_ (.A(_04060_),
    .Y(_04061_));
 sky130_fd_sc_hd__nor2_1 _09086_ (.A(_04056_),
    .B(_04060_),
    .Y(_04062_));
 sky130_fd_sc_hd__and3_1 _09087_ (.A(net171),
    .B(_04059_),
    .C(_04062_),
    .X(_04063_));
 sky130_fd_sc_hd__and2_1 _09088_ (.A(net266),
    .B(_04063_),
    .X(_04064_));
 sky130_fd_sc_hd__a22oi_2 _09089_ (.A1(net962),
    .A2(\dec.rInstrustion[6] ),
    .B1(net754),
    .B2(net62),
    .Y(_04065_));
 sky130_fd_sc_hd__a22o_1 _09090_ (.A1(net962),
    .A2(\dec.rInstrustion[6] ),
    .B1(net754),
    .B2(net62),
    .X(_04066_));
 sky130_fd_sc_hd__a22oi_1 _09091_ (.A1(net962),
    .A2(\dec.rInstrustion[4] ),
    .B1(net754),
    .B2(net60),
    .Y(_04067_));
 sky130_fd_sc_hd__a22o_1 _09092_ (.A1(net962),
    .A2(\dec.rInstrustion[4] ),
    .B1(net754),
    .B2(net60),
    .X(_04068_));
 sky130_fd_sc_hd__a22o_1 _09093_ (.A1(net963),
    .A2(\dec.rInstrustion[5] ),
    .B1(net754),
    .B2(net61),
    .X(_04069_));
 sky130_fd_sc_hd__and3_1 _09094_ (.A(net172),
    .B(_04068_),
    .C(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__a32o_1 _09095_ (.A1(_04064_),
    .A2(_04065_),
    .A3(_04070_),
    .B1(net257),
    .B2(\alu.r_type ),
    .X(_00039_));
 sky130_fd_sc_hd__o41a_1 _09096_ (.A1(\dec.op_memLd ),
    .A2(\dec.op_lui ),
    .A3(net740),
    .A4(_03218_),
    .B1(net1137),
    .X(_00040_));
 sky130_fd_sc_hd__a22o_1 _09097_ (.A1(net963),
    .A2(\dec.rInstrustion[12] ),
    .B1(net755),
    .B2(net37),
    .X(_04071_));
 sky130_fd_sc_hd__nand2_1 _09098_ (.A(net172),
    .B(_04071_),
    .Y(_04072_));
 sky130_fd_sc_hd__inv_2 _09099_ (.A(_04072_),
    .Y(_04073_));
 sky130_fd_sc_hd__a22o_1 _09100_ (.A1(net963),
    .A2(\dec.rInstrustion[13] ),
    .B1(net755),
    .B2(net38),
    .X(_04074_));
 sky130_fd_sc_hd__nor2_1 _09101_ (.A(_04072_),
    .B(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__or2_1 _09102_ (.A(_04066_),
    .B(_04069_),
    .X(_04076_));
 sky130_fd_sc_hd__nor2_1 _09103_ (.A(_04067_),
    .B(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__and4b_1 _09104_ (.A_N(net176),
    .B(_04047_),
    .C(_04077_),
    .D(_03217_),
    .X(_04078_));
 sky130_fd_sc_hd__and2_1 _09105_ (.A(net266),
    .B(_04078_),
    .X(_04079_));
 sky130_fd_sc_hd__nand2_1 _09106_ (.A(_04063_),
    .B(_04079_),
    .Y(_04080_));
 sky130_fd_sc_hd__a32o_1 _09107_ (.A1(_04063_),
    .A2(_04075_),
    .A3(_04079_),
    .B1(net259),
    .B2(net1447),
    .X(_00041_));
 sky130_fd_sc_hd__and3_1 _09108_ (.A(net172),
    .B(_04067_),
    .C(_04069_),
    .X(_04081_));
 sky130_fd_sc_hd__and3_2 _09109_ (.A(_04063_),
    .B(_04065_),
    .C(_04081_),
    .X(_04082_));
 sky130_fd_sc_hd__mux2_1 _09110_ (.A0(\dec.op_memSt ),
    .A1(_04082_),
    .S(net266),
    .X(_00042_));
 sky130_fd_sc_hd__a2bb2o_1 _09111_ (.A1_N(_04075_),
    .A2_N(_04080_),
    .B1(net1418),
    .B2(net259),
    .X(_00043_));
 sky130_fd_sc_hd__and2_1 _09112_ (.A(\dec.op_memLd ),
    .B(net257),
    .X(_04083_));
 sky130_fd_sc_hd__or2_1 _09113_ (.A(_04068_),
    .B(_04076_),
    .X(_04084_));
 sky130_fd_sc_hd__inv_2 _09114_ (.A(_04084_),
    .Y(_04085_));
 sky130_fd_sc_hd__a31o_1 _09115_ (.A1(net267),
    .A2(_04063_),
    .A3(_04085_),
    .B1(_04083_),
    .X(_00044_));
 sky130_fd_sc_hd__and4_1 _09116_ (.A(net172),
    .B(_04066_),
    .C(_04067_),
    .D(_04069_),
    .X(_04086_));
 sky130_fd_sc_hd__and4_1 _09117_ (.A(net171),
    .B(_04056_),
    .C(_04059_),
    .D(_04061_),
    .X(_04087_));
 sky130_fd_sc_hd__nor2_1 _09118_ (.A(_01208_),
    .B(net267),
    .Y(_04088_));
 sky130_fd_sc_hd__a31o_1 _09119_ (.A1(net267),
    .A2(_04086_),
    .A3(_04087_),
    .B1(_04088_),
    .X(_00045_));
 sky130_fd_sc_hd__and2_1 _09120_ (.A(_04056_),
    .B(_04060_),
    .X(_04089_));
 sky130_fd_sc_hd__and4_1 _09121_ (.A(net266),
    .B(net171),
    .C(_04059_),
    .D(_04089_),
    .X(_04090_));
 sky130_fd_sc_hd__a22o_1 _09122_ (.A1(net953),
    .A2(net258),
    .B1(_04086_),
    .B2(_04090_),
    .X(_00046_));
 sky130_fd_sc_hd__a22o_1 _09123_ (.A1(net951),
    .A2(net259),
    .B1(_04079_),
    .B2(_04087_),
    .X(_00047_));
 sky130_fd_sc_hd__and3_1 _09124_ (.A(net267),
    .B(_04065_),
    .C(_04070_),
    .X(_04091_));
 sky130_fd_sc_hd__a22o_1 _09125_ (.A1(net1339),
    .A2(net258),
    .B1(_04087_),
    .B2(_04091_),
    .X(_00048_));
 sky130_fd_sc_hd__a22o_1 _09126_ (.A1(net961),
    .A2(\dec.rInstrustion[20] ),
    .B1(net753),
    .B2(net46),
    .X(_04092_));
 sky130_fd_sc_hd__and3_1 _09127_ (.A(net266),
    .B(net171),
    .C(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__inv_2 _09128_ (.A(_04093_),
    .Y(_04094_));
 sky130_fd_sc_hd__a41o_1 _09129_ (.A1(net172),
    .A2(_04066_),
    .A3(_04068_),
    .A4(_04069_),
    .B1(_04078_),
    .X(_04095_));
 sky130_fd_sc_hd__and2_1 _09130_ (.A(_04063_),
    .B(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__and4_1 _09131_ (.A(net171),
    .B(_04059_),
    .C(_04085_),
    .D(_04089_),
    .X(_04097_));
 sky130_fd_sc_hd__a221o_1 _09132_ (.A1(_04063_),
    .A2(_04085_),
    .B1(_04086_),
    .B2(_04087_),
    .C1(_04097_),
    .X(_04098_));
 sky130_fd_sc_hd__nor2_2 _09133_ (.A(_04096_),
    .B(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__a22o_1 _09134_ (.A1(net964),
    .A2(\dec.rInstrustion[7] ),
    .B1(net753),
    .B2(net63),
    .X(_04100_));
 sky130_fd_sc_hd__a32o_1 _09135_ (.A1(net169),
    .A2(_04082_),
    .A3(_04100_),
    .B1(net256),
    .B2(\brancher.imm12_i_s[0] ),
    .X(_04101_));
 sky130_fd_sc_hd__o21bai_1 _09136_ (.A1(_04094_),
    .A2(_04099_),
    .B1_N(_04101_),
    .Y(_00049_));
 sky130_fd_sc_hd__a22o_1 _09137_ (.A1(\dec.rStall ),
    .A2(\dec.rInstrustion[21] ),
    .B1(net755),
    .B2(net47),
    .X(_04102_));
 sky130_fd_sc_hd__and3_1 _09138_ (.A(net266),
    .B(net171),
    .C(_04102_),
    .X(_04103_));
 sky130_fd_sc_hd__inv_2 _09139_ (.A(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__a22o_1 _09140_ (.A1(net961),
    .A2(\dec.rInstrustion[8] ),
    .B1(net753),
    .B2(net64),
    .X(_04105_));
 sky130_fd_sc_hd__a32o_1 _09141_ (.A1(net170),
    .A2(_04082_),
    .A3(_04105_),
    .B1(net256),
    .B2(\brancher.imm12_i_s[1] ),
    .X(_04106_));
 sky130_fd_sc_hd__o21bai_1 _09142_ (.A1(_04099_),
    .A2(_04104_),
    .B1_N(_04106_),
    .Y(_00050_));
 sky130_fd_sc_hd__a22o_1 _09143_ (.A1(net962),
    .A2(\dec.rInstrustion[22] ),
    .B1(net754),
    .B2(net48),
    .X(_04107_));
 sky130_fd_sc_hd__and3_1 _09144_ (.A(net266),
    .B(net171),
    .C(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__inv_2 _09145_ (.A(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__a22o_1 _09146_ (.A1(net962),
    .A2(\dec.rInstrustion[9] ),
    .B1(net755),
    .B2(net65),
    .X(_04110_));
 sky130_fd_sc_hd__a32o_1 _09147_ (.A1(net169),
    .A2(_04082_),
    .A3(_04110_),
    .B1(net257),
    .B2(\brancher.imm12_i_s[2] ),
    .X(_04111_));
 sky130_fd_sc_hd__o21bai_1 _09148_ (.A1(_04099_),
    .A2(_04109_),
    .B1_N(_04111_),
    .Y(_00051_));
 sky130_fd_sc_hd__a22o_1 _09149_ (.A1(net964),
    .A2(\dec.rInstrustion[23] ),
    .B1(net756),
    .B2(net49),
    .X(_04112_));
 sky130_fd_sc_hd__nand2_1 _09150_ (.A(net169),
    .B(_04112_),
    .Y(_04113_));
 sky130_fd_sc_hd__a22o_1 _09151_ (.A1(net964),
    .A2(\dec.rInstrustion[10] ),
    .B1(net756),
    .B2(net35),
    .X(_04114_));
 sky130_fd_sc_hd__and3_1 _09152_ (.A(_01251_),
    .B(net173),
    .C(_04114_),
    .X(_04115_));
 sky130_fd_sc_hd__a22oi_1 _09153_ (.A1(\brancher.imm12_i_s[3] ),
    .A2(net255),
    .B1(_04082_),
    .B2(_04115_),
    .Y(_04116_));
 sky130_fd_sc_hd__o21ai_1 _09154_ (.A1(_04099_),
    .A2(_04113_),
    .B1(_04116_),
    .Y(_00052_));
 sky130_fd_sc_hd__a22o_1 _09155_ (.A1(net961),
    .A2(\dec.rInstrustion[24] ),
    .B1(net753),
    .B2(net50),
    .X(_04117_));
 sky130_fd_sc_hd__and3_1 _09156_ (.A(net266),
    .B(net171),
    .C(_04117_),
    .X(_04118_));
 sky130_fd_sc_hd__inv_2 _09157_ (.A(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__a22o_1 _09158_ (.A1(net961),
    .A2(\dec.rInstrustion[11] ),
    .B1(net753),
    .B2(net36),
    .X(_04120_));
 sky130_fd_sc_hd__a32o_1 _09159_ (.A1(net169),
    .A2(_04082_),
    .A3(_04120_),
    .B1(net256),
    .B2(\brancher.imm12_i_s[4] ),
    .X(_04121_));
 sky130_fd_sc_hd__o21bai_1 _09160_ (.A1(_04099_),
    .A2(_04119_),
    .B1_N(_04121_),
    .Y(_00053_));
 sky130_fd_sc_hd__or3_4 _09161_ (.A(_04082_),
    .B(_04096_),
    .C(_04098_),
    .X(_04122_));
 sky130_fd_sc_hd__a22o_1 _09162_ (.A1(net964),
    .A2(\dec.rInstrustion[25] ),
    .B1(net756),
    .B2(net51),
    .X(_04123_));
 sky130_fd_sc_hd__and3_1 _09163_ (.A(net268),
    .B(net173),
    .C(_04123_),
    .X(_04124_));
 sky130_fd_sc_hd__a22o_1 _09164_ (.A1(\brancher.imm12_i_s[5] ),
    .A2(net250),
    .B1(_04122_),
    .B2(_04124_),
    .X(_00054_));
 sky130_fd_sc_hd__a22o_1 _09165_ (.A1(net964),
    .A2(\dec.rInstrustion[26] ),
    .B1(net756),
    .B2(net52),
    .X(_04125_));
 sky130_fd_sc_hd__and3_1 _09166_ (.A(net268),
    .B(net173),
    .C(_04125_),
    .X(_04126_));
 sky130_fd_sc_hd__a22o_1 _09167_ (.A1(\brancher.imm12_i_s[6] ),
    .A2(net250),
    .B1(_04122_),
    .B2(_04126_),
    .X(_00055_));
 sky130_fd_sc_hd__a22o_1 _09168_ (.A1(net964),
    .A2(\dec.rInstrustion[27] ),
    .B1(net756),
    .B2(net53),
    .X(_04127_));
 sky130_fd_sc_hd__and3_1 _09169_ (.A(net268),
    .B(net173),
    .C(_04127_),
    .X(_04128_));
 sky130_fd_sc_hd__a22o_1 _09170_ (.A1(\brancher.imm12_i_s[7] ),
    .A2(net250),
    .B1(_04122_),
    .B2(_04128_),
    .X(_00056_));
 sky130_fd_sc_hd__a22o_1 _09171_ (.A1(net964),
    .A2(\dec.rInstrustion[28] ),
    .B1(net756),
    .B2(net54),
    .X(_04129_));
 sky130_fd_sc_hd__and3_1 _09172_ (.A(net268),
    .B(net173),
    .C(_04129_),
    .X(_04130_));
 sky130_fd_sc_hd__a22o_1 _09173_ (.A1(\brancher.imm12_i_s[8] ),
    .A2(net250),
    .B1(_04122_),
    .B2(_04130_),
    .X(_00057_));
 sky130_fd_sc_hd__a22o_1 _09174_ (.A1(net964),
    .A2(\dec.rInstrustion[29] ),
    .B1(net756),
    .B2(net55),
    .X(_04131_));
 sky130_fd_sc_hd__and3_1 _09175_ (.A(net268),
    .B(net173),
    .C(_04131_),
    .X(_04132_));
 sky130_fd_sc_hd__a22o_1 _09176_ (.A1(\brancher.imm12_i_s[9] ),
    .A2(net251),
    .B1(_04122_),
    .B2(_04132_),
    .X(_00058_));
 sky130_fd_sc_hd__a22o_1 _09177_ (.A1(net962),
    .A2(\dec.rInstrustion[30] ),
    .B1(net754),
    .B2(net57),
    .X(_04133_));
 sky130_fd_sc_hd__and3_1 _09178_ (.A(net267),
    .B(net171),
    .C(_04133_),
    .X(_04134_));
 sky130_fd_sc_hd__a22o_1 _09179_ (.A1(\brancher.imm12_i_s[10] ),
    .A2(net259),
    .B1(_04122_),
    .B2(_04134_),
    .X(_00059_));
 sky130_fd_sc_hd__a22o_1 _09180_ (.A1(net964),
    .A2(\dec.rInstrustion[31] ),
    .B1(net756),
    .B2(net58),
    .X(_04135_));
 sky130_fd_sc_hd__and3_1 _09181_ (.A(net268),
    .B(net173),
    .C(_04135_),
    .X(_04136_));
 sky130_fd_sc_hd__a22o_1 _09182_ (.A1(net944),
    .A2(net252),
    .B1(_04122_),
    .B2(_04136_),
    .X(_00060_));
 sky130_fd_sc_hd__a22o_1 _09183_ (.A1(net1451),
    .A2(net963),
    .B1(net755),
    .B2(net39),
    .X(_04137_));
 sky130_fd_sc_hd__a22o_1 _09184_ (.A1(\brancher.funct3[2] ),
    .A2(net259),
    .B1(net170),
    .B2(_04137_),
    .X(_00061_));
 sky130_fd_sc_hd__a21o_1 _09185_ (.A1(net940),
    .A2(net256),
    .B1(_04118_),
    .X(_00062_));
 sky130_fd_sc_hd__a21o_1 _09186_ (.A1(net917),
    .A2(net256),
    .B1(_04093_),
    .X(_00063_));
 sky130_fd_sc_hd__a21o_1 _09187_ (.A1(net880),
    .A2(net257),
    .B1(_04103_),
    .X(_00064_));
 sky130_fd_sc_hd__a21o_1 _09188_ (.A1(net861),
    .A2(net257),
    .B1(_04108_),
    .X(_00065_));
 sky130_fd_sc_hd__o21ai_1 _09189_ (.A1(net790),
    .A2(_01251_),
    .B1(_04113_),
    .Y(_00066_));
 sky130_fd_sc_hd__mux2_1 _09190_ (.A0(\brancher.funct3[0] ),
    .A1(_04073_),
    .S(net267),
    .X(_00067_));
 sky130_fd_sc_hd__a22o_1 _09191_ (.A1(net846),
    .A2(net259),
    .B1(net170),
    .B2(_04074_),
    .X(_00068_));
 sky130_fd_sc_hd__a22o_1 _09192_ (.A1(\alu.b_type ),
    .A2(net257),
    .B1(_04064_),
    .B2(_04086_),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _09193_ (.A0(\brancher.pc_return[0] ),
    .A1(net1277),
    .S(net258),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _09194_ (.A0(\brancher.pc_return[1] ),
    .A1(net1284),
    .S(net255),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _09195_ (.A0(net1323),
    .A1(\brancher.rPc_current_reg2[2] ),
    .S(net255),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _09196_ (.A0(net1343),
    .A1(net1374),
    .S(net255),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _09197_ (.A0(net1324),
    .A1(\brancher.rPc_current_reg2[4] ),
    .S(net254),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _09198_ (.A0(net1326),
    .A1(\brancher.rPc_current_reg2[5] ),
    .S(net251),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _09199_ (.A0(net1309),
    .A1(\brancher.rPc_current_reg2[6] ),
    .S(net251),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _09200_ (.A0(\brancher.pc_return[7] ),
    .A1(net1281),
    .S(net251),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _09201_ (.A0(net1328),
    .A1(\brancher.rPc_current_reg2[8] ),
    .S(net251),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _09202_ (.A0(net1303),
    .A1(\brancher.rPc_current_reg2[9] ),
    .S(net252),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _09203_ (.A0(net1319),
    .A1(\brancher.rPc_current_reg2[10] ),
    .S(net252),
    .X(_00080_));
 sky130_fd_sc_hd__mux2_1 _09204_ (.A0(\brancher.pc_return[11] ),
    .A1(net1301),
    .S(net252),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _09205_ (.A0(net1311),
    .A1(\brancher.rPc_current_reg2[12] ),
    .S(net253),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _09206_ (.A0(net1296),
    .A1(\brancher.rPc_current_reg2[13] ),
    .S(net253),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _09207_ (.A0(net1294),
    .A1(\brancher.rPc_current_reg2[14] ),
    .S(net253),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _09208_ (.A0(net1299),
    .A1(\brancher.rPc_current_reg2[15] ),
    .S(net260),
    .X(_00085_));
 sky130_fd_sc_hd__mux2_1 _09209_ (.A0(net1300),
    .A1(\brancher.rPc_current_reg2[16] ),
    .S(net260),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _09210_ (.A0(net1295),
    .A1(\brancher.rPc_current_reg2[17] ),
    .S(net260),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _09211_ (.A0(net1313),
    .A1(\brancher.rPc_current_reg2[18] ),
    .S(net260),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _09212_ (.A0(net1306),
    .A1(\brancher.rPc_current_reg2[19] ),
    .S(net264),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _09213_ (.A0(net1341),
    .A1(\brancher.rPc_current_reg2[20] ),
    .S(net264),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _09214_ (.A0(\brancher.pc_return[21] ),
    .A1(net1334),
    .S(net261),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _09215_ (.A0(net1317),
    .A1(\brancher.rPc_current_reg2[22] ),
    .S(net261),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _09216_ (.A0(net1308),
    .A1(\brancher.rPc_current_reg2[23] ),
    .S(net261),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _09217_ (.A0(net1336),
    .A1(\brancher.rPc_current_reg2[24] ),
    .S(net262),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _09218_ (.A0(\brancher.pc_return[25] ),
    .A1(net1315),
    .S(net262),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_1 _09219_ (.A0(net1433),
    .A1(net1445),
    .S(net261),
    .X(_00096_));
 sky130_fd_sc_hd__mux2_1 _09220_ (.A0(net1344),
    .A1(\brancher.rPc_current_reg2[27] ),
    .S(net262),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _09221_ (.A0(net1330),
    .A1(\brancher.rPc_current_reg2[28] ),
    .S(net261),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _09222_ (.A0(net1332),
    .A1(\brancher.rPc_current_reg2[29] ),
    .S(net263),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _09223_ (.A0(net1255),
    .A1(net1305),
    .S(net263),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _09224_ (.A0(net1251),
    .A1(net1293),
    .S(net263),
    .X(_00101_));
 sky130_fd_sc_hd__nand3_1 _09225_ (.A(\rReg_d2[0] ),
    .B(net969),
    .C(net968),
    .Y(_04138_));
 sky130_fd_sc_hd__and4_1 _09226_ (.A(\rReg_d2[0] ),
    .B(net969),
    .C(net968),
    .D(net966),
    .X(_04139_));
 sky130_fd_sc_hd__and3_1 _09227_ (.A(\rReg_d2[4] ),
    .B(rRegWrEn2),
    .C(_04139_),
    .X(_04140_));
 sky130_fd_sc_hd__o21ai_1 _09228_ (.A1(net1446),
    .A2(net681),
    .B1(net1089),
    .Y(_04141_));
 sky130_fd_sc_hd__a21oi_1 _09229_ (.A1(_02685_),
    .A2(net681),
    .B1(_04141_),
    .Y(_00102_));
 sky130_fd_sc_hd__nand2_1 _09230_ (.A(net721),
    .B(net683),
    .Y(_04142_));
 sky130_fd_sc_hd__o211a_1 _09231_ (.A1(net1401),
    .A2(net683),
    .B1(_04142_),
    .C1(net1129),
    .X(_00103_));
 sky130_fd_sc_hd__nand2_1 _09232_ (.A(net713),
    .B(net680),
    .Y(_04143_));
 sky130_fd_sc_hd__o211a_1 _09233_ (.A1(net1393),
    .A2(net680),
    .B1(_04143_),
    .C1(net1108),
    .X(_00104_));
 sky130_fd_sc_hd__nand2_1 _09234_ (.A(net712),
    .B(net681),
    .Y(_04144_));
 sky130_fd_sc_hd__o211a_1 _09235_ (.A1(net1382),
    .A2(net681),
    .B1(_04144_),
    .C1(net1087),
    .X(_00105_));
 sky130_fd_sc_hd__nand2_1 _09236_ (.A(net723),
    .B(net683),
    .Y(_04145_));
 sky130_fd_sc_hd__o211a_1 _09237_ (.A1(net1388),
    .A2(net683),
    .B1(_04145_),
    .C1(net1126),
    .X(_00106_));
 sky130_fd_sc_hd__nand2_1 _09238_ (.A(net722),
    .B(net683),
    .Y(_04146_));
 sky130_fd_sc_hd__o211a_1 _09239_ (.A1(net1352),
    .A2(net683),
    .B1(_04146_),
    .C1(net1118),
    .X(_00107_));
 sky130_fd_sc_hd__nand2_1 _09240_ (.A(net725),
    .B(net681),
    .Y(_04147_));
 sky130_fd_sc_hd__o211a_1 _09241_ (.A1(net1419),
    .A2(net681),
    .B1(_04147_),
    .C1(net1071),
    .X(_00108_));
 sky130_fd_sc_hd__nand2_1 _09242_ (.A(net724),
    .B(net681),
    .Y(_04148_));
 sky130_fd_sc_hd__o211a_1 _09243_ (.A1(net1381),
    .A2(net681),
    .B1(_04148_),
    .C1(net1081),
    .X(_00109_));
 sky130_fd_sc_hd__nand2_1 _09244_ (.A(net689),
    .B(net683),
    .Y(_04149_));
 sky130_fd_sc_hd__o211a_1 _09245_ (.A1(net1367),
    .A2(net683),
    .B1(_04149_),
    .C1(net1121),
    .X(_00110_));
 sky130_fd_sc_hd__nand2_1 _09246_ (.A(net690),
    .B(net680),
    .Y(_04150_));
 sky130_fd_sc_hd__o211a_1 _09247_ (.A1(net1431),
    .A2(net680),
    .B1(_04150_),
    .C1(net1094),
    .X(_00111_));
 sky130_fd_sc_hd__nand2_1 _09248_ (.A(net692),
    .B(net681),
    .Y(_04151_));
 sky130_fd_sc_hd__o211a_1 _09249_ (.A1(net1407),
    .A2(net681),
    .B1(_04151_),
    .C1(net1075),
    .X(_00112_));
 sky130_fd_sc_hd__nand2_1 _09250_ (.A(net691),
    .B(net680),
    .Y(_04152_));
 sky130_fd_sc_hd__o211a_1 _09251_ (.A1(net1394),
    .A2(net680),
    .B1(_04152_),
    .C1(net1099),
    .X(_00113_));
 sky130_fd_sc_hd__nand2_1 _09252_ (.A(net693),
    .B(net680),
    .Y(_04153_));
 sky130_fd_sc_hd__o211a_1 _09253_ (.A1(net1411),
    .A2(net680),
    .B1(_04153_),
    .C1(net1103),
    .X(_00114_));
 sky130_fd_sc_hd__nand2_1 _09254_ (.A(net694),
    .B(net680),
    .Y(_04154_));
 sky130_fd_sc_hd__o211a_1 _09255_ (.A1(net1420),
    .A2(net680),
    .B1(_04154_),
    .C1(net1097),
    .X(_00115_));
 sky130_fd_sc_hd__nand2_1 _09256_ (.A(net696),
    .B(net682),
    .Y(_04155_));
 sky130_fd_sc_hd__o211a_1 _09257_ (.A1(net1378),
    .A2(net682),
    .B1(_04155_),
    .C1(net1115),
    .X(_00116_));
 sky130_fd_sc_hd__nand2_1 _09258_ (.A(net695),
    .B(net685),
    .Y(_04156_));
 sky130_fd_sc_hd__o211a_1 _09259_ (.A1(net1440),
    .A2(net685),
    .B1(_04156_),
    .C1(net1153),
    .X(_00117_));
 sky130_fd_sc_hd__nand2_1 _09260_ (.A(_02938_),
    .B(net686),
    .Y(_04157_));
 sky130_fd_sc_hd__o211a_1 _09261_ (.A1(net1415),
    .A2(net686),
    .B1(_04157_),
    .C1(net1202),
    .X(_00118_));
 sky130_fd_sc_hd__nand2_1 _09262_ (.A(net697),
    .B(net685),
    .Y(_04158_));
 sky130_fd_sc_hd__o211a_1 _09263_ (.A1(net1412),
    .A2(net685),
    .B1(_04158_),
    .C1(net1140),
    .X(_00119_));
 sky130_fd_sc_hd__nand2_1 _09264_ (.A(net700),
    .B(net685),
    .Y(_04159_));
 sky130_fd_sc_hd__o211a_1 _09265_ (.A1(net1430),
    .A2(net685),
    .B1(_04159_),
    .C1(net1100),
    .X(_00120_));
 sky130_fd_sc_hd__nand2_1 _09266_ (.A(net699),
    .B(net684),
    .Y(_04160_));
 sky130_fd_sc_hd__o211a_1 _09267_ (.A1(net1441),
    .A2(net684),
    .B1(_04160_),
    .C1(net1149),
    .X(_00121_));
 sky130_fd_sc_hd__nand2_1 _09268_ (.A(net702),
    .B(net682),
    .Y(_04161_));
 sky130_fd_sc_hd__o211a_1 _09269_ (.A1(net1351),
    .A2(net682),
    .B1(_04161_),
    .C1(net1113),
    .X(_00122_));
 sky130_fd_sc_hd__nand2_1 _09270_ (.A(net701),
    .B(net687),
    .Y(_04162_));
 sky130_fd_sc_hd__o211a_1 _09271_ (.A1(net1434),
    .A2(net687),
    .B1(_04162_),
    .C1(net1207),
    .X(_00123_));
 sky130_fd_sc_hd__nand2_1 _09272_ (.A(net704),
    .B(net686),
    .Y(_04163_));
 sky130_fd_sc_hd__o211a_1 _09273_ (.A1(net1442),
    .A2(net686),
    .B1(_04163_),
    .C1(net1195),
    .X(_00124_));
 sky130_fd_sc_hd__nand2_1 _09274_ (.A(net703),
    .B(net684),
    .Y(_04164_));
 sky130_fd_sc_hd__o211a_1 _09275_ (.A1(net1405),
    .A2(net684),
    .B1(_04164_),
    .C1(net1164),
    .X(_00125_));
 sky130_fd_sc_hd__nand2_1 _09276_ (.A(net705),
    .B(net685),
    .Y(_04165_));
 sky130_fd_sc_hd__o211a_1 _09277_ (.A1(net1402),
    .A2(net686),
    .B1(_04165_),
    .C1(net1182),
    .X(_00126_));
 sky130_fd_sc_hd__nand2_1 _09278_ (.A(net706),
    .B(net684),
    .Y(_04166_));
 sky130_fd_sc_hd__o211a_1 _09279_ (.A1(net1372),
    .A2(net684),
    .B1(_04166_),
    .C1(net1171),
    .X(_00127_));
 sky130_fd_sc_hd__nand2_1 _09280_ (.A(net708),
    .B(net685),
    .Y(_04167_));
 sky130_fd_sc_hd__o211a_1 _09281_ (.A1(net1413),
    .A2(net685),
    .B1(_04167_),
    .C1(net1158),
    .X(_00128_));
 sky130_fd_sc_hd__nand2_1 _09282_ (.A(_02800_),
    .B(net684),
    .Y(_04168_));
 sky130_fd_sc_hd__o211a_1 _09283_ (.A1(net1376),
    .A2(net684),
    .B1(_04168_),
    .C1(net1164),
    .X(_00129_));
 sky130_fd_sc_hd__nand2_1 _09284_ (.A(net710),
    .B(net684),
    .Y(_04169_));
 sky130_fd_sc_hd__o211a_1 _09285_ (.A1(net1371),
    .A2(net684),
    .B1(_04169_),
    .C1(net1170),
    .X(_00130_));
 sky130_fd_sc_hd__nand2_1 _09286_ (.A(net709),
    .B(net686),
    .Y(_04170_));
 sky130_fd_sc_hd__o211a_1 _09287_ (.A1(net1426),
    .A2(net686),
    .B1(_04170_),
    .C1(net1175),
    .X(_00131_));
 sky130_fd_sc_hd__nand2_1 _09288_ (.A(_02742_),
    .B(net686),
    .Y(_04171_));
 sky130_fd_sc_hd__o211a_1 _09289_ (.A1(net1365),
    .A2(net686),
    .B1(_04171_),
    .C1(net1192),
    .X(_00132_));
 sky130_fd_sc_hd__nand2_1 _09290_ (.A(net574),
    .B(net687),
    .Y(_04172_));
 sky130_fd_sc_hd__o211a_1 _09291_ (.A1(net1414),
    .A2(net687),
    .B1(_04172_),
    .C1(net1204),
    .X(_00133_));
 sky130_fd_sc_hd__xnor2_1 _09292_ (.A(\rReg_d2[4] ),
    .B(_04139_),
    .Y(_04173_));
 sky130_fd_sc_hd__and2b_2 _09293_ (.A_N(_04173_),
    .B(_01974_),
    .X(_04174_));
 sky130_fd_sc_hd__nand2b_4 _09294_ (.A_N(_04173_),
    .B(_01974_),
    .Y(_04175_));
 sky130_fd_sc_hd__and3_1 _09295_ (.A(_01213_),
    .B(net970),
    .C(\rReg_d2[2] ),
    .X(_04176_));
 sky130_fd_sc_hd__nand3_4 _09296_ (.A(net966),
    .B(net536),
    .C(net674),
    .Y(_04177_));
 sky130_fd_sc_hd__or2_2 _09297_ (.A(net965),
    .B(_04138_),
    .X(_04178_));
 sky130_fd_sc_hd__nand2_1 _09298_ (.A(net965),
    .B(_04138_),
    .Y(_04179_));
 sky130_fd_sc_hd__and2_2 _09299_ (.A(_04178_),
    .B(_04179_),
    .X(_04180_));
 sky130_fd_sc_hd__nor2_1 _09300_ (.A(_02685_),
    .B(net505),
    .Y(_04181_));
 sky130_fd_sc_hd__a32o_1 _09301_ (.A1(net515),
    .A2(net672),
    .A3(net418),
    .B1(net419),
    .B2(\reg_module.gprf[32] ),
    .X(_04182_));
 sky130_fd_sc_hd__and2_1 _09302_ (.A(net1089),
    .B(_04182_),
    .X(_00134_));
 sky130_fd_sc_hd__nor2_1 _09303_ (.A(_02673_),
    .B(net506),
    .Y(_04183_));
 sky130_fd_sc_hd__a32o_1 _09304_ (.A1(net533),
    .A2(net679),
    .A3(net417),
    .B1(net420),
    .B2(\reg_module.gprf[33] ),
    .X(_04184_));
 sky130_fd_sc_hd__and2_1 _09305_ (.A(net1129),
    .B(_04184_),
    .X(_00135_));
 sky130_fd_sc_hd__nor2_1 _09306_ (.A(net713),
    .B(net506),
    .Y(_04185_));
 sky130_fd_sc_hd__a32o_1 _09307_ (.A1(net524),
    .A2(net671),
    .A3(net416),
    .B1(net420),
    .B2(\reg_module.gprf[34] ),
    .X(_04186_));
 sky130_fd_sc_hd__and2_1 _09308_ (.A(net1108),
    .B(_04186_),
    .X(_00136_));
 sky130_fd_sc_hd__nor2_1 _09309_ (.A(net712),
    .B(net505),
    .Y(_04187_));
 sky130_fd_sc_hd__a32o_1 _09310_ (.A1(net511),
    .A2(net672),
    .A3(net415),
    .B1(net419),
    .B2(\reg_module.gprf[35] ),
    .X(_04188_));
 sky130_fd_sc_hd__and2_1 _09311_ (.A(net1077),
    .B(_04188_),
    .X(_00137_));
 sky130_fd_sc_hd__nor2_1 _09312_ (.A(net723),
    .B(net506),
    .Y(_04189_));
 sky130_fd_sc_hd__a32o_1 _09313_ (.A1(net535),
    .A2(net674),
    .A3(net414),
    .B1(net420),
    .B2(\reg_module.gprf[36] ),
    .X(_04190_));
 sky130_fd_sc_hd__and2_1 _09314_ (.A(net1126),
    .B(_04190_),
    .X(_00138_));
 sky130_fd_sc_hd__nor2_1 _09315_ (.A(net722),
    .B(net506),
    .Y(_04191_));
 sky130_fd_sc_hd__a32o_1 _09316_ (.A1(net529),
    .A2(net674),
    .A3(net413),
    .B1(net420),
    .B2(\reg_module.gprf[37] ),
    .X(_04192_));
 sky130_fd_sc_hd__and2_1 _09317_ (.A(net1118),
    .B(_04192_),
    .X(_00139_));
 sky130_fd_sc_hd__nor2_1 _09318_ (.A(net725),
    .B(net505),
    .Y(_04193_));
 sky130_fd_sc_hd__a32o_1 _09319_ (.A1(net509),
    .A2(net672),
    .A3(net412),
    .B1(net419),
    .B2(\reg_module.gprf[38] ),
    .X(_04194_));
 sky130_fd_sc_hd__and2_1 _09320_ (.A(net1071),
    .B(_04194_),
    .X(_00140_));
 sky130_fd_sc_hd__nor2_1 _09321_ (.A(net724),
    .B(net505),
    .Y(_04195_));
 sky130_fd_sc_hd__a32o_1 _09322_ (.A1(net513),
    .A2(net672),
    .A3(net411),
    .B1(net419),
    .B2(\reg_module.gprf[39] ),
    .X(_04196_));
 sky130_fd_sc_hd__and2_1 _09323_ (.A(net1081),
    .B(_04196_),
    .X(_00141_));
 sky130_fd_sc_hd__nor2_1 _09324_ (.A(net689),
    .B(net506),
    .Y(_04197_));
 sky130_fd_sc_hd__a32o_1 _09325_ (.A1(net530),
    .A2(net674),
    .A3(net410),
    .B1(net420),
    .B2(\reg_module.gprf[40] ),
    .X(_04198_));
 sky130_fd_sc_hd__and2_1 _09326_ (.A(net1121),
    .B(_04198_),
    .X(_00142_));
 sky130_fd_sc_hd__nor2_1 _09327_ (.A(net690),
    .B(net505),
    .Y(_04199_));
 sky130_fd_sc_hd__a32o_1 _09328_ (.A1(net518),
    .A2(net671),
    .A3(_04199_),
    .B1(net419),
    .B2(\reg_module.gprf[41] ),
    .X(_04200_));
 sky130_fd_sc_hd__and2_1 _09329_ (.A(net1094),
    .B(_04200_),
    .X(_00143_));
 sky130_fd_sc_hd__nor2_1 _09330_ (.A(net692),
    .B(net505),
    .Y(_04201_));
 sky130_fd_sc_hd__a32o_1 _09331_ (.A1(net512),
    .A2(net672),
    .A3(_04201_),
    .B1(net419),
    .B2(\reg_module.gprf[42] ),
    .X(_04202_));
 sky130_fd_sc_hd__and2_1 _09332_ (.A(net1077),
    .B(_04202_),
    .X(_00144_));
 sky130_fd_sc_hd__nor2_1 _09333_ (.A(_03044_),
    .B(net505),
    .Y(_04203_));
 sky130_fd_sc_hd__a32o_1 _09334_ (.A1(net520),
    .A2(net671),
    .A3(net407),
    .B1(net419),
    .B2(\reg_module.gprf[43] ),
    .X(_04204_));
 sky130_fd_sc_hd__and2_1 _09335_ (.A(net1099),
    .B(_04204_),
    .X(_00145_));
 sky130_fd_sc_hd__nor2_1 _09336_ (.A(net693),
    .B(net505),
    .Y(_04205_));
 sky130_fd_sc_hd__a32o_1 _09337_ (.A1(net521),
    .A2(net671),
    .A3(net406),
    .B1(net420),
    .B2(\reg_module.gprf[44] ),
    .X(_04206_));
 sky130_fd_sc_hd__and2_1 _09338_ (.A(net1102),
    .B(_04206_),
    .X(_00146_));
 sky130_fd_sc_hd__nor2_1 _09339_ (.A(net694),
    .B(net505),
    .Y(_04207_));
 sky130_fd_sc_hd__a32o_1 _09340_ (.A1(net523),
    .A2(net671),
    .A3(net405),
    .B1(net419),
    .B2(\reg_module.gprf[45] ),
    .X(_04208_));
 sky130_fd_sc_hd__and2_1 _09341_ (.A(net1097),
    .B(_04208_),
    .X(_00147_));
 sky130_fd_sc_hd__nor2_1 _09342_ (.A(net696),
    .B(net506),
    .Y(_04209_));
 sky130_fd_sc_hd__a32o_1 _09343_ (.A1(net527),
    .A2(net673),
    .A3(net404),
    .B1(net419),
    .B2(\reg_module.gprf[46] ),
    .X(_04210_));
 sky130_fd_sc_hd__and2_1 _09344_ (.A(net1115),
    .B(_04210_),
    .X(_00148_));
 sky130_fd_sc_hd__nor2_1 _09345_ (.A(net695),
    .B(net507),
    .Y(_04211_));
 sky130_fd_sc_hd__a32o_1 _09346_ (.A1(net543),
    .A2(net676),
    .A3(net403),
    .B1(net421),
    .B2(\reg_module.gprf[47] ),
    .X(_04212_));
 sky130_fd_sc_hd__and2_1 _09347_ (.A(net1152),
    .B(_04212_),
    .X(_00149_));
 sky130_fd_sc_hd__nor2_1 _09348_ (.A(net698),
    .B(net508),
    .Y(_04213_));
 sky130_fd_sc_hd__a32o_1 _09349_ (.A1(net559),
    .A2(net677),
    .A3(net402),
    .B1(net422),
    .B2(\reg_module.gprf[48] ),
    .X(_04214_));
 sky130_fd_sc_hd__and2_1 _09350_ (.A(net1202),
    .B(_04214_),
    .X(_00150_));
 sky130_fd_sc_hd__nor2_1 _09351_ (.A(net697),
    .B(net507),
    .Y(_04215_));
 sky130_fd_sc_hd__a32o_1 _09352_ (.A1(net538),
    .A2(net676),
    .A3(net401),
    .B1(net421),
    .B2(\reg_module.gprf[49] ),
    .X(_04216_));
 sky130_fd_sc_hd__and2_1 _09353_ (.A(net1140),
    .B(_04216_),
    .X(_00151_));
 sky130_fd_sc_hd__nor2_1 _09354_ (.A(_02909_),
    .B(net507),
    .Y(_04217_));
 sky130_fd_sc_hd__a32o_1 _09355_ (.A1(net520),
    .A2(net676),
    .A3(net400),
    .B1(net421),
    .B2(\reg_module.gprf[50] ),
    .X(_04218_));
 sky130_fd_sc_hd__and2_1 _09356_ (.A(net1100),
    .B(_04218_),
    .X(_00152_));
 sky130_fd_sc_hd__nor2_1 _09357_ (.A(net699),
    .B(net508),
    .Y(_04219_));
 sky130_fd_sc_hd__a32o_1 _09358_ (.A1(net541),
    .A2(net675),
    .A3(net399),
    .B1(net422),
    .B2(\reg_module.gprf[51] ),
    .X(_04220_));
 sky130_fd_sc_hd__and2_1 _09359_ (.A(net1149),
    .B(_04220_),
    .X(_00153_));
 sky130_fd_sc_hd__nor2_1 _09360_ (.A(net702),
    .B(net505),
    .Y(_04221_));
 sky130_fd_sc_hd__a32o_1 _09361_ (.A1(net526),
    .A2(net671),
    .A3(net398),
    .B1(net419),
    .B2(\reg_module.gprf[52] ),
    .X(_04222_));
 sky130_fd_sc_hd__and2_1 _09362_ (.A(net1108),
    .B(_04222_),
    .X(_00154_));
 sky130_fd_sc_hd__nor2_1 _09363_ (.A(net701),
    .B(net508),
    .Y(_04223_));
 sky130_fd_sc_hd__a32o_1 _09364_ (.A1(net561),
    .A2(net677),
    .A3(net397),
    .B1(net422),
    .B2(\reg_module.gprf[53] ),
    .X(_04224_));
 sky130_fd_sc_hd__and2_1 _09365_ (.A(net1204),
    .B(_04224_),
    .X(_00155_));
 sky130_fd_sc_hd__nor2_1 _09366_ (.A(net704),
    .B(net508),
    .Y(_04225_));
 sky130_fd_sc_hd__a32o_1 _09367_ (.A1(net557),
    .A2(net677),
    .A3(_04225_),
    .B1(net422),
    .B2(\reg_module.gprf[54] ),
    .X(_04226_));
 sky130_fd_sc_hd__and2_1 _09368_ (.A(net1195),
    .B(_04226_),
    .X(_00156_));
 sky130_fd_sc_hd__nor2_1 _09369_ (.A(net703),
    .B(net507),
    .Y(_04227_));
 sky130_fd_sc_hd__a32o_1 _09370_ (.A1(net547),
    .A2(net675),
    .A3(net395),
    .B1(net421),
    .B2(\reg_module.gprf[55] ),
    .X(_04228_));
 sky130_fd_sc_hd__and2_1 _09371_ (.A(net1166),
    .B(_04228_),
    .X(_00157_));
 sky130_fd_sc_hd__nor2_1 _09372_ (.A(net705),
    .B(net507),
    .Y(_04229_));
 sky130_fd_sc_hd__a32o_1 _09373_ (.A1(net554),
    .A2(net676),
    .A3(_04229_),
    .B1(net421),
    .B2(\reg_module.gprf[56] ),
    .X(_04230_));
 sky130_fd_sc_hd__and2_1 _09374_ (.A(net1182),
    .B(_04230_),
    .X(_00158_));
 sky130_fd_sc_hd__nor2_1 _09375_ (.A(net706),
    .B(net507),
    .Y(_04231_));
 sky130_fd_sc_hd__a32o_1 _09376_ (.A1(net550),
    .A2(net675),
    .A3(net393),
    .B1(net421),
    .B2(\reg_module.gprf[57] ),
    .X(_04232_));
 sky130_fd_sc_hd__and2_1 _09377_ (.A(net1171),
    .B(_04232_),
    .X(_00159_));
 sky130_fd_sc_hd__nor2_1 _09378_ (.A(net708),
    .B(net507),
    .Y(_04233_));
 sky130_fd_sc_hd__a32o_1 _09379_ (.A1(net545),
    .A2(net676),
    .A3(net392),
    .B1(net421),
    .B2(\reg_module.gprf[58] ),
    .X(_04234_));
 sky130_fd_sc_hd__and2_1 _09380_ (.A(net1158),
    .B(_04234_),
    .X(_00160_));
 sky130_fd_sc_hd__nor2_1 _09381_ (.A(net707),
    .B(net507),
    .Y(_04235_));
 sky130_fd_sc_hd__a32o_1 _09382_ (.A1(net547),
    .A2(net675),
    .A3(net391),
    .B1(net421),
    .B2(\reg_module.gprf[59] ),
    .X(_04236_));
 sky130_fd_sc_hd__and2_1 _09383_ (.A(net1146),
    .B(_04236_),
    .X(_00161_));
 sky130_fd_sc_hd__nor2_1 _09384_ (.A(net710),
    .B(net507),
    .Y(_04237_));
 sky130_fd_sc_hd__a32o_1 _09385_ (.A1(net549),
    .A2(net675),
    .A3(net390),
    .B1(net421),
    .B2(\reg_module.gprf[60] ),
    .X(_04238_));
 sky130_fd_sc_hd__and2_1 _09386_ (.A(net1170),
    .B(_04238_),
    .X(_00162_));
 sky130_fd_sc_hd__nor2_1 _09387_ (.A(net709),
    .B(net507),
    .Y(_04239_));
 sky130_fd_sc_hd__a32o_1 _09388_ (.A1(net551),
    .A2(net675),
    .A3(net389),
    .B1(net421),
    .B2(\reg_module.gprf[61] ),
    .X(_04240_));
 sky130_fd_sc_hd__and2_1 _09389_ (.A(net1159),
    .B(_04240_),
    .X(_00163_));
 sky130_fd_sc_hd__nor2_1 _09390_ (.A(net711),
    .B(net508),
    .Y(_04241_));
 sky130_fd_sc_hd__a32o_1 _09391_ (.A1(net558),
    .A2(net677),
    .A3(_04241_),
    .B1(net422),
    .B2(\reg_module.gprf[62] ),
    .X(_04242_));
 sky130_fd_sc_hd__and2_1 _09392_ (.A(net1192),
    .B(_04242_),
    .X(_00164_));
 sky130_fd_sc_hd__nor2_1 _09393_ (.A(net574),
    .B(net508),
    .Y(_04243_));
 sky130_fd_sc_hd__a32o_1 _09394_ (.A1(net560),
    .A2(net677),
    .A3(net387),
    .B1(net422),
    .B2(\reg_module.gprf[63] ),
    .X(_04244_));
 sky130_fd_sc_hd__and2_1 _09395_ (.A(net1204),
    .B(_04244_),
    .X(_00165_));
 sky130_fd_sc_hd__and3b_4 _09396_ (.A_N(net970),
    .B(net968),
    .C(\rReg_d2[0] ),
    .X(_04245_));
 sky130_fd_sc_hd__nand3_4 _09397_ (.A(net965),
    .B(net536),
    .C(net748),
    .Y(_04246_));
 sky130_fd_sc_hd__a32o_1 _09398_ (.A1(net515),
    .A2(net418),
    .A3(net745),
    .B1(net383),
    .B2(\reg_module.gprf[64] ),
    .X(_04247_));
 sky130_fd_sc_hd__and2_1 _09399_ (.A(net1089),
    .B(_04247_),
    .X(_00166_));
 sky130_fd_sc_hd__a32o_1 _09400_ (.A1(net534),
    .A2(net417),
    .A3(net748),
    .B1(net384),
    .B2(\reg_module.gprf[65] ),
    .X(_04248_));
 sky130_fd_sc_hd__and2_1 _09401_ (.A(net1130),
    .B(_04248_),
    .X(_00167_));
 sky130_fd_sc_hd__a32o_1 _09402_ (.A1(net524),
    .A2(net416),
    .A3(net746),
    .B1(net384),
    .B2(\reg_module.gprf[66] ),
    .X(_04249_));
 sky130_fd_sc_hd__and2_1 _09403_ (.A(net1108),
    .B(_04249_),
    .X(_00168_));
 sky130_fd_sc_hd__a32o_1 _09404_ (.A1(net512),
    .A2(net415),
    .A3(net745),
    .B1(net383),
    .B2(\reg_module.gprf[67] ),
    .X(_04250_));
 sky130_fd_sc_hd__and2_1 _09405_ (.A(net1077),
    .B(_04250_),
    .X(_00169_));
 sky130_fd_sc_hd__a32o_1 _09406_ (.A1(net535),
    .A2(net414),
    .A3(net748),
    .B1(net384),
    .B2(\reg_module.gprf[68] ),
    .X(_04251_));
 sky130_fd_sc_hd__and2_1 _09407_ (.A(net1126),
    .B(_04251_),
    .X(_00170_));
 sky130_fd_sc_hd__a32o_1 _09408_ (.A1(net529),
    .A2(net413),
    .A3(net745),
    .B1(net383),
    .B2(\reg_module.gprf[69] ),
    .X(_04252_));
 sky130_fd_sc_hd__and2_1 _09409_ (.A(net1084),
    .B(_04252_),
    .X(_00171_));
 sky130_fd_sc_hd__a32o_1 _09410_ (.A1(net509),
    .A2(net412),
    .A3(net745),
    .B1(net383),
    .B2(\reg_module.gprf[70] ),
    .X(_04253_));
 sky130_fd_sc_hd__and2_1 _09411_ (.A(net1071),
    .B(_04253_),
    .X(_00172_));
 sky130_fd_sc_hd__a32o_1 _09412_ (.A1(net513),
    .A2(net411),
    .A3(net747),
    .B1(net383),
    .B2(\reg_module.gprf[71] ),
    .X(_04254_));
 sky130_fd_sc_hd__and2_1 _09413_ (.A(net1084),
    .B(_04254_),
    .X(_00173_));
 sky130_fd_sc_hd__a32o_1 _09414_ (.A1(net530),
    .A2(net410),
    .A3(net748),
    .B1(net384),
    .B2(\reg_module.gprf[72] ),
    .X(_04255_));
 sky130_fd_sc_hd__and2_1 _09415_ (.A(net1118),
    .B(_04255_),
    .X(_00174_));
 sky130_fd_sc_hd__a32o_1 _09416_ (.A1(net518),
    .A2(net409),
    .A3(net746),
    .B1(net383),
    .B2(\reg_module.gprf[73] ),
    .X(_04256_));
 sky130_fd_sc_hd__and2_1 _09417_ (.A(net1095),
    .B(_04256_),
    .X(_00175_));
 sky130_fd_sc_hd__a32o_1 _09418_ (.A1(net511),
    .A2(net408),
    .A3(net745),
    .B1(net383),
    .B2(\reg_module.gprf[74] ),
    .X(_04257_));
 sky130_fd_sc_hd__and2_1 _09419_ (.A(net1074),
    .B(_04257_),
    .X(_00176_));
 sky130_fd_sc_hd__a32o_1 _09420_ (.A1(net522),
    .A2(_04203_),
    .A3(net746),
    .B1(net383),
    .B2(\reg_module.gprf[75] ),
    .X(_04258_));
 sky130_fd_sc_hd__and2_1 _09421_ (.A(net1099),
    .B(_04258_),
    .X(_00177_));
 sky130_fd_sc_hd__a32o_1 _09422_ (.A1(net521),
    .A2(net406),
    .A3(net746),
    .B1(net383),
    .B2(\reg_module.gprf[76] ),
    .X(_04259_));
 sky130_fd_sc_hd__and2_1 _09423_ (.A(net1103),
    .B(_04259_),
    .X(_00178_));
 sky130_fd_sc_hd__a32o_1 _09424_ (.A1(net519),
    .A2(net405),
    .A3(net746),
    .B1(net384),
    .B2(\reg_module.gprf[77] ),
    .X(_04260_));
 sky130_fd_sc_hd__and2_1 _09425_ (.A(net1097),
    .B(_04260_),
    .X(_00179_));
 sky130_fd_sc_hd__a32o_1 _09426_ (.A1(net527),
    .A2(_04209_),
    .A3(net746),
    .B1(net383),
    .B2(\reg_module.gprf[78] ),
    .X(_04261_));
 sky130_fd_sc_hd__and2_1 _09427_ (.A(net1115),
    .B(_04261_),
    .X(_00180_));
 sky130_fd_sc_hd__a32o_1 _09428_ (.A1(net543),
    .A2(net403),
    .A3(net750),
    .B1(net385),
    .B2(\reg_module.gprf[79] ),
    .X(_04262_));
 sky130_fd_sc_hd__and2_1 _09429_ (.A(net1152),
    .B(_04262_),
    .X(_00181_));
 sky130_fd_sc_hd__a32o_1 _09430_ (.A1(net563),
    .A2(net402),
    .A3(net751),
    .B1(net386),
    .B2(\reg_module.gprf[80] ),
    .X(_04263_));
 sky130_fd_sc_hd__and2_1 _09431_ (.A(net1201),
    .B(_04263_),
    .X(_00182_));
 sky130_fd_sc_hd__a32o_1 _09432_ (.A1(net538),
    .A2(net401),
    .A3(net750),
    .B1(net385),
    .B2(\reg_module.gprf[81] ),
    .X(_04264_));
 sky130_fd_sc_hd__and2_1 _09433_ (.A(net1140),
    .B(_04264_),
    .X(_00183_));
 sky130_fd_sc_hd__a32o_1 _09434_ (.A1(net520),
    .A2(net400),
    .A3(net750),
    .B1(net385),
    .B2(\reg_module.gprf[82] ),
    .X(_04265_));
 sky130_fd_sc_hd__and2_1 _09435_ (.A(net1100),
    .B(_04265_),
    .X(_00184_));
 sky130_fd_sc_hd__a32o_1 _09436_ (.A1(net541),
    .A2(net399),
    .A3(net749),
    .B1(net386),
    .B2(\reg_module.gprf[83] ),
    .X(_04266_));
 sky130_fd_sc_hd__and2_1 _09437_ (.A(net1149),
    .B(_04266_),
    .X(_00185_));
 sky130_fd_sc_hd__a32o_1 _09438_ (.A1(net526),
    .A2(net398),
    .A3(net747),
    .B1(net384),
    .B2(\reg_module.gprf[84] ),
    .X(_04267_));
 sky130_fd_sc_hd__and2_1 _09439_ (.A(net1108),
    .B(_04267_),
    .X(_00186_));
 sky130_fd_sc_hd__a32o_1 _09440_ (.A1(net561),
    .A2(_04223_),
    .A3(net751),
    .B1(net386),
    .B2(\reg_module.gprf[85] ),
    .X(_04268_));
 sky130_fd_sc_hd__and2_1 _09441_ (.A(net1207),
    .B(_04268_),
    .X(_00187_));
 sky130_fd_sc_hd__a32o_1 _09442_ (.A1(net557),
    .A2(net396),
    .A3(net751),
    .B1(net386),
    .B2(\reg_module.gprf[86] ),
    .X(_04269_));
 sky130_fd_sc_hd__and2_1 _09443_ (.A(net1195),
    .B(_04269_),
    .X(_00188_));
 sky130_fd_sc_hd__a32o_1 _09444_ (.A1(net547),
    .A2(net395),
    .A3(net749),
    .B1(net385),
    .B2(\reg_module.gprf[87] ),
    .X(_04270_));
 sky130_fd_sc_hd__and2_1 _09445_ (.A(net1166),
    .B(_04270_),
    .X(_00189_));
 sky130_fd_sc_hd__a32o_1 _09446_ (.A1(net554),
    .A2(net394),
    .A3(net750),
    .B1(net385),
    .B2(\reg_module.gprf[88] ),
    .X(_04271_));
 sky130_fd_sc_hd__and2_1 _09447_ (.A(net1182),
    .B(_04271_),
    .X(_00190_));
 sky130_fd_sc_hd__a32o_1 _09448_ (.A1(net550),
    .A2(net393),
    .A3(net749),
    .B1(net385),
    .B2(\reg_module.gprf[89] ),
    .X(_04272_));
 sky130_fd_sc_hd__and2_1 _09449_ (.A(net1171),
    .B(_04272_),
    .X(_00191_));
 sky130_fd_sc_hd__a32o_1 _09450_ (.A1(net545),
    .A2(net392),
    .A3(net750),
    .B1(net385),
    .B2(\reg_module.gprf[90] ),
    .X(_04273_));
 sky130_fd_sc_hd__and2_1 _09451_ (.A(net1158),
    .B(_04273_),
    .X(_00192_));
 sky130_fd_sc_hd__a32o_1 _09452_ (.A1(net548),
    .A2(net391),
    .A3(net749),
    .B1(net385),
    .B2(\reg_module.gprf[91] ),
    .X(_04274_));
 sky130_fd_sc_hd__and2_1 _09453_ (.A(net1167),
    .B(_04274_),
    .X(_00193_));
 sky130_fd_sc_hd__a32o_1 _09454_ (.A1(net549),
    .A2(net390),
    .A3(net749),
    .B1(net385),
    .B2(\reg_module.gprf[92] ),
    .X(_04275_));
 sky130_fd_sc_hd__and2_1 _09455_ (.A(net1170),
    .B(_04275_),
    .X(_00194_));
 sky130_fd_sc_hd__a32o_1 _09456_ (.A1(net551),
    .A2(net389),
    .A3(net749),
    .B1(net385),
    .B2(\reg_module.gprf[93] ),
    .X(_04276_));
 sky130_fd_sc_hd__and2_1 _09457_ (.A(net1159),
    .B(_04276_),
    .X(_00195_));
 sky130_fd_sc_hd__a32o_1 _09458_ (.A1(net558),
    .A2(net388),
    .A3(net751),
    .B1(net386),
    .B2(\reg_module.gprf[94] ),
    .X(_04277_));
 sky130_fd_sc_hd__and2_1 _09459_ (.A(net1192),
    .B(_04277_),
    .X(_00196_));
 sky130_fd_sc_hd__a32o_1 _09460_ (.A1(net560),
    .A2(net387),
    .A3(net751),
    .B1(net386),
    .B2(\reg_module.gprf[95] ),
    .X(_04278_));
 sky130_fd_sc_hd__and2_1 _09461_ (.A(net1204),
    .B(_04278_),
    .X(_00197_));
 sky130_fd_sc_hd__nor3_4 _09462_ (.A(\rReg_d2[0] ),
    .B(net969),
    .C(_01214_),
    .Y(_04279_));
 sky130_fd_sc_hd__nand3_4 _09463_ (.A(net965),
    .B(net536),
    .C(net666),
    .Y(_04280_));
 sky130_fd_sc_hd__a32o_1 _09464_ (.A1(net516),
    .A2(net418),
    .A3(net663),
    .B1(net379),
    .B2(\reg_module.gprf[96] ),
    .X(_04281_));
 sky130_fd_sc_hd__and2_1 _09465_ (.A(net1090),
    .B(_04281_),
    .X(_00198_));
 sky130_fd_sc_hd__a32o_1 _09466_ (.A1(net534),
    .A2(net417),
    .A3(net666),
    .B1(net380),
    .B2(\reg_module.gprf[97] ),
    .X(_04282_));
 sky130_fd_sc_hd__and2_1 _09467_ (.A(net1130),
    .B(_04282_),
    .X(_00199_));
 sky130_fd_sc_hd__a32o_1 _09468_ (.A1(net524),
    .A2(_04185_),
    .A3(net664),
    .B1(net380),
    .B2(\reg_module.gprf[98] ),
    .X(_04283_));
 sky130_fd_sc_hd__and2_1 _09469_ (.A(net1108),
    .B(_04283_),
    .X(_00200_));
 sky130_fd_sc_hd__a32o_1 _09470_ (.A1(net515),
    .A2(net415),
    .A3(net663),
    .B1(net379),
    .B2(\reg_module.gprf[99] ),
    .X(_04284_));
 sky130_fd_sc_hd__and2_1 _09471_ (.A(net1087),
    .B(_04284_),
    .X(_00201_));
 sky130_fd_sc_hd__a32o_1 _09472_ (.A1(net535),
    .A2(net414),
    .A3(net666),
    .B1(net380),
    .B2(\reg_module.gprf[100] ),
    .X(_04285_));
 sky130_fd_sc_hd__and2_1 _09473_ (.A(net1126),
    .B(_04285_),
    .X(_00202_));
 sky130_fd_sc_hd__a32o_1 _09474_ (.A1(net529),
    .A2(net413),
    .A3(net666),
    .B1(net380),
    .B2(\reg_module.gprf[101] ),
    .X(_04286_));
 sky130_fd_sc_hd__and2_1 _09475_ (.A(net1085),
    .B(_04286_),
    .X(_00203_));
 sky130_fd_sc_hd__a32o_1 _09476_ (.A1(net509),
    .A2(net412),
    .A3(net663),
    .B1(net379),
    .B2(\reg_module.gprf[102] ),
    .X(_04287_));
 sky130_fd_sc_hd__and2_1 _09477_ (.A(net1071),
    .B(_04287_),
    .X(_00204_));
 sky130_fd_sc_hd__a32o_1 _09478_ (.A1(net513),
    .A2(net411),
    .A3(net663),
    .B1(net379),
    .B2(\reg_module.gprf[103] ),
    .X(_04288_));
 sky130_fd_sc_hd__and2_1 _09479_ (.A(net1083),
    .B(_04288_),
    .X(_00205_));
 sky130_fd_sc_hd__a32o_1 _09480_ (.A1(net530),
    .A2(net410),
    .A3(net666),
    .B1(net380),
    .B2(\reg_module.gprf[104] ),
    .X(_04289_));
 sky130_fd_sc_hd__and2_1 _09481_ (.A(net1121),
    .B(_04289_),
    .X(_00206_));
 sky130_fd_sc_hd__a32o_1 _09482_ (.A1(net518),
    .A2(net409),
    .A3(net664),
    .B1(net379),
    .B2(\reg_module.gprf[105] ),
    .X(_04290_));
 sky130_fd_sc_hd__and2_1 _09483_ (.A(net1095),
    .B(_04290_),
    .X(_00207_));
 sky130_fd_sc_hd__a32o_1 _09484_ (.A1(net511),
    .A2(_04201_),
    .A3(net663),
    .B1(net379),
    .B2(\reg_module.gprf[106] ),
    .X(_04291_));
 sky130_fd_sc_hd__and2_1 _09485_ (.A(net1075),
    .B(_04291_),
    .X(_00208_));
 sky130_fd_sc_hd__a32o_1 _09486_ (.A1(net520),
    .A2(net407),
    .A3(net664),
    .B1(net379),
    .B2(\reg_module.gprf[107] ),
    .X(_04292_));
 sky130_fd_sc_hd__and2_1 _09487_ (.A(net1100),
    .B(_04292_),
    .X(_00209_));
 sky130_fd_sc_hd__a32o_1 _09488_ (.A1(net521),
    .A2(net406),
    .A3(net664),
    .B1(net379),
    .B2(\reg_module.gprf[108] ),
    .X(_04293_));
 sky130_fd_sc_hd__and2_1 _09489_ (.A(net1103),
    .B(_04293_),
    .X(_00210_));
 sky130_fd_sc_hd__a32o_1 _09490_ (.A1(net519),
    .A2(net405),
    .A3(net664),
    .B1(net379),
    .B2(\reg_module.gprf[109] ),
    .X(_04294_));
 sky130_fd_sc_hd__and2_1 _09491_ (.A(net1098),
    .B(_04294_),
    .X(_00211_));
 sky130_fd_sc_hd__a32o_1 _09492_ (.A1(net527),
    .A2(_04209_),
    .A3(net665),
    .B1(net379),
    .B2(\reg_module.gprf[110] ),
    .X(_04295_));
 sky130_fd_sc_hd__and2_1 _09493_ (.A(net1115),
    .B(_04295_),
    .X(_00212_));
 sky130_fd_sc_hd__a32o_1 _09494_ (.A1(net543),
    .A2(net403),
    .A3(net668),
    .B1(net381),
    .B2(\reg_module.gprf[111] ),
    .X(_04296_));
 sky130_fd_sc_hd__and2_1 _09495_ (.A(net1153),
    .B(_04296_),
    .X(_00213_));
 sky130_fd_sc_hd__a32o_1 _09496_ (.A1(net559),
    .A2(net402),
    .A3(net669),
    .B1(net382),
    .B2(\reg_module.gprf[112] ),
    .X(_04297_));
 sky130_fd_sc_hd__and2_1 _09497_ (.A(net1199),
    .B(_04297_),
    .X(_00214_));
 sky130_fd_sc_hd__a32o_1 _09498_ (.A1(net538),
    .A2(net401),
    .A3(net668),
    .B1(net381),
    .B2(\reg_module.gprf[113] ),
    .X(_04298_));
 sky130_fd_sc_hd__and2_1 _09499_ (.A(net1140),
    .B(_04298_),
    .X(_00215_));
 sky130_fd_sc_hd__a32o_1 _09500_ (.A1(net538),
    .A2(net400),
    .A3(net668),
    .B1(net381),
    .B2(\reg_module.gprf[114] ),
    .X(_04299_));
 sky130_fd_sc_hd__and2_1 _09501_ (.A(net1139),
    .B(_04299_),
    .X(_00216_));
 sky130_fd_sc_hd__a32o_1 _09502_ (.A1(net540),
    .A2(net399),
    .A3(net667),
    .B1(net381),
    .B2(\reg_module.gprf[115] ),
    .X(_04300_));
 sky130_fd_sc_hd__and2_1 _09503_ (.A(net1149),
    .B(_04300_),
    .X(_00217_));
 sky130_fd_sc_hd__a32o_1 _09504_ (.A1(net526),
    .A2(net398),
    .A3(net664),
    .B1(net380),
    .B2(\reg_module.gprf[116] ),
    .X(_04301_));
 sky130_fd_sc_hd__and2_1 _09505_ (.A(net1113),
    .B(_04301_),
    .X(_00218_));
 sky130_fd_sc_hd__a32o_1 _09506_ (.A1(net561),
    .A2(net397),
    .A3(net669),
    .B1(net382),
    .B2(\reg_module.gprf[117] ),
    .X(_04302_));
 sky130_fd_sc_hd__and2_1 _09507_ (.A(net1204),
    .B(_04302_),
    .X(_00219_));
 sky130_fd_sc_hd__a32o_1 _09508_ (.A1(net557),
    .A2(net396),
    .A3(net669),
    .B1(net382),
    .B2(\reg_module.gprf[118] ),
    .X(_04303_));
 sky130_fd_sc_hd__and2_1 _09509_ (.A(net1195),
    .B(_04303_),
    .X(_00220_));
 sky130_fd_sc_hd__a32o_1 _09510_ (.A1(net548),
    .A2(net395),
    .A3(net667),
    .B1(net381),
    .B2(\reg_module.gprf[119] ),
    .X(_04304_));
 sky130_fd_sc_hd__and2_1 _09511_ (.A(net1165),
    .B(_04304_),
    .X(_00221_));
 sky130_fd_sc_hd__a32o_1 _09512_ (.A1(net554),
    .A2(net394),
    .A3(net667),
    .B1(net381),
    .B2(\reg_module.gprf[120] ),
    .X(_04305_));
 sky130_fd_sc_hd__and2_1 _09513_ (.A(net1182),
    .B(_04305_),
    .X(_00222_));
 sky130_fd_sc_hd__a32o_1 _09514_ (.A1(net550),
    .A2(net393),
    .A3(net667),
    .B1(net381),
    .B2(\reg_module.gprf[121] ),
    .X(_04306_));
 sky130_fd_sc_hd__and2_1 _09515_ (.A(net1171),
    .B(_04306_),
    .X(_00223_));
 sky130_fd_sc_hd__a32o_1 _09516_ (.A1(net545),
    .A2(net392),
    .A3(net668),
    .B1(net381),
    .B2(\reg_module.gprf[122] ),
    .X(_04307_));
 sky130_fd_sc_hd__and2_1 _09517_ (.A(net1158),
    .B(_04307_),
    .X(_00224_));
 sky130_fd_sc_hd__a32o_1 _09518_ (.A1(net547),
    .A2(net391),
    .A3(net667),
    .B1(net381),
    .B2(\reg_module.gprf[123] ),
    .X(_04308_));
 sky130_fd_sc_hd__and2_1 _09519_ (.A(net1166),
    .B(_04308_),
    .X(_00225_));
 sky130_fd_sc_hd__a32o_1 _09520_ (.A1(net549),
    .A2(net390),
    .A3(net667),
    .B1(net381),
    .B2(\reg_module.gprf[124] ),
    .X(_04309_));
 sky130_fd_sc_hd__and2_1 _09521_ (.A(net1170),
    .B(_04309_),
    .X(_00226_));
 sky130_fd_sc_hd__a32o_1 _09522_ (.A1(net551),
    .A2(net389),
    .A3(net668),
    .B1(net382),
    .B2(\reg_module.gprf[125] ),
    .X(_04310_));
 sky130_fd_sc_hd__and2_1 _09523_ (.A(net1175),
    .B(_04310_),
    .X(_00227_));
 sky130_fd_sc_hd__a32o_1 _09524_ (.A1(net558),
    .A2(_04241_),
    .A3(net669),
    .B1(net382),
    .B2(\reg_module.gprf[126] ),
    .X(_04311_));
 sky130_fd_sc_hd__and2_1 _09525_ (.A(net1192),
    .B(_04311_),
    .X(_00228_));
 sky130_fd_sc_hd__a32o_1 _09526_ (.A1(net560),
    .A2(net387),
    .A3(net669),
    .B1(net382),
    .B2(\reg_module.gprf[127] ),
    .X(_04312_));
 sky130_fd_sc_hd__and2_1 _09527_ (.A(net1204),
    .B(_04312_),
    .X(_00229_));
 sky130_fd_sc_hd__and3_4 _09528_ (.A(\rReg_d2[0] ),
    .B(net969),
    .C(_01214_),
    .X(_04313_));
 sky130_fd_sc_hd__nand3_4 _09529_ (.A(net967),
    .B(net536),
    .C(net658),
    .Y(_04314_));
 sky130_fd_sc_hd__a32o_1 _09530_ (.A1(net515),
    .A2(net418),
    .A3(net657),
    .B1(net375),
    .B2(\reg_module.gprf[128] ),
    .X(_04315_));
 sky130_fd_sc_hd__and2_1 _09531_ (.A(net1089),
    .B(_04315_),
    .X(_00230_));
 sky130_fd_sc_hd__a32o_1 _09532_ (.A1(net534),
    .A2(net417),
    .A3(net658),
    .B1(net376),
    .B2(\reg_module.gprf[129] ),
    .X(_04316_));
 sky130_fd_sc_hd__and2_1 _09533_ (.A(net1126),
    .B(_04316_),
    .X(_00231_));
 sky130_fd_sc_hd__a32o_1 _09534_ (.A1(net524),
    .A2(net416),
    .A3(net656),
    .B1(net375),
    .B2(\reg_module.gprf[130] ),
    .X(_04317_));
 sky130_fd_sc_hd__and2_1 _09535_ (.A(net1106),
    .B(_04317_),
    .X(_00232_));
 sky130_fd_sc_hd__a32o_1 _09536_ (.A1(net512),
    .A2(net415),
    .A3(net655),
    .B1(net375),
    .B2(\reg_module.gprf[131] ),
    .X(_04318_));
 sky130_fd_sc_hd__and2_1 _09537_ (.A(net1077),
    .B(_04318_),
    .X(_00233_));
 sky130_fd_sc_hd__a32o_1 _09538_ (.A1(net535),
    .A2(net414),
    .A3(net658),
    .B1(net376),
    .B2(\reg_module.gprf[132] ),
    .X(_04319_));
 sky130_fd_sc_hd__and2_1 _09539_ (.A(net1126),
    .B(_04319_),
    .X(_00234_));
 sky130_fd_sc_hd__a32o_1 _09540_ (.A1(net529),
    .A2(net413),
    .A3(net658),
    .B1(net376),
    .B2(\reg_module.gprf[133] ),
    .X(_04320_));
 sky130_fd_sc_hd__and2_1 _09541_ (.A(net1118),
    .B(_04320_),
    .X(_00235_));
 sky130_fd_sc_hd__a32o_1 _09542_ (.A1(net509),
    .A2(net412),
    .A3(net655),
    .B1(net375),
    .B2(\reg_module.gprf[134] ),
    .X(_04321_));
 sky130_fd_sc_hd__and2_1 _09543_ (.A(net1072),
    .B(_04321_),
    .X(_00236_));
 sky130_fd_sc_hd__a32o_1 _09544_ (.A1(net513),
    .A2(net411),
    .A3(net655),
    .B1(net375),
    .B2(\reg_module.gprf[135] ),
    .X(_04322_));
 sky130_fd_sc_hd__and2_1 _09545_ (.A(net1083),
    .B(_04322_),
    .X(_00237_));
 sky130_fd_sc_hd__a32o_1 _09546_ (.A1(net530),
    .A2(net410),
    .A3(_04313_),
    .B1(net376),
    .B2(\reg_module.gprf[136] ),
    .X(_04323_));
 sky130_fd_sc_hd__and2_1 _09547_ (.A(net1121),
    .B(_04323_),
    .X(_00238_));
 sky130_fd_sc_hd__a32o_1 _09548_ (.A1(net519),
    .A2(net409),
    .A3(net656),
    .B1(net375),
    .B2(\reg_module.gprf[137] ),
    .X(_04324_));
 sky130_fd_sc_hd__and2_1 _09549_ (.A(net1097),
    .B(_04324_),
    .X(_00239_));
 sky130_fd_sc_hd__a32o_1 _09550_ (.A1(net510),
    .A2(net408),
    .A3(net655),
    .B1(net375),
    .B2(\reg_module.gprf[138] ),
    .X(_04325_));
 sky130_fd_sc_hd__and2_1 _09551_ (.A(net1073),
    .B(_04325_),
    .X(_00240_));
 sky130_fd_sc_hd__a32o_1 _09552_ (.A1(net521),
    .A2(net407),
    .A3(net656),
    .B1(net375),
    .B2(\reg_module.gprf[139] ),
    .X(_04326_));
 sky130_fd_sc_hd__and2_1 _09553_ (.A(net1102),
    .B(_04326_),
    .X(_00241_));
 sky130_fd_sc_hd__a32o_1 _09554_ (.A1(net521),
    .A2(net406),
    .A3(net656),
    .B1(net376),
    .B2(\reg_module.gprf[140] ),
    .X(_04327_));
 sky130_fd_sc_hd__and2_1 _09555_ (.A(net1102),
    .B(_04327_),
    .X(_00242_));
 sky130_fd_sc_hd__a32o_1 _09556_ (.A1(net519),
    .A2(_04207_),
    .A3(net656),
    .B1(net375),
    .B2(\reg_module.gprf[141] ),
    .X(_04328_));
 sky130_fd_sc_hd__and2_1 _09557_ (.A(net1098),
    .B(_04328_),
    .X(_00243_));
 sky130_fd_sc_hd__a32o_1 _09558_ (.A1(net525),
    .A2(net404),
    .A3(net656),
    .B1(net375),
    .B2(\reg_module.gprf[142] ),
    .X(_04329_));
 sky130_fd_sc_hd__and2_1 _09559_ (.A(net1110),
    .B(_04329_),
    .X(_00244_));
 sky130_fd_sc_hd__a32o_1 _09560_ (.A1(net544),
    .A2(net403),
    .A3(net661),
    .B1(net377),
    .B2(\reg_module.gprf[143] ),
    .X(_04330_));
 sky130_fd_sc_hd__and2_1 _09561_ (.A(net1155),
    .B(_04330_),
    .X(_00245_));
 sky130_fd_sc_hd__a32o_1 _09562_ (.A1(net559),
    .A2(net402),
    .A3(net662),
    .B1(net378),
    .B2(\reg_module.gprf[144] ),
    .X(_04331_));
 sky130_fd_sc_hd__and2_1 _09563_ (.A(net1200),
    .B(_04331_),
    .X(_00246_));
 sky130_fd_sc_hd__a32o_1 _09564_ (.A1(net539),
    .A2(net401),
    .A3(net659),
    .B1(net377),
    .B2(\reg_module.gprf[145] ),
    .X(_04332_));
 sky130_fd_sc_hd__and2_1 _09565_ (.A(net1142),
    .B(_04332_),
    .X(_00247_));
 sky130_fd_sc_hd__a32o_1 _09566_ (.A1(net542),
    .A2(net400),
    .A3(net659),
    .B1(net377),
    .B2(\reg_module.gprf[146] ),
    .X(_04333_));
 sky130_fd_sc_hd__and2_1 _09567_ (.A(net1143),
    .B(_04333_),
    .X(_00248_));
 sky130_fd_sc_hd__a32o_1 _09568_ (.A1(net541),
    .A2(net399),
    .A3(net659),
    .B1(net377),
    .B2(\reg_module.gprf[147] ),
    .X(_04334_));
 sky130_fd_sc_hd__and2_1 _09569_ (.A(net1148),
    .B(_04334_),
    .X(_00249_));
 sky130_fd_sc_hd__a32o_1 _09570_ (.A1(net526),
    .A2(net398),
    .A3(net657),
    .B1(net376),
    .B2(\reg_module.gprf[148] ),
    .X(_04335_));
 sky130_fd_sc_hd__and2_1 _09571_ (.A(net1109),
    .B(_04335_),
    .X(_00250_));
 sky130_fd_sc_hd__a32o_1 _09572_ (.A1(net561),
    .A2(net397),
    .A3(net662),
    .B1(net378),
    .B2(\reg_module.gprf[149] ),
    .X(_04336_));
 sky130_fd_sc_hd__and2_1 _09573_ (.A(net1204),
    .B(_04336_),
    .X(_00251_));
 sky130_fd_sc_hd__a32o_1 _09574_ (.A1(net557),
    .A2(_04225_),
    .A3(net662),
    .B1(net378),
    .B2(\reg_module.gprf[150] ),
    .X(_04337_));
 sky130_fd_sc_hd__and2_1 _09575_ (.A(net1192),
    .B(_04337_),
    .X(_00252_));
 sky130_fd_sc_hd__a32o_1 _09576_ (.A1(net548),
    .A2(net395),
    .A3(net660),
    .B1(net377),
    .B2(\reg_module.gprf[151] ),
    .X(_04338_));
 sky130_fd_sc_hd__and2_1 _09577_ (.A(net1167),
    .B(_04338_),
    .X(_00253_));
 sky130_fd_sc_hd__a32o_1 _09578_ (.A1(net552),
    .A2(net394),
    .A3(net660),
    .B1(net377),
    .B2(\reg_module.gprf[152] ),
    .X(_04339_));
 sky130_fd_sc_hd__and2_1 _09579_ (.A(net1181),
    .B(_04339_),
    .X(_00254_));
 sky130_fd_sc_hd__a32o_1 _09580_ (.A1(net552),
    .A2(net393),
    .A3(net660),
    .B1(net377),
    .B2(\reg_module.gprf[153] ),
    .X(_04340_));
 sky130_fd_sc_hd__and2_1 _09581_ (.A(net1181),
    .B(_04340_),
    .X(_00255_));
 sky130_fd_sc_hd__a32o_1 _09582_ (.A1(net545),
    .A2(net392),
    .A3(net659),
    .B1(net377),
    .B2(\reg_module.gprf[154] ),
    .X(_04341_));
 sky130_fd_sc_hd__and2_1 _09583_ (.A(net1161),
    .B(_04341_),
    .X(_00256_));
 sky130_fd_sc_hd__a32o_1 _09584_ (.A1(net540),
    .A2(net391),
    .A3(net659),
    .B1(net377),
    .B2(\reg_module.gprf[155] ),
    .X(_04342_));
 sky130_fd_sc_hd__and2_1 _09585_ (.A(net1145),
    .B(_04342_),
    .X(_00257_));
 sky130_fd_sc_hd__a32o_1 _09586_ (.A1(net550),
    .A2(_04237_),
    .A3(net660),
    .B1(net377),
    .B2(\reg_module.gprf[156] ),
    .X(_04343_));
 sky130_fd_sc_hd__and2_1 _09587_ (.A(net1171),
    .B(_04343_),
    .X(_00258_));
 sky130_fd_sc_hd__a32o_1 _09588_ (.A1(net551),
    .A2(net389),
    .A3(net660),
    .B1(net378),
    .B2(\reg_module.gprf[157] ),
    .X(_04344_));
 sky130_fd_sc_hd__and2_1 _09589_ (.A(net1159),
    .B(_04344_),
    .X(_00259_));
 sky130_fd_sc_hd__a32o_1 _09590_ (.A1(net558),
    .A2(net388),
    .A3(net662),
    .B1(net378),
    .B2(\reg_module.gprf[158] ),
    .X(_04345_));
 sky130_fd_sc_hd__and2_1 _09591_ (.A(net1192),
    .B(_04345_),
    .X(_00260_));
 sky130_fd_sc_hd__a32o_1 _09592_ (.A1(net560),
    .A2(net387),
    .A3(net662),
    .B1(net378),
    .B2(\reg_module.gprf[159] ),
    .X(_04346_));
 sky130_fd_sc_hd__and2_1 _09593_ (.A(net1195),
    .B(_04346_),
    .X(_00261_));
 sky130_fd_sc_hd__and3_1 _09594_ (.A(_01213_),
    .B(net970),
    .C(_01214_),
    .X(_04347_));
 sky130_fd_sc_hd__nand3_4 _09595_ (.A(net967),
    .B(net536),
    .C(net650),
    .Y(_04348_));
 sky130_fd_sc_hd__a32o_1 _09596_ (.A1(net515),
    .A2(net418),
    .A3(net649),
    .B1(net371),
    .B2(\reg_module.gprf[160] ),
    .X(_04349_));
 sky130_fd_sc_hd__and2_1 _09597_ (.A(net1089),
    .B(_04349_),
    .X(_00262_));
 sky130_fd_sc_hd__a32o_1 _09598_ (.A1(net534),
    .A2(net417),
    .A3(net650),
    .B1(net372),
    .B2(\reg_module.gprf[161] ),
    .X(_04350_));
 sky130_fd_sc_hd__and2_1 _09599_ (.A(net1126),
    .B(_04350_),
    .X(_00263_));
 sky130_fd_sc_hd__a32o_1 _09600_ (.A1(net524),
    .A2(net416),
    .A3(net649),
    .B1(net371),
    .B2(\reg_module.gprf[162] ),
    .X(_04351_));
 sky130_fd_sc_hd__and2_1 _09601_ (.A(net1106),
    .B(_04351_),
    .X(_00264_));
 sky130_fd_sc_hd__a32o_1 _09602_ (.A1(net512),
    .A2(net415),
    .A3(net647),
    .B1(net371),
    .B2(\reg_module.gprf[163] ),
    .X(_04352_));
 sky130_fd_sc_hd__and2_1 _09603_ (.A(net1077),
    .B(_04352_),
    .X(_00265_));
 sky130_fd_sc_hd__a32o_1 _09604_ (.A1(net535),
    .A2(net414),
    .A3(net654),
    .B1(net372),
    .B2(\reg_module.gprf[164] ),
    .X(_04353_));
 sky130_fd_sc_hd__and2_1 _09605_ (.A(net1127),
    .B(_04353_),
    .X(_00266_));
 sky130_fd_sc_hd__a32o_1 _09606_ (.A1(net529),
    .A2(net413),
    .A3(net650),
    .B1(net372),
    .B2(\reg_module.gprf[165] ),
    .X(_04354_));
 sky130_fd_sc_hd__and2_1 _09607_ (.A(net1118),
    .B(_04354_),
    .X(_00267_));
 sky130_fd_sc_hd__a32o_1 _09608_ (.A1(net509),
    .A2(net412),
    .A3(net647),
    .B1(net371),
    .B2(\reg_module.gprf[166] ),
    .X(_04355_));
 sky130_fd_sc_hd__and2_1 _09609_ (.A(net1071),
    .B(_04355_),
    .X(_00268_));
 sky130_fd_sc_hd__a32o_1 _09610_ (.A1(net513),
    .A2(net411),
    .A3(net647),
    .B1(net371),
    .B2(\reg_module.gprf[167] ),
    .X(_04356_));
 sky130_fd_sc_hd__and2_1 _09611_ (.A(net1083),
    .B(_04356_),
    .X(_00269_));
 sky130_fd_sc_hd__a32o_1 _09612_ (.A1(net530),
    .A2(net410),
    .A3(net650),
    .B1(net372),
    .B2(\reg_module.gprf[168] ),
    .X(_04357_));
 sky130_fd_sc_hd__and2_1 _09613_ (.A(net1121),
    .B(_04357_),
    .X(_00270_));
 sky130_fd_sc_hd__a32o_1 _09614_ (.A1(net518),
    .A2(_04199_),
    .A3(net648),
    .B1(net372),
    .B2(\reg_module.gprf[169] ),
    .X(_04358_));
 sky130_fd_sc_hd__and2_1 _09615_ (.A(net1094),
    .B(_04358_),
    .X(_00271_));
 sky130_fd_sc_hd__a32o_1 _09616_ (.A1(net510),
    .A2(net408),
    .A3(net647),
    .B1(net371),
    .B2(\reg_module.gprf[170] ),
    .X(_04359_));
 sky130_fd_sc_hd__and2_1 _09617_ (.A(net1073),
    .B(_04359_),
    .X(_00272_));
 sky130_fd_sc_hd__a32o_1 _09618_ (.A1(net520),
    .A2(_04203_),
    .A3(net648),
    .B1(net371),
    .B2(\reg_module.gprf[171] ),
    .X(_04360_));
 sky130_fd_sc_hd__and2_1 _09619_ (.A(net1100),
    .B(_04360_),
    .X(_00273_));
 sky130_fd_sc_hd__a32o_1 _09620_ (.A1(net521),
    .A2(net406),
    .A3(net648),
    .B1(net372),
    .B2(\reg_module.gprf[172] ),
    .X(_04361_));
 sky130_fd_sc_hd__and2_1 _09621_ (.A(net1102),
    .B(_04361_),
    .X(_00274_));
 sky130_fd_sc_hd__a32o_1 _09622_ (.A1(net519),
    .A2(net405),
    .A3(net648),
    .B1(net371),
    .B2(\reg_module.gprf[173] ),
    .X(_04362_));
 sky130_fd_sc_hd__and2_1 _09623_ (.A(net1097),
    .B(_04362_),
    .X(_00275_));
 sky130_fd_sc_hd__a32o_1 _09624_ (.A1(net525),
    .A2(net404),
    .A3(net649),
    .B1(net371),
    .B2(\reg_module.gprf[174] ),
    .X(_04363_));
 sky130_fd_sc_hd__and2_1 _09625_ (.A(net1110),
    .B(_04363_),
    .X(_00276_));
 sky130_fd_sc_hd__a32o_1 _09626_ (.A1(net544),
    .A2(net403),
    .A3(net652),
    .B1(net373),
    .B2(\reg_module.gprf[175] ),
    .X(_04364_));
 sky130_fd_sc_hd__and2_1 _09627_ (.A(net1155),
    .B(_04364_),
    .X(_00277_));
 sky130_fd_sc_hd__a32o_1 _09628_ (.A1(net559),
    .A2(net402),
    .A3(net653),
    .B1(net374),
    .B2(\reg_module.gprf[176] ),
    .X(_04365_));
 sky130_fd_sc_hd__and2_1 _09629_ (.A(net1200),
    .B(_04365_),
    .X(_00278_));
 sky130_fd_sc_hd__a32o_1 _09630_ (.A1(net539),
    .A2(net401),
    .A3(net652),
    .B1(net373),
    .B2(\reg_module.gprf[177] ),
    .X(_04366_));
 sky130_fd_sc_hd__and2_1 _09631_ (.A(net1142),
    .B(_04366_),
    .X(_00279_));
 sky130_fd_sc_hd__a32o_1 _09632_ (.A1(net521),
    .A2(net400),
    .A3(net648),
    .B1(net371),
    .B2(\reg_module.gprf[178] ),
    .X(_04367_));
 sky130_fd_sc_hd__and2_1 _09633_ (.A(net1103),
    .B(_04367_),
    .X(_00280_));
 sky130_fd_sc_hd__a32o_1 _09634_ (.A1(net541),
    .A2(_04219_),
    .A3(net652),
    .B1(net373),
    .B2(\reg_module.gprf[179] ),
    .X(_04368_));
 sky130_fd_sc_hd__and2_1 _09635_ (.A(net1148),
    .B(_04368_),
    .X(_00281_));
 sky130_fd_sc_hd__a32o_1 _09636_ (.A1(net526),
    .A2(net398),
    .A3(net649),
    .B1(net372),
    .B2(\reg_module.gprf[180] ),
    .X(_04369_));
 sky130_fd_sc_hd__and2_1 _09637_ (.A(net1109),
    .B(_04369_),
    .X(_00282_));
 sky130_fd_sc_hd__a32o_1 _09638_ (.A1(net561),
    .A2(net397),
    .A3(net653),
    .B1(net374),
    .B2(\reg_module.gprf[181] ),
    .X(_04370_));
 sky130_fd_sc_hd__and2_1 _09639_ (.A(net1204),
    .B(_04370_),
    .X(_00283_));
 sky130_fd_sc_hd__a32o_1 _09640_ (.A1(net557),
    .A2(net396),
    .A3(net653),
    .B1(net374),
    .B2(\reg_module.gprf[182] ),
    .X(_04371_));
 sky130_fd_sc_hd__and2_1 _09641_ (.A(net1192),
    .B(_04371_),
    .X(_00284_));
 sky130_fd_sc_hd__a32o_1 _09642_ (.A1(net548),
    .A2(net395),
    .A3(net651),
    .B1(net373),
    .B2(\reg_module.gprf[183] ),
    .X(_04372_));
 sky130_fd_sc_hd__and2_1 _09643_ (.A(net1167),
    .B(_04372_),
    .X(_00285_));
 sky130_fd_sc_hd__a32o_1 _09644_ (.A1(net552),
    .A2(net394),
    .A3(net651),
    .B1(net373),
    .B2(\reg_module.gprf[184] ),
    .X(_04373_));
 sky130_fd_sc_hd__and2_1 _09645_ (.A(net1181),
    .B(_04373_),
    .X(_00286_));
 sky130_fd_sc_hd__a32o_1 _09646_ (.A1(net552),
    .A2(net393),
    .A3(net651),
    .B1(net373),
    .B2(\reg_module.gprf[185] ),
    .X(_04374_));
 sky130_fd_sc_hd__and2_1 _09647_ (.A(net1181),
    .B(_04374_),
    .X(_00287_));
 sky130_fd_sc_hd__a32o_1 _09648_ (.A1(net545),
    .A2(net392),
    .A3(net652),
    .B1(net373),
    .B2(\reg_module.gprf[186] ),
    .X(_04375_));
 sky130_fd_sc_hd__and2_1 _09649_ (.A(net1161),
    .B(_04375_),
    .X(_00288_));
 sky130_fd_sc_hd__a32o_1 _09650_ (.A1(net540),
    .A2(net391),
    .A3(net652),
    .B1(net373),
    .B2(\reg_module.gprf[187] ),
    .X(_04376_));
 sky130_fd_sc_hd__and2_1 _09651_ (.A(net1145),
    .B(_04376_),
    .X(_00289_));
 sky130_fd_sc_hd__a32o_1 _09652_ (.A1(net549),
    .A2(net390),
    .A3(net651),
    .B1(net373),
    .B2(\reg_module.gprf[188] ),
    .X(_04377_));
 sky130_fd_sc_hd__and2_1 _09653_ (.A(net1170),
    .B(_04377_),
    .X(_00290_));
 sky130_fd_sc_hd__a32o_1 _09654_ (.A1(net548),
    .A2(net389),
    .A3(net651),
    .B1(net373),
    .B2(\reg_module.gprf[189] ),
    .X(_04378_));
 sky130_fd_sc_hd__and2_1 _09655_ (.A(net1167),
    .B(_04378_),
    .X(_00291_));
 sky130_fd_sc_hd__a32o_1 _09656_ (.A1(net558),
    .A2(net388),
    .A3(net654),
    .B1(net374),
    .B2(\reg_module.gprf[190] ),
    .X(_04379_));
 sky130_fd_sc_hd__and2_1 _09657_ (.A(net1182),
    .B(_04379_),
    .X(_00292_));
 sky130_fd_sc_hd__a32o_1 _09658_ (.A1(net560),
    .A2(net387),
    .A3(net653),
    .B1(net374),
    .B2(\reg_module.gprf[191] ),
    .X(_04380_));
 sky130_fd_sc_hd__and2_1 _09659_ (.A(net1204),
    .B(_04380_),
    .X(_00293_));
 sky130_fd_sc_hd__or4b_4 _09660_ (.A(_01213_),
    .B(net969),
    .C(net968),
    .D_N(net967),
    .X(_04381_));
 sky130_fd_sc_hd__or2_2 _09661_ (.A(_04175_),
    .B(net644),
    .X(_04382_));
 sky130_fd_sc_hd__nor2_1 _09662_ (.A(_02685_),
    .B(net643),
    .Y(_04383_));
 sky130_fd_sc_hd__a22o_1 _09663_ (.A1(\reg_module.gprf[192] ),
    .A2(net367),
    .B1(_04383_),
    .B2(net516),
    .X(_04384_));
 sky130_fd_sc_hd__and2_1 _09664_ (.A(net1090),
    .B(_04384_),
    .X(_00294_));
 sky130_fd_sc_hd__nor2_1 _09665_ (.A(_02673_),
    .B(net644),
    .Y(_04385_));
 sky130_fd_sc_hd__a22o_1 _09666_ (.A1(\reg_module.gprf[193] ),
    .A2(net368),
    .B1(_04385_),
    .B2(net534),
    .X(_04386_));
 sky130_fd_sc_hd__and2_1 _09667_ (.A(net1128),
    .B(_04386_),
    .X(_00295_));
 sky130_fd_sc_hd__nor2_1 _09668_ (.A(net713),
    .B(net644),
    .Y(_04387_));
 sky130_fd_sc_hd__a22o_1 _09669_ (.A1(\reg_module.gprf[194] ),
    .A2(net368),
    .B1(_04387_),
    .B2(net524),
    .X(_04388_));
 sky130_fd_sc_hd__and2_1 _09670_ (.A(net1106),
    .B(_04388_),
    .X(_00296_));
 sky130_fd_sc_hd__nor2_1 _09671_ (.A(net712),
    .B(net643),
    .Y(_04389_));
 sky130_fd_sc_hd__a22o_1 _09672_ (.A1(\reg_module.gprf[195] ),
    .A2(net367),
    .B1(_04389_),
    .B2(net515),
    .X(_04390_));
 sky130_fd_sc_hd__and2_1 _09673_ (.A(net1078),
    .B(_04390_),
    .X(_00297_));
 sky130_fd_sc_hd__nor2_1 _09674_ (.A(net723),
    .B(net644),
    .Y(_04391_));
 sky130_fd_sc_hd__a22o_1 _09675_ (.A1(\reg_module.gprf[196] ),
    .A2(net368),
    .B1(_04391_),
    .B2(net535),
    .X(_04392_));
 sky130_fd_sc_hd__and2_1 _09676_ (.A(net1128),
    .B(_04392_),
    .X(_00298_));
 sky130_fd_sc_hd__nor2_1 _09677_ (.A(net722),
    .B(net644),
    .Y(_04393_));
 sky130_fd_sc_hd__a22o_1 _09678_ (.A1(\reg_module.gprf[197] ),
    .A2(net368),
    .B1(_04393_),
    .B2(net531),
    .X(_04394_));
 sky130_fd_sc_hd__and2_1 _09679_ (.A(net1120),
    .B(_04394_),
    .X(_00299_));
 sky130_fd_sc_hd__nor2_1 _09680_ (.A(net725),
    .B(net643),
    .Y(_04395_));
 sky130_fd_sc_hd__a22o_1 _09681_ (.A1(\reg_module.gprf[198] ),
    .A2(net367),
    .B1(_04395_),
    .B2(net510),
    .X(_04396_));
 sky130_fd_sc_hd__and2_1 _09682_ (.A(net1072),
    .B(_04396_),
    .X(_00300_));
 sky130_fd_sc_hd__nor2_1 _09683_ (.A(net724),
    .B(net643),
    .Y(_04397_));
 sky130_fd_sc_hd__a22o_1 _09684_ (.A1(\reg_module.gprf[199] ),
    .A2(net367),
    .B1(_04397_),
    .B2(net513),
    .X(_04398_));
 sky130_fd_sc_hd__and2_1 _09685_ (.A(net1082),
    .B(_04398_),
    .X(_00301_));
 sky130_fd_sc_hd__nor2_1 _09686_ (.A(_03077_),
    .B(net644),
    .Y(_04399_));
 sky130_fd_sc_hd__a22o_1 _09687_ (.A1(\reg_module.gprf[200] ),
    .A2(net368),
    .B1(_04399_),
    .B2(net531),
    .X(_04400_));
 sky130_fd_sc_hd__and2_1 _09688_ (.A(net1122),
    .B(_04400_),
    .X(_00302_));
 sky130_fd_sc_hd__nor2_1 _09689_ (.A(net690),
    .B(net643),
    .Y(_04401_));
 sky130_fd_sc_hd__a22o_1 _09690_ (.A1(\reg_module.gprf[201] ),
    .A2(net367),
    .B1(_04401_),
    .B2(net518),
    .X(_04402_));
 sky130_fd_sc_hd__and2_1 _09691_ (.A(net1096),
    .B(_04402_),
    .X(_00303_));
 sky130_fd_sc_hd__nor2_1 _09692_ (.A(_03030_),
    .B(net643),
    .Y(_04403_));
 sky130_fd_sc_hd__a22o_1 _09693_ (.A1(\reg_module.gprf[202] ),
    .A2(net367),
    .B1(_04403_),
    .B2(net509),
    .X(_04404_));
 sky130_fd_sc_hd__and2_1 _09694_ (.A(net1073),
    .B(_04404_),
    .X(_00304_));
 sky130_fd_sc_hd__nor2_1 _09695_ (.A(net691),
    .B(net643),
    .Y(_04405_));
 sky130_fd_sc_hd__a22o_1 _09696_ (.A1(\reg_module.gprf[203] ),
    .A2(net367),
    .B1(_04405_),
    .B2(net520),
    .X(_04406_));
 sky130_fd_sc_hd__and2_1 _09697_ (.A(net1100),
    .B(_04406_),
    .X(_00305_));
 sky130_fd_sc_hd__nor2_1 _09698_ (.A(net693),
    .B(net643),
    .Y(_04407_));
 sky130_fd_sc_hd__a22o_1 _09699_ (.A1(\reg_module.gprf[204] ),
    .A2(net367),
    .B1(_04407_),
    .B2(net521),
    .X(_04408_));
 sky130_fd_sc_hd__and2_1 _09700_ (.A(net1102),
    .B(_04408_),
    .X(_00306_));
 sky130_fd_sc_hd__nor2_1 _09701_ (.A(net694),
    .B(net643),
    .Y(_04409_));
 sky130_fd_sc_hd__a22o_1 _09702_ (.A1(\reg_module.gprf[205] ),
    .A2(net367),
    .B1(_04409_),
    .B2(net519),
    .X(_04410_));
 sky130_fd_sc_hd__and2_1 _09703_ (.A(net1098),
    .B(_04410_),
    .X(_00307_));
 sky130_fd_sc_hd__nor2_1 _09704_ (.A(net696),
    .B(net643),
    .Y(_04411_));
 sky130_fd_sc_hd__a22o_1 _09705_ (.A1(\reg_module.gprf[206] ),
    .A2(net367),
    .B1(_04411_),
    .B2(net527),
    .X(_04412_));
 sky130_fd_sc_hd__and2_1 _09706_ (.A(net1115),
    .B(_04412_),
    .X(_00308_));
 sky130_fd_sc_hd__nor2_1 _09707_ (.A(net695),
    .B(net645),
    .Y(_04413_));
 sky130_fd_sc_hd__a22o_1 _09708_ (.A1(\reg_module.gprf[207] ),
    .A2(net369),
    .B1(_04413_),
    .B2(net544),
    .X(_04414_));
 sky130_fd_sc_hd__and2_1 _09709_ (.A(net1155),
    .B(_04414_),
    .X(_00309_));
 sky130_fd_sc_hd__nor2_1 _09710_ (.A(net698),
    .B(net646),
    .Y(_04415_));
 sky130_fd_sc_hd__a22o_1 _09711_ (.A1(\reg_module.gprf[208] ),
    .A2(net370),
    .B1(_04415_),
    .B2(net563),
    .X(_04416_));
 sky130_fd_sc_hd__and2_1 _09712_ (.A(net1199),
    .B(_04416_),
    .X(_00310_));
 sky130_fd_sc_hd__nor2_1 _09713_ (.A(net697),
    .B(net645),
    .Y(_04417_));
 sky130_fd_sc_hd__a22o_1 _09714_ (.A1(\reg_module.gprf[209] ),
    .A2(net369),
    .B1(_04417_),
    .B2(net539),
    .X(_04418_));
 sky130_fd_sc_hd__and2_1 _09715_ (.A(net1142),
    .B(_04418_),
    .X(_00311_));
 sky130_fd_sc_hd__nor2_1 _09716_ (.A(net700),
    .B(net645),
    .Y(_04419_));
 sky130_fd_sc_hd__a22o_1 _09717_ (.A1(\reg_module.gprf[210] ),
    .A2(net369),
    .B1(_04419_),
    .B2(net542),
    .X(_04420_));
 sky130_fd_sc_hd__and2_1 _09718_ (.A(net1143),
    .B(_04420_),
    .X(_00312_));
 sky130_fd_sc_hd__nor2_1 _09719_ (.A(net699),
    .B(net645),
    .Y(_04421_));
 sky130_fd_sc_hd__a22o_1 _09720_ (.A1(\reg_module.gprf[211] ),
    .A2(net369),
    .B1(_04421_),
    .B2(net541),
    .X(_04422_));
 sky130_fd_sc_hd__and2_1 _09721_ (.A(net1148),
    .B(_04422_),
    .X(_00313_));
 sky130_fd_sc_hd__nor2_1 _09722_ (.A(net702),
    .B(net644),
    .Y(_04423_));
 sky130_fd_sc_hd__a22o_1 _09723_ (.A1(\reg_module.gprf[212] ),
    .A2(net368),
    .B1(_04423_),
    .B2(net526),
    .X(_04424_));
 sky130_fd_sc_hd__and2_1 _09724_ (.A(net1113),
    .B(_04424_),
    .X(_00314_));
 sky130_fd_sc_hd__nor2_1 _09725_ (.A(net701),
    .B(net646),
    .Y(_04425_));
 sky130_fd_sc_hd__a22o_1 _09726_ (.A1(\reg_module.gprf[213] ),
    .A2(net370),
    .B1(_04425_),
    .B2(net561),
    .X(_04426_));
 sky130_fd_sc_hd__and2_1 _09727_ (.A(net1206),
    .B(_04426_),
    .X(_00315_));
 sky130_fd_sc_hd__nor2_1 _09728_ (.A(net704),
    .B(net646),
    .Y(_04427_));
 sky130_fd_sc_hd__a22o_1 _09729_ (.A1(\reg_module.gprf[214] ),
    .A2(net370),
    .B1(_04427_),
    .B2(net557),
    .X(_04428_));
 sky130_fd_sc_hd__and2_1 _09730_ (.A(net1192),
    .B(_04428_),
    .X(_00316_));
 sky130_fd_sc_hd__nor2_1 _09731_ (.A(_02864_),
    .B(net645),
    .Y(_04429_));
 sky130_fd_sc_hd__a22o_1 _09732_ (.A1(\reg_module.gprf[215] ),
    .A2(net369),
    .B1(_04429_),
    .B2(net548),
    .X(_04430_));
 sky130_fd_sc_hd__and2_1 _09733_ (.A(net1168),
    .B(_04430_),
    .X(_00317_));
 sky130_fd_sc_hd__nor2_1 _09734_ (.A(net705),
    .B(net645),
    .Y(_04431_));
 sky130_fd_sc_hd__a22o_1 _09735_ (.A1(\reg_module.gprf[216] ),
    .A2(net369),
    .B1(_04431_),
    .B2(net552),
    .X(_04432_));
 sky130_fd_sc_hd__and2_1 _09736_ (.A(net1181),
    .B(_04432_),
    .X(_00318_));
 sky130_fd_sc_hd__nor2_1 _09737_ (.A(net706),
    .B(net645),
    .Y(_04433_));
 sky130_fd_sc_hd__a22o_1 _09738_ (.A1(\reg_module.gprf[217] ),
    .A2(net369),
    .B1(_04433_),
    .B2(net552),
    .X(_04434_));
 sky130_fd_sc_hd__and2_1 _09739_ (.A(net1173),
    .B(_04434_),
    .X(_00319_));
 sky130_fd_sc_hd__nor2_1 _09740_ (.A(net708),
    .B(net645),
    .Y(_04435_));
 sky130_fd_sc_hd__a22o_1 _09741_ (.A1(\reg_module.gprf[218] ),
    .A2(net369),
    .B1(_04435_),
    .B2(net545),
    .X(_04436_));
 sky130_fd_sc_hd__and2_1 _09742_ (.A(net1161),
    .B(_04436_),
    .X(_00320_));
 sky130_fd_sc_hd__nor2_1 _09743_ (.A(net707),
    .B(net646),
    .Y(_04437_));
 sky130_fd_sc_hd__a22o_1 _09744_ (.A1(\reg_module.gprf[219] ),
    .A2(net370),
    .B1(_04437_),
    .B2(net541),
    .X(_04438_));
 sky130_fd_sc_hd__and2_1 _09745_ (.A(net1149),
    .B(_04438_),
    .X(_00321_));
 sky130_fd_sc_hd__nor2_1 _09746_ (.A(net710),
    .B(net646),
    .Y(_04439_));
 sky130_fd_sc_hd__a22o_1 _09747_ (.A1(\reg_module.gprf[220] ),
    .A2(net369),
    .B1(_04439_),
    .B2(net550),
    .X(_04440_));
 sky130_fd_sc_hd__and2_1 _09748_ (.A(net1171),
    .B(_04440_),
    .X(_00322_));
 sky130_fd_sc_hd__nor2_1 _09749_ (.A(net709),
    .B(net645),
    .Y(_04441_));
 sky130_fd_sc_hd__a22o_1 _09750_ (.A1(\reg_module.gprf[221] ),
    .A2(net370),
    .B1(_04441_),
    .B2(net551),
    .X(_04442_));
 sky130_fd_sc_hd__and2_1 _09751_ (.A(net1175),
    .B(_04442_),
    .X(_00323_));
 sky130_fd_sc_hd__nor2_1 _09752_ (.A(net711),
    .B(net645),
    .Y(_04443_));
 sky130_fd_sc_hd__a22o_1 _09753_ (.A1(\reg_module.gprf[222] ),
    .A2(net369),
    .B1(_04443_),
    .B2(net554),
    .X(_04444_));
 sky130_fd_sc_hd__and2_1 _09754_ (.A(net1182),
    .B(_04444_),
    .X(_00324_));
 sky130_fd_sc_hd__nor2_1 _09755_ (.A(net574),
    .B(net646),
    .Y(_04445_));
 sky130_fd_sc_hd__a22o_1 _09756_ (.A1(\reg_module.gprf[223] ),
    .A2(net370),
    .B1(_04445_),
    .B2(net560),
    .X(_04446_));
 sky130_fd_sc_hd__and2_1 _09757_ (.A(net1195),
    .B(_04446_),
    .X(_00325_));
 sky130_fd_sc_hd__nand3_4 _09758_ (.A(net967),
    .B(net777),
    .C(net536),
    .Y(_04447_));
 sky130_fd_sc_hd__a32o_1 _09759_ (.A1(net776),
    .A2(net516),
    .A3(net418),
    .B1(net363),
    .B2(\reg_module.gprf[224] ),
    .X(_04448_));
 sky130_fd_sc_hd__and2_1 _09760_ (.A(net1090),
    .B(_04448_),
    .X(_00326_));
 sky130_fd_sc_hd__a32o_1 _09761_ (.A1(_01253_),
    .A2(net533),
    .A3(net417),
    .B1(net364),
    .B2(\reg_module.gprf[225] ),
    .X(_04449_));
 sky130_fd_sc_hd__and2_1 _09762_ (.A(net1128),
    .B(_04449_),
    .X(_00327_));
 sky130_fd_sc_hd__a32o_1 _09763_ (.A1(net775),
    .A2(net524),
    .A3(_04185_),
    .B1(net363),
    .B2(\reg_module.gprf[226] ),
    .X(_04450_));
 sky130_fd_sc_hd__and2_1 _09764_ (.A(net1106),
    .B(_04450_),
    .X(_00328_));
 sky130_fd_sc_hd__a32o_1 _09765_ (.A1(net774),
    .A2(net512),
    .A3(net415),
    .B1(net363),
    .B2(\reg_module.gprf[227] ),
    .X(_04451_));
 sky130_fd_sc_hd__and2_1 _09766_ (.A(net1078),
    .B(_04451_),
    .X(_00329_));
 sky130_fd_sc_hd__a32o_1 _09767_ (.A1(net777),
    .A2(net535),
    .A3(_04189_),
    .B1(net364),
    .B2(\reg_module.gprf[228] ),
    .X(_04452_));
 sky130_fd_sc_hd__and2_1 _09768_ (.A(net1128),
    .B(_04452_),
    .X(_00330_));
 sky130_fd_sc_hd__a32o_1 _09769_ (.A1(net777),
    .A2(net531),
    .A3(net413),
    .B1(net364),
    .B2(\reg_module.gprf[229] ),
    .X(_04453_));
 sky130_fd_sc_hd__and2_1 _09770_ (.A(net1120),
    .B(_04453_),
    .X(_00331_));
 sky130_fd_sc_hd__a32o_1 _09771_ (.A1(net774),
    .A2(net509),
    .A3(_04193_),
    .B1(net363),
    .B2(\reg_module.gprf[230] ),
    .X(_04454_));
 sky130_fd_sc_hd__and2_1 _09772_ (.A(net1072),
    .B(_04454_),
    .X(_00332_));
 sky130_fd_sc_hd__a32o_1 _09773_ (.A1(net774),
    .A2(net513),
    .A3(_04195_),
    .B1(net363),
    .B2(\reg_module.gprf[231] ),
    .X(_04455_));
 sky130_fd_sc_hd__and2_1 _09774_ (.A(net1082),
    .B(_04455_),
    .X(_00333_));
 sky130_fd_sc_hd__a32o_1 _09775_ (.A1(net777),
    .A2(net530),
    .A3(net410),
    .B1(net364),
    .B2(\reg_module.gprf[232] ),
    .X(_04456_));
 sky130_fd_sc_hd__and2_1 _09776_ (.A(net1122),
    .B(_04456_),
    .X(_00334_));
 sky130_fd_sc_hd__a32o_1 _09777_ (.A1(net775),
    .A2(net518),
    .A3(net409),
    .B1(net364),
    .B2(\reg_module.gprf[233] ),
    .X(_04457_));
 sky130_fd_sc_hd__and2_1 _09778_ (.A(net1095),
    .B(_04457_),
    .X(_00335_));
 sky130_fd_sc_hd__a32o_1 _09779_ (.A1(net774),
    .A2(net511),
    .A3(net408),
    .B1(net363),
    .B2(\reg_module.gprf[234] ),
    .X(_04458_));
 sky130_fd_sc_hd__and2_1 _09780_ (.A(net1074),
    .B(_04458_),
    .X(_00336_));
 sky130_fd_sc_hd__a32o_1 _09781_ (.A1(net775),
    .A2(net522),
    .A3(net407),
    .B1(net363),
    .B2(\reg_module.gprf[235] ),
    .X(_04459_));
 sky130_fd_sc_hd__and2_1 _09782_ (.A(net1103),
    .B(_04459_),
    .X(_00337_));
 sky130_fd_sc_hd__a32o_1 _09783_ (.A1(net775),
    .A2(net521),
    .A3(net406),
    .B1(net364),
    .B2(\reg_module.gprf[236] ),
    .X(_04460_));
 sky130_fd_sc_hd__and2_1 _09784_ (.A(net1102),
    .B(_04460_),
    .X(_00338_));
 sky130_fd_sc_hd__a32o_1 _09785_ (.A1(net775),
    .A2(net519),
    .A3(net405),
    .B1(net363),
    .B2(\reg_module.gprf[237] ),
    .X(_04461_));
 sky130_fd_sc_hd__and2_1 _09786_ (.A(net1098),
    .B(_04461_),
    .X(_00339_));
 sky130_fd_sc_hd__a32o_1 _09787_ (.A1(net775),
    .A2(net527),
    .A3(net404),
    .B1(net363),
    .B2(\reg_module.gprf[238] ),
    .X(_04462_));
 sky130_fd_sc_hd__and2_1 _09788_ (.A(net1110),
    .B(_04462_),
    .X(_00340_));
 sky130_fd_sc_hd__a32o_1 _09789_ (.A1(net778),
    .A2(net544),
    .A3(net403),
    .B1(net365),
    .B2(\reg_module.gprf[239] ),
    .X(_04463_));
 sky130_fd_sc_hd__and2_1 _09790_ (.A(net1156),
    .B(_04463_),
    .X(_00341_));
 sky130_fd_sc_hd__a32o_1 _09791_ (.A1(net781),
    .A2(net559),
    .A3(_04213_),
    .B1(net366),
    .B2(\reg_module.gprf[240] ),
    .X(_04464_));
 sky130_fd_sc_hd__and2_1 _09792_ (.A(net1199),
    .B(_04464_),
    .X(_00342_));
 sky130_fd_sc_hd__a32o_1 _09793_ (.A1(net778),
    .A2(net539),
    .A3(net401),
    .B1(net365),
    .B2(\reg_module.gprf[241] ),
    .X(_04465_));
 sky130_fd_sc_hd__and2_1 _09794_ (.A(net1142),
    .B(_04465_),
    .X(_00343_));
 sky130_fd_sc_hd__a32o_1 _09795_ (.A1(net778),
    .A2(net538),
    .A3(_04217_),
    .B1(net365),
    .B2(\reg_module.gprf[242] ),
    .X(_04466_));
 sky130_fd_sc_hd__and2_1 _09796_ (.A(net1141),
    .B(_04466_),
    .X(_00344_));
 sky130_fd_sc_hd__a32o_1 _09797_ (.A1(net778),
    .A2(net541),
    .A3(_04219_),
    .B1(net365),
    .B2(\reg_module.gprf[243] ),
    .X(_04467_));
 sky130_fd_sc_hd__and2_1 _09798_ (.A(net1149),
    .B(_04467_),
    .X(_00345_));
 sky130_fd_sc_hd__a32o_1 _09799_ (.A1(net776),
    .A2(net526),
    .A3(net398),
    .B1(net363),
    .B2(\reg_module.gprf[244] ),
    .X(_04468_));
 sky130_fd_sc_hd__and2_1 _09800_ (.A(net1113),
    .B(_04468_),
    .X(_00346_));
 sky130_fd_sc_hd__a32o_1 _09801_ (.A1(net781),
    .A2(net562),
    .A3(_04223_),
    .B1(net366),
    .B2(\reg_module.gprf[245] ),
    .X(_04469_));
 sky130_fd_sc_hd__and2_1 _09802_ (.A(net1206),
    .B(_04469_),
    .X(_00347_));
 sky130_fd_sc_hd__a32o_1 _09803_ (.A1(net781),
    .A2(net557),
    .A3(net396),
    .B1(net366),
    .B2(\reg_module.gprf[246] ),
    .X(_04470_));
 sky130_fd_sc_hd__and2_1 _09804_ (.A(net1194),
    .B(_04470_),
    .X(_00348_));
 sky130_fd_sc_hd__a32o_1 _09805_ (.A1(net779),
    .A2(net548),
    .A3(net395),
    .B1(net365),
    .B2(\reg_module.gprf[247] ),
    .X(_04471_));
 sky130_fd_sc_hd__and2_1 _09806_ (.A(net1167),
    .B(_04471_),
    .X(_00349_));
 sky130_fd_sc_hd__a32o_1 _09807_ (.A1(net780),
    .A2(net552),
    .A3(_04229_),
    .B1(net365),
    .B2(\reg_module.gprf[248] ),
    .X(_04472_));
 sky130_fd_sc_hd__and2_1 _09808_ (.A(net1181),
    .B(_04472_),
    .X(_00350_));
 sky130_fd_sc_hd__a32o_1 _09809_ (.A1(net779),
    .A2(net552),
    .A3(net393),
    .B1(net365),
    .B2(\reg_module.gprf[249] ),
    .X(_04473_));
 sky130_fd_sc_hd__and2_1 _09810_ (.A(net1181),
    .B(_04473_),
    .X(_00351_));
 sky130_fd_sc_hd__a32o_1 _09811_ (.A1(net778),
    .A2(net545),
    .A3(net392),
    .B1(net365),
    .B2(\reg_module.gprf[250] ),
    .X(_04474_));
 sky130_fd_sc_hd__and2_1 _09812_ (.A(net1161),
    .B(_04474_),
    .X(_00352_));
 sky130_fd_sc_hd__a32o_1 _09813_ (.A1(net778),
    .A2(net540),
    .A3(net391),
    .B1(net365),
    .B2(\reg_module.gprf[251] ),
    .X(_04475_));
 sky130_fd_sc_hd__and2_1 _09814_ (.A(net1146),
    .B(_04475_),
    .X(_00353_));
 sky130_fd_sc_hd__a32o_1 _09815_ (.A1(net779),
    .A2(net549),
    .A3(net390),
    .B1(net365),
    .B2(\reg_module.gprf[252] ),
    .X(_04476_));
 sky130_fd_sc_hd__and2_1 _09816_ (.A(net1170),
    .B(_04476_),
    .X(_00354_));
 sky130_fd_sc_hd__a32o_1 _09817_ (.A1(net779),
    .A2(net548),
    .A3(net389),
    .B1(net366),
    .B2(\reg_module.gprf[253] ),
    .X(_04477_));
 sky130_fd_sc_hd__and2_1 _09818_ (.A(net1167),
    .B(_04477_),
    .X(_00355_));
 sky130_fd_sc_hd__a32o_1 _09819_ (.A1(net780),
    .A2(net555),
    .A3(net388),
    .B1(net366),
    .B2(\reg_module.gprf[254] ),
    .X(_04478_));
 sky130_fd_sc_hd__and2_1 _09820_ (.A(net1182),
    .B(_04478_),
    .X(_00356_));
 sky130_fd_sc_hd__a32o_1 _09821_ (.A1(net781),
    .A2(net560),
    .A3(net387),
    .B1(net366),
    .B2(\reg_module.gprf[255] ),
    .X(_04479_));
 sky130_fd_sc_hd__and2_1 _09822_ (.A(net1195),
    .B(_04479_),
    .X(_00357_));
 sky130_fd_sc_hd__nor2_4 _09823_ (.A(_04175_),
    .B(_04178_),
    .Y(_04480_));
 sky130_fd_sc_hd__or2_1 _09824_ (.A(\reg_module.gprf[256] ),
    .B(net358),
    .X(_04481_));
 sky130_fd_sc_hd__o311a_1 _09825_ (.A1(_02686_),
    .A2(_04175_),
    .A3(_04178_),
    .B1(_04481_),
    .C1(net1125),
    .X(_00358_));
 sky130_fd_sc_hd__nand2_1 _09826_ (.A(net721),
    .B(net358),
    .Y(_04482_));
 sky130_fd_sc_hd__o211a_1 _09827_ (.A1(net1387),
    .A2(net358),
    .B1(_04482_),
    .C1(net1129),
    .X(_00359_));
 sky130_fd_sc_hd__nand2_1 _09828_ (.A(net713),
    .B(net357),
    .Y(_04483_));
 sky130_fd_sc_hd__o211a_1 _09829_ (.A1(net1346),
    .A2(net357),
    .B1(_04483_),
    .C1(net1109),
    .X(_00360_));
 sky130_fd_sc_hd__nand2_1 _09830_ (.A(net712),
    .B(net356),
    .Y(_04484_));
 sky130_fd_sc_hd__o211a_1 _09831_ (.A1(net1392),
    .A2(net356),
    .B1(_04484_),
    .C1(net1088),
    .X(_00361_));
 sky130_fd_sc_hd__nand2_1 _09832_ (.A(net723),
    .B(net358),
    .Y(_04485_));
 sky130_fd_sc_hd__o211a_1 _09833_ (.A1(net1386),
    .A2(net358),
    .B1(_04485_),
    .C1(net1126),
    .X(_00362_));
 sky130_fd_sc_hd__nand2_1 _09834_ (.A(net722),
    .B(net358),
    .Y(_04486_));
 sky130_fd_sc_hd__o211a_1 _09835_ (.A1(net1385),
    .A2(_04480_),
    .B1(_04486_),
    .C1(net1118),
    .X(_00363_));
 sky130_fd_sc_hd__nand2_1 _09836_ (.A(net725),
    .B(net356),
    .Y(_04487_));
 sky130_fd_sc_hd__o211a_1 _09837_ (.A1(net1404),
    .A2(net356),
    .B1(_04487_),
    .C1(net1071),
    .X(_00364_));
 sky130_fd_sc_hd__nand2_1 _09838_ (.A(net724),
    .B(net356),
    .Y(_04488_));
 sky130_fd_sc_hd__o211a_1 _09839_ (.A1(net1362),
    .A2(net356),
    .B1(_04488_),
    .C1(net1084),
    .X(_00365_));
 sky130_fd_sc_hd__nand2_1 _09840_ (.A(net689),
    .B(net358),
    .Y(_04489_));
 sky130_fd_sc_hd__o211a_1 _09841_ (.A1(net1384),
    .A2(net358),
    .B1(_04489_),
    .C1(net1121),
    .X(_00366_));
 sky130_fd_sc_hd__nand2_1 _09842_ (.A(net690),
    .B(net357),
    .Y(_04490_));
 sky130_fd_sc_hd__o211a_1 _09843_ (.A1(net1428),
    .A2(net357),
    .B1(_04490_),
    .C1(net1094),
    .X(_00367_));
 sky130_fd_sc_hd__nand2_1 _09844_ (.A(net692),
    .B(net356),
    .Y(_04491_));
 sky130_fd_sc_hd__o211a_1 _09845_ (.A1(net1355),
    .A2(net356),
    .B1(_04491_),
    .C1(net1074),
    .X(_00368_));
 sky130_fd_sc_hd__nand2_1 _09846_ (.A(net691),
    .B(net357),
    .Y(_04492_));
 sky130_fd_sc_hd__o211a_1 _09847_ (.A1(net1406),
    .A2(net357),
    .B1(_04492_),
    .C1(net1099),
    .X(_00369_));
 sky130_fd_sc_hd__nand2_1 _09848_ (.A(net693),
    .B(net359),
    .Y(_04493_));
 sky130_fd_sc_hd__o211a_1 _09849_ (.A1(net1380),
    .A2(net359),
    .B1(_04493_),
    .C1(net1103),
    .X(_00370_));
 sky130_fd_sc_hd__nand2_1 _09850_ (.A(_03000_),
    .B(net356),
    .Y(_04494_));
 sky130_fd_sc_hd__o211a_1 _09851_ (.A1(net1348),
    .A2(net356),
    .B1(_04494_),
    .C1(net1106),
    .X(_00371_));
 sky130_fd_sc_hd__nand2_1 _09852_ (.A(net696),
    .B(net361),
    .Y(_04495_));
 sky130_fd_sc_hd__o211a_1 _09853_ (.A1(net1379),
    .A2(net359),
    .B1(_04495_),
    .C1(net1155),
    .X(_00372_));
 sky130_fd_sc_hd__nand2_1 _09854_ (.A(net695),
    .B(net359),
    .Y(_04496_));
 sky130_fd_sc_hd__o211a_1 _09855_ (.A1(net1435),
    .A2(net361),
    .B1(_04496_),
    .C1(net1154),
    .X(_00373_));
 sky130_fd_sc_hd__nand2_1 _09856_ (.A(net698),
    .B(net362),
    .Y(_04497_));
 sky130_fd_sc_hd__o211a_1 _09857_ (.A1(net1417),
    .A2(net362),
    .B1(_04497_),
    .C1(net1202),
    .X(_00374_));
 sky130_fd_sc_hd__nand2_1 _09858_ (.A(net697),
    .B(net359),
    .Y(_04498_));
 sky130_fd_sc_hd__o211a_1 _09859_ (.A1(net1409),
    .A2(net359),
    .B1(_04498_),
    .C1(net1140),
    .X(_00375_));
 sky130_fd_sc_hd__nand2_1 _09860_ (.A(net700),
    .B(net359),
    .Y(_04499_));
 sky130_fd_sc_hd__o211a_1 _09861_ (.A1(net1353),
    .A2(net359),
    .B1(_04499_),
    .C1(net1139),
    .X(_00376_));
 sky130_fd_sc_hd__nand2_1 _09862_ (.A(net699),
    .B(net359),
    .Y(_04500_));
 sky130_fd_sc_hd__o211a_1 _09863_ (.A1(net1396),
    .A2(net359),
    .B1(_04500_),
    .C1(net1159),
    .X(_00377_));
 sky130_fd_sc_hd__nand2_1 _09864_ (.A(net702),
    .B(net357),
    .Y(_04501_));
 sky130_fd_sc_hd__o211a_1 _09865_ (.A1(net1422),
    .A2(net357),
    .B1(_04501_),
    .C1(net1114),
    .X(_00378_));
 sky130_fd_sc_hd__nand2_1 _09866_ (.A(net701),
    .B(net362),
    .Y(_04502_));
 sky130_fd_sc_hd__o211a_1 _09867_ (.A1(net1383),
    .A2(net362),
    .B1(_04502_),
    .C1(net1207),
    .X(_00379_));
 sky130_fd_sc_hd__nand2_1 _09868_ (.A(net704),
    .B(net362),
    .Y(_04503_));
 sky130_fd_sc_hd__o211a_1 _09869_ (.A1(net1375),
    .A2(net362),
    .B1(_04503_),
    .C1(net1193),
    .X(_00380_));
 sky130_fd_sc_hd__nand2_1 _09870_ (.A(net703),
    .B(net360),
    .Y(_04504_));
 sky130_fd_sc_hd__o211a_1 _09871_ (.A1(net1369),
    .A2(net360),
    .B1(_04504_),
    .C1(net1165),
    .X(_00381_));
 sky130_fd_sc_hd__nand2_1 _09872_ (.A(net705),
    .B(net360),
    .Y(_04505_));
 sky130_fd_sc_hd__o211a_1 _09873_ (.A1(net1408),
    .A2(net360),
    .B1(_04505_),
    .C1(net1180),
    .X(_00382_));
 sky130_fd_sc_hd__nand2_1 _09874_ (.A(net706),
    .B(net360),
    .Y(_04506_));
 sky130_fd_sc_hd__o211a_1 _09875_ (.A1(net1403),
    .A2(net360),
    .B1(_04506_),
    .C1(net1180),
    .X(_00383_));
 sky130_fd_sc_hd__nand2_1 _09876_ (.A(net708),
    .B(net361),
    .Y(_04507_));
 sky130_fd_sc_hd__o211a_1 _09877_ (.A1(net1423),
    .A2(net361),
    .B1(_04507_),
    .C1(net1159),
    .X(_00384_));
 sky130_fd_sc_hd__nand2_1 _09878_ (.A(net707),
    .B(net360),
    .Y(_04508_));
 sky130_fd_sc_hd__o211a_1 _09879_ (.A1(net1368),
    .A2(net360),
    .B1(_04508_),
    .C1(net1164),
    .X(_00385_));
 sky130_fd_sc_hd__nand2_1 _09880_ (.A(net710),
    .B(net360),
    .Y(_04509_));
 sky130_fd_sc_hd__o211a_1 _09881_ (.A1(net1360),
    .A2(net360),
    .B1(_04509_),
    .C1(net1170),
    .X(_00386_));
 sky130_fd_sc_hd__nand2_1 _09882_ (.A(net709),
    .B(net361),
    .Y(_04510_));
 sky130_fd_sc_hd__o211a_1 _09883_ (.A1(net1398),
    .A2(net361),
    .B1(_04510_),
    .C1(net1178),
    .X(_00387_));
 sky130_fd_sc_hd__nand2_1 _09884_ (.A(net711),
    .B(_04480_),
    .Y(_04511_));
 sky130_fd_sc_hd__o211a_1 _09885_ (.A1(net1399),
    .A2(net362),
    .B1(_04511_),
    .C1(net1193),
    .X(_00388_));
 sky130_fd_sc_hd__nand2_1 _09886_ (.A(net574),
    .B(net362),
    .Y(_04512_));
 sky130_fd_sc_hd__o211a_1 _09887_ (.A1(net1424),
    .A2(net362),
    .B1(_04512_),
    .C1(net1205),
    .X(_00389_));
 sky130_fd_sc_hd__nand2b_4 _09888_ (.A_N(net965),
    .B(net674),
    .Y(_04513_));
 sky130_fd_sc_hd__or2_1 _09889_ (.A(_04175_),
    .B(net502),
    .X(_04514_));
 sky130_fd_sc_hd__nor2_1 _09890_ (.A(_02685_),
    .B(net502),
    .Y(_04515_));
 sky130_fd_sc_hd__a22o_1 _09891_ (.A1(\reg_module.gprf[288] ),
    .A2(net355),
    .B1(_04515_),
    .B2(net532),
    .X(_04516_));
 sky130_fd_sc_hd__and2_1 _09892_ (.A(net1124),
    .B(_04516_),
    .X(_00390_));
 sky130_fd_sc_hd__nor2_1 _09893_ (.A(net721),
    .B(net502),
    .Y(_04517_));
 sky130_fd_sc_hd__a22o_1 _09894_ (.A1(\reg_module.gprf[289] ),
    .A2(net352),
    .B1(_04517_),
    .B2(net533),
    .X(_04518_));
 sky130_fd_sc_hd__and2_1 _09895_ (.A(net1129),
    .B(_04518_),
    .X(_00391_));
 sky130_fd_sc_hd__nor2_1 _09896_ (.A(net713),
    .B(net501),
    .Y(_04519_));
 sky130_fd_sc_hd__a22o_1 _09897_ (.A1(\reg_module.gprf[290] ),
    .A2(net352),
    .B1(_04519_),
    .B2(net525),
    .X(_04520_));
 sky130_fd_sc_hd__and2_1 _09898_ (.A(net1109),
    .B(_04520_),
    .X(_00392_));
 sky130_fd_sc_hd__nor2_1 _09899_ (.A(net712),
    .B(net501),
    .Y(_04521_));
 sky130_fd_sc_hd__a22o_1 _09900_ (.A1(\reg_module.gprf[291] ),
    .A2(net352),
    .B1(_04521_),
    .B2(net515),
    .X(_04522_));
 sky130_fd_sc_hd__and2_1 _09901_ (.A(net1087),
    .B(_04522_),
    .X(_00393_));
 sky130_fd_sc_hd__nor2_1 _09902_ (.A(net723),
    .B(net502),
    .Y(_04523_));
 sky130_fd_sc_hd__a22o_1 _09903_ (.A1(\reg_module.gprf[292] ),
    .A2(net355),
    .B1(_04523_),
    .B2(net533),
    .X(_04524_));
 sky130_fd_sc_hd__and2_1 _09904_ (.A(net1127),
    .B(_04524_),
    .X(_00394_));
 sky130_fd_sc_hd__nor2_1 _09905_ (.A(net722),
    .B(net502),
    .Y(_04525_));
 sky130_fd_sc_hd__a22o_1 _09906_ (.A1(\reg_module.gprf[293] ),
    .A2(net355),
    .B1(_04525_),
    .B2(net529),
    .X(_04526_));
 sky130_fd_sc_hd__and2_1 _09907_ (.A(net1118),
    .B(_04526_),
    .X(_00395_));
 sky130_fd_sc_hd__nor2_1 _09908_ (.A(net725),
    .B(net501),
    .Y(_04527_));
 sky130_fd_sc_hd__a22o_1 _09909_ (.A1(\reg_module.gprf[294] ),
    .A2(net352),
    .B1(_04527_),
    .B2(net509),
    .X(_04528_));
 sky130_fd_sc_hd__and2_1 _09910_ (.A(net1071),
    .B(_04528_),
    .X(_00396_));
 sky130_fd_sc_hd__nor2_1 _09911_ (.A(net724),
    .B(net501),
    .Y(_04529_));
 sky130_fd_sc_hd__a22o_1 _09912_ (.A1(\reg_module.gprf[295] ),
    .A2(net352),
    .B1(_04529_),
    .B2(net514),
    .X(_04530_));
 sky130_fd_sc_hd__and2_1 _09913_ (.A(net1084),
    .B(_04530_),
    .X(_00397_));
 sky130_fd_sc_hd__nor2_1 _09914_ (.A(net689),
    .B(net502),
    .Y(_04531_));
 sky130_fd_sc_hd__a22o_1 _09915_ (.A1(\reg_module.gprf[296] ),
    .A2(net355),
    .B1(_04531_),
    .B2(net530),
    .X(_04532_));
 sky130_fd_sc_hd__and2_1 _09916_ (.A(net1121),
    .B(_04532_),
    .X(_00398_));
 sky130_fd_sc_hd__nor2_1 _09917_ (.A(net690),
    .B(net501),
    .Y(_04533_));
 sky130_fd_sc_hd__a22o_1 _09918_ (.A1(\reg_module.gprf[297] ),
    .A2(net352),
    .B1(_04533_),
    .B2(net518),
    .X(_04534_));
 sky130_fd_sc_hd__and2_1 _09919_ (.A(net1094),
    .B(_04534_),
    .X(_00399_));
 sky130_fd_sc_hd__nor2_1 _09920_ (.A(net692),
    .B(net501),
    .Y(_04535_));
 sky130_fd_sc_hd__a22o_1 _09921_ (.A1(\reg_module.gprf[298] ),
    .A2(net352),
    .B1(_04535_),
    .B2(net511),
    .X(_04536_));
 sky130_fd_sc_hd__and2_1 _09922_ (.A(net1074),
    .B(_04536_),
    .X(_00400_));
 sky130_fd_sc_hd__nor2_1 _09923_ (.A(net691),
    .B(net501),
    .Y(_04537_));
 sky130_fd_sc_hd__a22o_1 _09924_ (.A1(\reg_module.gprf[299] ),
    .A2(net352),
    .B1(_04537_),
    .B2(net520),
    .X(_04538_));
 sky130_fd_sc_hd__and2_1 _09925_ (.A(net1099),
    .B(_04538_),
    .X(_00401_));
 sky130_fd_sc_hd__nor2_1 _09926_ (.A(net693),
    .B(net503),
    .Y(_04539_));
 sky130_fd_sc_hd__a22o_1 _09927_ (.A1(\reg_module.gprf[300] ),
    .A2(net353),
    .B1(_04539_),
    .B2(net521),
    .X(_04540_));
 sky130_fd_sc_hd__and2_1 _09928_ (.A(net1104),
    .B(_04540_),
    .X(_00402_));
 sky130_fd_sc_hd__nor2_1 _09929_ (.A(net694),
    .B(net501),
    .Y(_04541_));
 sky130_fd_sc_hd__a22o_1 _09930_ (.A1(\reg_module.gprf[301] ),
    .A2(net352),
    .B1(_04541_),
    .B2(net515),
    .X(_04542_));
 sky130_fd_sc_hd__and2_1 _09931_ (.A(net1088),
    .B(_04542_),
    .X(_00403_));
 sky130_fd_sc_hd__nor2_1 _09932_ (.A(net696),
    .B(net501),
    .Y(_04543_));
 sky130_fd_sc_hd__a22o_1 _09933_ (.A1(\reg_module.gprf[302] ),
    .A2(net353),
    .B1(_04543_),
    .B2(net527),
    .X(_04544_));
 sky130_fd_sc_hd__and2_1 _09934_ (.A(net1116),
    .B(_04544_),
    .X(_00404_));
 sky130_fd_sc_hd__nor2_1 _09935_ (.A(net695),
    .B(net503),
    .Y(_04545_));
 sky130_fd_sc_hd__a22o_1 _09936_ (.A1(\reg_module.gprf[303] ),
    .A2(net353),
    .B1(_04545_),
    .B2(net543),
    .X(_04546_));
 sky130_fd_sc_hd__and2_1 _09937_ (.A(net1154),
    .B(_04546_),
    .X(_00405_));
 sky130_fd_sc_hd__nor2_1 _09938_ (.A(net698),
    .B(net504),
    .Y(_04547_));
 sky130_fd_sc_hd__a22o_1 _09939_ (.A1(\reg_module.gprf[304] ),
    .A2(net354),
    .B1(_04547_),
    .B2(net559),
    .X(_04548_));
 sky130_fd_sc_hd__and2_1 _09940_ (.A(net1202),
    .B(_04548_),
    .X(_00406_));
 sky130_fd_sc_hd__nor2_1 _09941_ (.A(net697),
    .B(net503),
    .Y(_04549_));
 sky130_fd_sc_hd__a22o_1 _09942_ (.A1(\reg_module.gprf[305] ),
    .A2(net353),
    .B1(_04549_),
    .B2(net538),
    .X(_04550_));
 sky130_fd_sc_hd__and2_1 _09943_ (.A(net1140),
    .B(_04550_),
    .X(_00407_));
 sky130_fd_sc_hd__nor2_1 _09944_ (.A(net700),
    .B(net503),
    .Y(_04551_));
 sky130_fd_sc_hd__a22o_1 _09945_ (.A1(\reg_module.gprf[306] ),
    .A2(net353),
    .B1(_04551_),
    .B2(net538),
    .X(_04552_));
 sky130_fd_sc_hd__and2_1 _09946_ (.A(net1139),
    .B(_04552_),
    .X(_00408_));
 sky130_fd_sc_hd__nor2_1 _09947_ (.A(net699),
    .B(net503),
    .Y(_04553_));
 sky130_fd_sc_hd__a22o_1 _09948_ (.A1(\reg_module.gprf[307] ),
    .A2(net353),
    .B1(_04553_),
    .B2(net546),
    .X(_04554_));
 sky130_fd_sc_hd__and2_1 _09949_ (.A(net1159),
    .B(_04554_),
    .X(_00409_));
 sky130_fd_sc_hd__nor2_1 _09950_ (.A(net702),
    .B(net501),
    .Y(_04555_));
 sky130_fd_sc_hd__a22o_1 _09951_ (.A1(\reg_module.gprf[308] ),
    .A2(net352),
    .B1(_04555_),
    .B2(net526),
    .X(_04556_));
 sky130_fd_sc_hd__and2_1 _09952_ (.A(net1113),
    .B(_04556_),
    .X(_00410_));
 sky130_fd_sc_hd__nor2_1 _09953_ (.A(net701),
    .B(net504),
    .Y(_04557_));
 sky130_fd_sc_hd__a22o_1 _09954_ (.A1(\reg_module.gprf[309] ),
    .A2(net354),
    .B1(_04557_),
    .B2(net561),
    .X(_04558_));
 sky130_fd_sc_hd__and2_1 _09955_ (.A(net1207),
    .B(_04558_),
    .X(_00411_));
 sky130_fd_sc_hd__nor2_1 _09956_ (.A(net704),
    .B(net504),
    .Y(_04559_));
 sky130_fd_sc_hd__a22o_1 _09957_ (.A1(\reg_module.gprf[310] ),
    .A2(net354),
    .B1(_04559_),
    .B2(net557),
    .X(_04560_));
 sky130_fd_sc_hd__and2_1 _09958_ (.A(net1196),
    .B(_04560_),
    .X(_00412_));
 sky130_fd_sc_hd__nor2_1 _09959_ (.A(net703),
    .B(net504),
    .Y(_04561_));
 sky130_fd_sc_hd__a22o_1 _09960_ (.A1(\reg_module.gprf[311] ),
    .A2(net353),
    .B1(_04561_),
    .B2(net547),
    .X(_04562_));
 sky130_fd_sc_hd__and2_1 _09961_ (.A(net1165),
    .B(_04562_),
    .X(_00413_));
 sky130_fd_sc_hd__nor2_1 _09962_ (.A(net705),
    .B(net503),
    .Y(_04563_));
 sky130_fd_sc_hd__a22o_1 _09963_ (.A1(\reg_module.gprf[312] ),
    .A2(net353),
    .B1(_04563_),
    .B2(net553),
    .X(_04564_));
 sky130_fd_sc_hd__and2_1 _09964_ (.A(net1180),
    .B(_04564_),
    .X(_00414_));
 sky130_fd_sc_hd__nor2_1 _09965_ (.A(net706),
    .B(net503),
    .Y(_04565_));
 sky130_fd_sc_hd__a22o_1 _09966_ (.A1(\reg_module.gprf[313] ),
    .A2(net353),
    .B1(_04565_),
    .B2(net550),
    .X(_04566_));
 sky130_fd_sc_hd__and2_1 _09967_ (.A(net1172),
    .B(_04566_),
    .X(_00415_));
 sky130_fd_sc_hd__nor2_1 _09968_ (.A(net708),
    .B(net503),
    .Y(_04567_));
 sky130_fd_sc_hd__a22o_1 _09969_ (.A1(\reg_module.gprf[314] ),
    .A2(net353),
    .B1(_04567_),
    .B2(net546),
    .X(_04568_));
 sky130_fd_sc_hd__and2_1 _09970_ (.A(net1162),
    .B(_04568_),
    .X(_00416_));
 sky130_fd_sc_hd__nor2_1 _09971_ (.A(net707),
    .B(net503),
    .Y(_04569_));
 sky130_fd_sc_hd__a22o_1 _09972_ (.A1(\reg_module.gprf[315] ),
    .A2(net354),
    .B1(_04569_),
    .B2(net540),
    .X(_04570_));
 sky130_fd_sc_hd__and2_1 _09973_ (.A(net1146),
    .B(_04570_),
    .X(_00417_));
 sky130_fd_sc_hd__nor2_1 _09974_ (.A(net710),
    .B(net504),
    .Y(_04571_));
 sky130_fd_sc_hd__a22o_1 _09975_ (.A1(\reg_module.gprf[316] ),
    .A2(net354),
    .B1(_04571_),
    .B2(net549),
    .X(_04572_));
 sky130_fd_sc_hd__and2_1 _09976_ (.A(net1170),
    .B(_04572_),
    .X(_00418_));
 sky130_fd_sc_hd__nor2_1 _09977_ (.A(net709),
    .B(net503),
    .Y(_04573_));
 sky130_fd_sc_hd__a22o_1 _09978_ (.A1(\reg_module.gprf[317] ),
    .A2(net354),
    .B1(_04573_),
    .B2(net551),
    .X(_04574_));
 sky130_fd_sc_hd__and2_1 _09979_ (.A(net1178),
    .B(_04574_),
    .X(_00419_));
 sky130_fd_sc_hd__nor2_1 _09980_ (.A(net711),
    .B(net504),
    .Y(_04575_));
 sky130_fd_sc_hd__a22o_1 _09981_ (.A1(\reg_module.gprf[318] ),
    .A2(net354),
    .B1(_04575_),
    .B2(net558),
    .X(_04576_));
 sky130_fd_sc_hd__and2_1 _09982_ (.A(net1192),
    .B(_04576_),
    .X(_00420_));
 sky130_fd_sc_hd__nor2_1 _09983_ (.A(net574),
    .B(net504),
    .Y(_04577_));
 sky130_fd_sc_hd__a22o_1 _09984_ (.A1(\reg_module.gprf[319] ),
    .A2(net354),
    .B1(_04577_),
    .B2(net562),
    .X(_04578_));
 sky130_fd_sc_hd__and2_1 _09985_ (.A(net1205),
    .B(_04578_),
    .X(_00421_));
 sky130_fd_sc_hd__nand2b_4 _09986_ (.A_N(net965),
    .B(net748),
    .Y(_04579_));
 sky130_fd_sc_hd__or2_4 _09987_ (.A(_04175_),
    .B(net640),
    .X(_04580_));
 sky130_fd_sc_hd__nor2_1 _09988_ (.A(_02685_),
    .B(net640),
    .Y(_04581_));
 sky130_fd_sc_hd__a22o_1 _09989_ (.A1(\reg_module.gprf[320] ),
    .A2(net349),
    .B1(_04581_),
    .B2(net532),
    .X(_04582_));
 sky130_fd_sc_hd__and2_1 _09990_ (.A(net1124),
    .B(_04582_),
    .X(_00422_));
 sky130_fd_sc_hd__nor2_1 _09991_ (.A(net721),
    .B(net640),
    .Y(_04583_));
 sky130_fd_sc_hd__a22o_1 _09992_ (.A1(\reg_module.gprf[321] ),
    .A2(net349),
    .B1(_04583_),
    .B2(net533),
    .X(_04584_));
 sky130_fd_sc_hd__and2_1 _09993_ (.A(net1129),
    .B(_04584_),
    .X(_00423_));
 sky130_fd_sc_hd__nor2_1 _09994_ (.A(net713),
    .B(net639),
    .Y(_04585_));
 sky130_fd_sc_hd__a22o_1 _09995_ (.A1(\reg_module.gprf[322] ),
    .A2(net348),
    .B1(_04585_),
    .B2(net525),
    .X(_04586_));
 sky130_fd_sc_hd__and2_1 _09996_ (.A(net1110),
    .B(_04586_),
    .X(_00424_));
 sky130_fd_sc_hd__nor2_1 _09997_ (.A(net712),
    .B(net639),
    .Y(_04587_));
 sky130_fd_sc_hd__a22o_1 _09998_ (.A1(\reg_module.gprf[323] ),
    .A2(net348),
    .B1(_04587_),
    .B2(net515),
    .X(_04588_));
 sky130_fd_sc_hd__and2_1 _09999_ (.A(net1088),
    .B(_04588_),
    .X(_00425_));
 sky130_fd_sc_hd__nor2_1 _10000_ (.A(net723),
    .B(net640),
    .Y(_04589_));
 sky130_fd_sc_hd__a22o_1 _10001_ (.A1(\reg_module.gprf[324] ),
    .A2(net349),
    .B1(_04589_),
    .B2(net533),
    .X(_04590_));
 sky130_fd_sc_hd__and2_1 _10002_ (.A(net1127),
    .B(_04590_),
    .X(_00426_));
 sky130_fd_sc_hd__nor2_1 _10003_ (.A(net722),
    .B(net640),
    .Y(_04591_));
 sky130_fd_sc_hd__a22o_1 _10004_ (.A1(\reg_module.gprf[325] ),
    .A2(net349),
    .B1(_04591_),
    .B2(net529),
    .X(_04592_));
 sky130_fd_sc_hd__and2_1 _10005_ (.A(net1118),
    .B(_04592_),
    .X(_00427_));
 sky130_fd_sc_hd__nor2_1 _10006_ (.A(net725),
    .B(net639),
    .Y(_04593_));
 sky130_fd_sc_hd__a22o_1 _10007_ (.A1(\reg_module.gprf[326] ),
    .A2(net348),
    .B1(_04593_),
    .B2(net509),
    .X(_04594_));
 sky130_fd_sc_hd__and2_1 _10008_ (.A(net1071),
    .B(_04594_),
    .X(_00428_));
 sky130_fd_sc_hd__nor2_1 _10009_ (.A(net724),
    .B(net639),
    .Y(_04595_));
 sky130_fd_sc_hd__a22o_1 _10010_ (.A1(\reg_module.gprf[327] ),
    .A2(net348),
    .B1(_04595_),
    .B2(net514),
    .X(_04596_));
 sky130_fd_sc_hd__and2_1 _10011_ (.A(net1084),
    .B(_04596_),
    .X(_00429_));
 sky130_fd_sc_hd__nor2_1 _10012_ (.A(net689),
    .B(net640),
    .Y(_04597_));
 sky130_fd_sc_hd__a22o_1 _10013_ (.A1(\reg_module.gprf[328] ),
    .A2(net349),
    .B1(_04597_),
    .B2(net530),
    .X(_04598_));
 sky130_fd_sc_hd__and2_1 _10014_ (.A(net1121),
    .B(_04598_),
    .X(_00430_));
 sky130_fd_sc_hd__nor2_1 _10015_ (.A(net690),
    .B(net639),
    .Y(_04599_));
 sky130_fd_sc_hd__a22o_1 _10016_ (.A1(\reg_module.gprf[329] ),
    .A2(net348),
    .B1(_04599_),
    .B2(net518),
    .X(_04600_));
 sky130_fd_sc_hd__and2_1 _10017_ (.A(net1094),
    .B(_04600_),
    .X(_00431_));
 sky130_fd_sc_hd__nor2_1 _10018_ (.A(net692),
    .B(net639),
    .Y(_04601_));
 sky130_fd_sc_hd__a22o_1 _10019_ (.A1(\reg_module.gprf[330] ),
    .A2(net348),
    .B1(_04601_),
    .B2(net511),
    .X(_04602_));
 sky130_fd_sc_hd__and2_1 _10020_ (.A(net1074),
    .B(_04602_),
    .X(_00432_));
 sky130_fd_sc_hd__nor2_1 _10021_ (.A(net691),
    .B(net639),
    .Y(_04603_));
 sky130_fd_sc_hd__a22o_1 _10022_ (.A1(\reg_module.gprf[331] ),
    .A2(net348),
    .B1(_04603_),
    .B2(net520),
    .X(_04604_));
 sky130_fd_sc_hd__and2_1 _10023_ (.A(net1099),
    .B(_04604_),
    .X(_00433_));
 sky130_fd_sc_hd__nor2_1 _10024_ (.A(net693),
    .B(net641),
    .Y(_04605_));
 sky130_fd_sc_hd__a22o_1 _10025_ (.A1(\reg_module.gprf[332] ),
    .A2(net350),
    .B1(_04605_),
    .B2(net539),
    .X(_04606_));
 sky130_fd_sc_hd__and2_1 _10026_ (.A(net1143),
    .B(_04606_),
    .X(_00434_));
 sky130_fd_sc_hd__nor2_1 _10027_ (.A(net694),
    .B(net639),
    .Y(_04607_));
 sky130_fd_sc_hd__a22o_1 _10028_ (.A1(\reg_module.gprf[333] ),
    .A2(net348),
    .B1(_04607_),
    .B2(net524),
    .X(_04608_));
 sky130_fd_sc_hd__and2_1 _10029_ (.A(net1106),
    .B(_04608_),
    .X(_00435_));
 sky130_fd_sc_hd__nor2_1 _10030_ (.A(_02969_),
    .B(net639),
    .Y(_04609_));
 sky130_fd_sc_hd__a22o_1 _10031_ (.A1(\reg_module.gprf[334] ),
    .A2(net348),
    .B1(_04609_),
    .B2(net544),
    .X(_04610_));
 sky130_fd_sc_hd__and2_1 _10032_ (.A(net1155),
    .B(_04610_),
    .X(_00436_));
 sky130_fd_sc_hd__nor2_1 _10033_ (.A(net695),
    .B(net641),
    .Y(_04611_));
 sky130_fd_sc_hd__a22o_1 _10034_ (.A1(\reg_module.gprf[335] ),
    .A2(net350),
    .B1(_04611_),
    .B2(net543),
    .X(_04612_));
 sky130_fd_sc_hd__and2_1 _10035_ (.A(net1153),
    .B(_04612_),
    .X(_00437_));
 sky130_fd_sc_hd__nor2_1 _10036_ (.A(net698),
    .B(net642),
    .Y(_04613_));
 sky130_fd_sc_hd__a22o_1 _10037_ (.A1(\reg_module.gprf[336] ),
    .A2(net351),
    .B1(_04613_),
    .B2(net559),
    .X(_04614_));
 sky130_fd_sc_hd__and2_1 _10038_ (.A(net1201),
    .B(_04614_),
    .X(_00438_));
 sky130_fd_sc_hd__nor2_1 _10039_ (.A(net697),
    .B(net641),
    .Y(_04615_));
 sky130_fd_sc_hd__a22o_1 _10040_ (.A1(\reg_module.gprf[337] ),
    .A2(net350),
    .B1(_04615_),
    .B2(net539),
    .X(_04616_));
 sky130_fd_sc_hd__and2_1 _10041_ (.A(net1140),
    .B(_04616_),
    .X(_00439_));
 sky130_fd_sc_hd__nor2_1 _10042_ (.A(net700),
    .B(net641),
    .Y(_04617_));
 sky130_fd_sc_hd__a22o_1 _10043_ (.A1(\reg_module.gprf[338] ),
    .A2(net350),
    .B1(_04617_),
    .B2(net538),
    .X(_04618_));
 sky130_fd_sc_hd__and2_1 _10044_ (.A(net1139),
    .B(_04618_),
    .X(_00440_));
 sky130_fd_sc_hd__nor2_1 _10045_ (.A(net699),
    .B(net641),
    .Y(_04619_));
 sky130_fd_sc_hd__a22o_1 _10046_ (.A1(\reg_module.gprf[339] ),
    .A2(net350),
    .B1(_04619_),
    .B2(net546),
    .X(_04620_));
 sky130_fd_sc_hd__and2_1 _10047_ (.A(net1159),
    .B(_04620_),
    .X(_00441_));
 sky130_fd_sc_hd__nor2_1 _10048_ (.A(net702),
    .B(net639),
    .Y(_04621_));
 sky130_fd_sc_hd__a22o_1 _10049_ (.A1(\reg_module.gprf[340] ),
    .A2(net348),
    .B1(_04621_),
    .B2(net527),
    .X(_04622_));
 sky130_fd_sc_hd__and2_1 _10050_ (.A(net1114),
    .B(_04622_),
    .X(_00442_));
 sky130_fd_sc_hd__nor2_1 _10051_ (.A(net701),
    .B(net642),
    .Y(_04623_));
 sky130_fd_sc_hd__a22o_1 _10052_ (.A1(\reg_module.gprf[341] ),
    .A2(net351),
    .B1(_04623_),
    .B2(net562),
    .X(_04624_));
 sky130_fd_sc_hd__and2_1 _10053_ (.A(net1208),
    .B(_04624_),
    .X(_00443_));
 sky130_fd_sc_hd__nor2_1 _10054_ (.A(net704),
    .B(net642),
    .Y(_04625_));
 sky130_fd_sc_hd__a22o_1 _10055_ (.A1(\reg_module.gprf[342] ),
    .A2(net351),
    .B1(_04625_),
    .B2(net557),
    .X(_04626_));
 sky130_fd_sc_hd__and2_1 _10056_ (.A(net1193),
    .B(_04626_),
    .X(_00444_));
 sky130_fd_sc_hd__nor2_1 _10057_ (.A(net703),
    .B(net642),
    .Y(_04627_));
 sky130_fd_sc_hd__a22o_1 _10058_ (.A1(\reg_module.gprf[343] ),
    .A2(net351),
    .B1(_04627_),
    .B2(net547),
    .X(_04628_));
 sky130_fd_sc_hd__and2_1 _10059_ (.A(net1165),
    .B(_04628_),
    .X(_00445_));
 sky130_fd_sc_hd__nor2_1 _10060_ (.A(net705),
    .B(net641),
    .Y(_04629_));
 sky130_fd_sc_hd__a22o_1 _10061_ (.A1(\reg_module.gprf[344] ),
    .A2(net350),
    .B1(_04629_),
    .B2(net552),
    .X(_04630_));
 sky130_fd_sc_hd__and2_1 _10062_ (.A(net1180),
    .B(_04630_),
    .X(_00446_));
 sky130_fd_sc_hd__nor2_1 _10063_ (.A(net706),
    .B(net641),
    .Y(_04631_));
 sky130_fd_sc_hd__a22o_1 _10064_ (.A1(\reg_module.gprf[345] ),
    .A2(net350),
    .B1(_04631_),
    .B2(net553),
    .X(_04632_));
 sky130_fd_sc_hd__and2_1 _10065_ (.A(net1172),
    .B(_04632_),
    .X(_00447_));
 sky130_fd_sc_hd__nor2_1 _10066_ (.A(net708),
    .B(net641),
    .Y(_04633_));
 sky130_fd_sc_hd__a22o_1 _10067_ (.A1(\reg_module.gprf[346] ),
    .A2(net350),
    .B1(_04633_),
    .B2(net546),
    .X(_04634_));
 sky130_fd_sc_hd__and2_1 _10068_ (.A(net1159),
    .B(_04634_),
    .X(_00448_));
 sky130_fd_sc_hd__nor2_1 _10069_ (.A(net707),
    .B(net642),
    .Y(_04635_));
 sky130_fd_sc_hd__a22o_1 _10070_ (.A1(\reg_module.gprf[347] ),
    .A2(net350),
    .B1(_04635_),
    .B2(net547),
    .X(_04636_));
 sky130_fd_sc_hd__and2_1 _10071_ (.A(net1164),
    .B(_04636_),
    .X(_00449_));
 sky130_fd_sc_hd__nor2_1 _10072_ (.A(net710),
    .B(net641),
    .Y(_04637_));
 sky130_fd_sc_hd__a22o_1 _10073_ (.A1(\reg_module.gprf[348] ),
    .A2(net351),
    .B1(_04637_),
    .B2(net549),
    .X(_04638_));
 sky130_fd_sc_hd__and2_1 _10074_ (.A(net1170),
    .B(_04638_),
    .X(_00450_));
 sky130_fd_sc_hd__nor2_1 _10075_ (.A(net709),
    .B(net641),
    .Y(_04639_));
 sky130_fd_sc_hd__a22o_1 _10076_ (.A1(\reg_module.gprf[349] ),
    .A2(net350),
    .B1(_04639_),
    .B2(net551),
    .X(_04640_));
 sky130_fd_sc_hd__and2_1 _10077_ (.A(net1178),
    .B(_04640_),
    .X(_00451_));
 sky130_fd_sc_hd__nor2_1 _10078_ (.A(net711),
    .B(net642),
    .Y(_04641_));
 sky130_fd_sc_hd__a22o_1 _10079_ (.A1(\reg_module.gprf[350] ),
    .A2(net351),
    .B1(_04641_),
    .B2(net558),
    .X(_04642_));
 sky130_fd_sc_hd__and2_1 _10080_ (.A(net1193),
    .B(_04642_),
    .X(_00452_));
 sky130_fd_sc_hd__nor2_1 _10081_ (.A(net574),
    .B(net642),
    .Y(_04643_));
 sky130_fd_sc_hd__a22o_1 _10082_ (.A1(\reg_module.gprf[351] ),
    .A2(net351),
    .B1(_04643_),
    .B2(net560),
    .X(_04644_));
 sky130_fd_sc_hd__and2_1 _10083_ (.A(net1205),
    .B(_04644_),
    .X(_00453_));
 sky130_fd_sc_hd__or4_4 _10084_ (.A(\rReg_d2[0] ),
    .B(net970),
    .C(_01214_),
    .D(net967),
    .X(_04645_));
 sky130_fd_sc_hd__or2_1 _10085_ (.A(_04175_),
    .B(net636),
    .X(_04646_));
 sky130_fd_sc_hd__nor2_1 _10086_ (.A(_02685_),
    .B(net636),
    .Y(_04647_));
 sky130_fd_sc_hd__a22o_1 _10087_ (.A1(\reg_module.gprf[352] ),
    .A2(net347),
    .B1(_04647_),
    .B2(net532),
    .X(_04648_));
 sky130_fd_sc_hd__and2_1 _10088_ (.A(net1124),
    .B(_04648_),
    .X(_00454_));
 sky130_fd_sc_hd__nor2_1 _10089_ (.A(net721),
    .B(net636),
    .Y(_04649_));
 sky130_fd_sc_hd__a22o_1 _10090_ (.A1(\reg_module.gprf[353] ),
    .A2(net347),
    .B1(_04649_),
    .B2(net533),
    .X(_04650_));
 sky130_fd_sc_hd__and2_1 _10091_ (.A(net1129),
    .B(_04650_),
    .X(_00455_));
 sky130_fd_sc_hd__nor2_1 _10092_ (.A(net713),
    .B(net635),
    .Y(_04651_));
 sky130_fd_sc_hd__a22o_1 _10093_ (.A1(\reg_module.gprf[354] ),
    .A2(net344),
    .B1(_04651_),
    .B2(net524),
    .X(_04652_));
 sky130_fd_sc_hd__and2_1 _10094_ (.A(net1109),
    .B(_04652_),
    .X(_00456_));
 sky130_fd_sc_hd__nor2_1 _10095_ (.A(net712),
    .B(net635),
    .Y(_04653_));
 sky130_fd_sc_hd__a22o_1 _10096_ (.A1(\reg_module.gprf[355] ),
    .A2(net344),
    .B1(_04653_),
    .B2(net515),
    .X(_04654_));
 sky130_fd_sc_hd__and2_1 _10097_ (.A(net1088),
    .B(_04654_),
    .X(_00457_));
 sky130_fd_sc_hd__nor2_1 _10098_ (.A(net723),
    .B(net636),
    .Y(_04655_));
 sky130_fd_sc_hd__a22o_1 _10099_ (.A1(\reg_module.gprf[356] ),
    .A2(net347),
    .B1(_04655_),
    .B2(net533),
    .X(_04656_));
 sky130_fd_sc_hd__and2_1 _10100_ (.A(net1127),
    .B(_04656_),
    .X(_00458_));
 sky130_fd_sc_hd__nor2_1 _10101_ (.A(net722),
    .B(net636),
    .Y(_04657_));
 sky130_fd_sc_hd__a22o_1 _10102_ (.A1(\reg_module.gprf[357] ),
    .A2(net344),
    .B1(_04657_),
    .B2(net529),
    .X(_04658_));
 sky130_fd_sc_hd__and2_1 _10103_ (.A(net1118),
    .B(_04658_),
    .X(_00459_));
 sky130_fd_sc_hd__nor2_1 _10104_ (.A(net725),
    .B(net635),
    .Y(_04659_));
 sky130_fd_sc_hd__a22o_1 _10105_ (.A1(\reg_module.gprf[358] ),
    .A2(net344),
    .B1(_04659_),
    .B2(net509),
    .X(_04660_));
 sky130_fd_sc_hd__and2_1 _10106_ (.A(net1071),
    .B(_04660_),
    .X(_00460_));
 sky130_fd_sc_hd__nor2_1 _10107_ (.A(net724),
    .B(net635),
    .Y(_04661_));
 sky130_fd_sc_hd__a22o_1 _10108_ (.A1(\reg_module.gprf[359] ),
    .A2(net344),
    .B1(_04661_),
    .B2(net514),
    .X(_04662_));
 sky130_fd_sc_hd__and2_1 _10109_ (.A(net1084),
    .B(_04662_),
    .X(_00461_));
 sky130_fd_sc_hd__nor2_1 _10110_ (.A(net689),
    .B(net636),
    .Y(_04663_));
 sky130_fd_sc_hd__a22o_1 _10111_ (.A1(\reg_module.gprf[360] ),
    .A2(net347),
    .B1(_04663_),
    .B2(net535),
    .X(_04664_));
 sky130_fd_sc_hd__and2_1 _10112_ (.A(net1121),
    .B(_04664_),
    .X(_00462_));
 sky130_fd_sc_hd__nor2_1 _10113_ (.A(net690),
    .B(net635),
    .Y(_04665_));
 sky130_fd_sc_hd__a22o_1 _10114_ (.A1(\reg_module.gprf[361] ),
    .A2(net344),
    .B1(_04665_),
    .B2(net518),
    .X(_04666_));
 sky130_fd_sc_hd__and2_1 _10115_ (.A(net1094),
    .B(_04666_),
    .X(_00463_));
 sky130_fd_sc_hd__nor2_1 _10116_ (.A(net692),
    .B(net635),
    .Y(_04667_));
 sky130_fd_sc_hd__a22o_1 _10117_ (.A1(\reg_module.gprf[362] ),
    .A2(net344),
    .B1(_04667_),
    .B2(net511),
    .X(_04668_));
 sky130_fd_sc_hd__and2_1 _10118_ (.A(net1075),
    .B(_04668_),
    .X(_00464_));
 sky130_fd_sc_hd__nor2_1 _10119_ (.A(net691),
    .B(net635),
    .Y(_04669_));
 sky130_fd_sc_hd__a22o_1 _10120_ (.A1(\reg_module.gprf[363] ),
    .A2(net344),
    .B1(_04669_),
    .B2(net520),
    .X(_04670_));
 sky130_fd_sc_hd__and2_1 _10121_ (.A(net1099),
    .B(_04670_),
    .X(_00465_));
 sky130_fd_sc_hd__nor2_1 _10122_ (.A(net693),
    .B(net637),
    .Y(_04671_));
 sky130_fd_sc_hd__a22o_1 _10123_ (.A1(\reg_module.gprf[364] ),
    .A2(net345),
    .B1(_04671_),
    .B2(net539),
    .X(_04672_));
 sky130_fd_sc_hd__and2_1 _10124_ (.A(net1142),
    .B(_04672_),
    .X(_00466_));
 sky130_fd_sc_hd__nor2_1 _10125_ (.A(net694),
    .B(net635),
    .Y(_04673_));
 sky130_fd_sc_hd__a22o_1 _10126_ (.A1(\reg_module.gprf[365] ),
    .A2(net344),
    .B1(_04673_),
    .B2(net524),
    .X(_04674_));
 sky130_fd_sc_hd__and2_1 _10127_ (.A(net1106),
    .B(_04674_),
    .X(_00467_));
 sky130_fd_sc_hd__nor2_1 _10128_ (.A(_02969_),
    .B(net635),
    .Y(_04675_));
 sky130_fd_sc_hd__a22o_1 _10129_ (.A1(\reg_module.gprf[366] ),
    .A2(net345),
    .B1(_04675_),
    .B2(net544),
    .X(_04676_));
 sky130_fd_sc_hd__and2_1 _10130_ (.A(net1155),
    .B(_04676_),
    .X(_00468_));
 sky130_fd_sc_hd__nor2_1 _10131_ (.A(net695),
    .B(net637),
    .Y(_04677_));
 sky130_fd_sc_hd__a22o_1 _10132_ (.A1(\reg_module.gprf[367] ),
    .A2(net345),
    .B1(_04677_),
    .B2(net546),
    .X(_04678_));
 sky130_fd_sc_hd__and2_1 _10133_ (.A(net1158),
    .B(_04678_),
    .X(_00469_));
 sky130_fd_sc_hd__nor2_1 _10134_ (.A(net698),
    .B(net638),
    .Y(_04679_));
 sky130_fd_sc_hd__a22o_1 _10135_ (.A1(\reg_module.gprf[368] ),
    .A2(net346),
    .B1(_04679_),
    .B2(net559),
    .X(_04680_));
 sky130_fd_sc_hd__and2_1 _10136_ (.A(net1201),
    .B(_04680_),
    .X(_00470_));
 sky130_fd_sc_hd__nor2_1 _10137_ (.A(net697),
    .B(net637),
    .Y(_04681_));
 sky130_fd_sc_hd__a22o_1 _10138_ (.A1(\reg_module.gprf[369] ),
    .A2(net345),
    .B1(_04681_),
    .B2(net540),
    .X(_04682_));
 sky130_fd_sc_hd__and2_1 _10139_ (.A(net1145),
    .B(_04682_),
    .X(_00471_));
 sky130_fd_sc_hd__nor2_1 _10140_ (.A(net700),
    .B(net637),
    .Y(_04683_));
 sky130_fd_sc_hd__a22o_1 _10141_ (.A1(\reg_module.gprf[370] ),
    .A2(net345),
    .B1(_04683_),
    .B2(net538),
    .X(_04684_));
 sky130_fd_sc_hd__and2_1 _10142_ (.A(net1139),
    .B(_04684_),
    .X(_00472_));
 sky130_fd_sc_hd__nor2_1 _10143_ (.A(net699),
    .B(net637),
    .Y(_04685_));
 sky130_fd_sc_hd__a22o_1 _10144_ (.A1(\reg_module.gprf[371] ),
    .A2(net345),
    .B1(_04685_),
    .B2(net546),
    .X(_04686_));
 sky130_fd_sc_hd__and2_1 _10145_ (.A(net1159),
    .B(_04686_),
    .X(_00473_));
 sky130_fd_sc_hd__nor2_1 _10146_ (.A(net702),
    .B(net635),
    .Y(_04687_));
 sky130_fd_sc_hd__a22o_1 _10147_ (.A1(\reg_module.gprf[372] ),
    .A2(net344),
    .B1(_04687_),
    .B2(net526),
    .X(_04688_));
 sky130_fd_sc_hd__and2_1 _10148_ (.A(net1114),
    .B(_04688_),
    .X(_00474_));
 sky130_fd_sc_hd__nor2_1 _10149_ (.A(net701),
    .B(net638),
    .Y(_04689_));
 sky130_fd_sc_hd__a22o_1 _10150_ (.A1(\reg_module.gprf[373] ),
    .A2(net346),
    .B1(_04689_),
    .B2(net561),
    .X(_04690_));
 sky130_fd_sc_hd__and2_1 _10151_ (.A(net1208),
    .B(_04690_),
    .X(_00475_));
 sky130_fd_sc_hd__nor2_1 _10152_ (.A(net704),
    .B(net638),
    .Y(_04691_));
 sky130_fd_sc_hd__a22o_1 _10153_ (.A1(\reg_module.gprf[374] ),
    .A2(net346),
    .B1(_04691_),
    .B2(net564),
    .X(_04692_));
 sky130_fd_sc_hd__and2_1 _10154_ (.A(net1193),
    .B(_04692_),
    .X(_00476_));
 sky130_fd_sc_hd__nor2_1 _10155_ (.A(net703),
    .B(net638),
    .Y(_04693_));
 sky130_fd_sc_hd__a22o_1 _10156_ (.A1(\reg_module.gprf[375] ),
    .A2(net346),
    .B1(_04693_),
    .B2(net549),
    .X(_04694_));
 sky130_fd_sc_hd__and2_1 _10157_ (.A(net1165),
    .B(_04694_),
    .X(_00477_));
 sky130_fd_sc_hd__nor2_1 _10158_ (.A(net705),
    .B(net637),
    .Y(_04695_));
 sky130_fd_sc_hd__a22o_1 _10159_ (.A1(\reg_module.gprf[376] ),
    .A2(net345),
    .B1(_04695_),
    .B2(net553),
    .X(_04696_));
 sky130_fd_sc_hd__and2_1 _10160_ (.A(net1185),
    .B(_04696_),
    .X(_00478_));
 sky130_fd_sc_hd__nor2_1 _10161_ (.A(net706),
    .B(net637),
    .Y(_04697_));
 sky130_fd_sc_hd__a22o_1 _10162_ (.A1(\reg_module.gprf[377] ),
    .A2(net345),
    .B1(_04697_),
    .B2(net553),
    .X(_04698_));
 sky130_fd_sc_hd__and2_1 _10163_ (.A(net1172),
    .B(_04698_),
    .X(_00479_));
 sky130_fd_sc_hd__nor2_1 _10164_ (.A(net708),
    .B(net637),
    .Y(_04699_));
 sky130_fd_sc_hd__a22o_1 _10165_ (.A1(\reg_module.gprf[378] ),
    .A2(net345),
    .B1(_04699_),
    .B2(net546),
    .X(_04700_));
 sky130_fd_sc_hd__and2_1 _10166_ (.A(net1162),
    .B(_04700_),
    .X(_00480_));
 sky130_fd_sc_hd__nor2_1 _10167_ (.A(net707),
    .B(net637),
    .Y(_04701_));
 sky130_fd_sc_hd__a22o_1 _10168_ (.A1(\reg_module.gprf[379] ),
    .A2(net345),
    .B1(_04701_),
    .B2(net547),
    .X(_04702_));
 sky130_fd_sc_hd__and2_1 _10169_ (.A(net1164),
    .B(_04702_),
    .X(_00481_));
 sky130_fd_sc_hd__nor2_1 _10170_ (.A(net710),
    .B(net638),
    .Y(_04703_));
 sky130_fd_sc_hd__a22o_1 _10171_ (.A1(\reg_module.gprf[380] ),
    .A2(net346),
    .B1(_04703_),
    .B2(net549),
    .X(_04704_));
 sky130_fd_sc_hd__and2_1 _10172_ (.A(net1170),
    .B(_04704_),
    .X(_00482_));
 sky130_fd_sc_hd__nor2_1 _10173_ (.A(_02770_),
    .B(net637),
    .Y(_04705_));
 sky130_fd_sc_hd__a22o_1 _10174_ (.A1(\reg_module.gprf[381] ),
    .A2(net346),
    .B1(_04705_),
    .B2(net551),
    .X(_04706_));
 sky130_fd_sc_hd__and2_1 _10175_ (.A(net1178),
    .B(_04706_),
    .X(_00483_));
 sky130_fd_sc_hd__nor2_1 _10176_ (.A(net711),
    .B(net638),
    .Y(_04707_));
 sky130_fd_sc_hd__a22o_1 _10177_ (.A1(\reg_module.gprf[382] ),
    .A2(net346),
    .B1(_04707_),
    .B2(net554),
    .X(_04708_));
 sky130_fd_sc_hd__and2_1 _10178_ (.A(net1183),
    .B(_04708_),
    .X(_00484_));
 sky130_fd_sc_hd__nor2_1 _10179_ (.A(net574),
    .B(net638),
    .Y(_04709_));
 sky130_fd_sc_hd__a22o_1 _10180_ (.A1(\reg_module.gprf[383] ),
    .A2(net346),
    .B1(_04709_),
    .B2(net560),
    .X(_04710_));
 sky130_fd_sc_hd__and2_1 _10181_ (.A(net1205),
    .B(_04710_),
    .X(_00485_));
 sky130_fd_sc_hd__nand2b_4 _10182_ (.A_N(net965),
    .B(net658),
    .Y(_04711_));
 sky130_fd_sc_hd__or2_4 _10183_ (.A(_04175_),
    .B(net498),
    .X(_04712_));
 sky130_fd_sc_hd__nor2_1 _10184_ (.A(_02685_),
    .B(net498),
    .Y(_04713_));
 sky130_fd_sc_hd__a22o_1 _10185_ (.A1(\reg_module.gprf[384] ),
    .A2(net341),
    .B1(_04713_),
    .B2(net532),
    .X(_04714_));
 sky130_fd_sc_hd__and2_1 _10186_ (.A(net1089),
    .B(_04714_),
    .X(_00486_));
 sky130_fd_sc_hd__nor2_1 _10187_ (.A(net721),
    .B(net498),
    .Y(_04715_));
 sky130_fd_sc_hd__a22o_1 _10188_ (.A1(\reg_module.gprf[385] ),
    .A2(net341),
    .B1(_04715_),
    .B2(net536),
    .X(_04716_));
 sky130_fd_sc_hd__and2_1 _10189_ (.A(net1132),
    .B(_04716_),
    .X(_00487_));
 sky130_fd_sc_hd__nor2_1 _10190_ (.A(net713),
    .B(net497),
    .Y(_04717_));
 sky130_fd_sc_hd__a22o_1 _10191_ (.A1(\reg_module.gprf[386] ),
    .A2(net341),
    .B1(_04717_),
    .B2(net525),
    .X(_04718_));
 sky130_fd_sc_hd__and2_1 _10192_ (.A(net1110),
    .B(_04718_),
    .X(_00488_));
 sky130_fd_sc_hd__nor2_1 _10193_ (.A(net712),
    .B(net497),
    .Y(_04719_));
 sky130_fd_sc_hd__a22o_1 _10194_ (.A1(\reg_module.gprf[387] ),
    .A2(net340),
    .B1(_04719_),
    .B2(net516),
    .X(_04720_));
 sky130_fd_sc_hd__and2_1 _10195_ (.A(net1087),
    .B(_04720_),
    .X(_00489_));
 sky130_fd_sc_hd__nor2_1 _10196_ (.A(_02642_),
    .B(net498),
    .Y(_04721_));
 sky130_fd_sc_hd__a22o_1 _10197_ (.A1(\reg_module.gprf[388] ),
    .A2(net341),
    .B1(_04721_),
    .B2(net534),
    .X(_04722_));
 sky130_fd_sc_hd__and2_1 _10198_ (.A(net1130),
    .B(_04722_),
    .X(_00490_));
 sky130_fd_sc_hd__nor2_1 _10199_ (.A(net722),
    .B(net498),
    .Y(_04723_));
 sky130_fd_sc_hd__a22o_1 _10200_ (.A1(\reg_module.gprf[389] ),
    .A2(net341),
    .B1(_04723_),
    .B2(net531),
    .X(_04724_));
 sky130_fd_sc_hd__and2_1 _10201_ (.A(net1120),
    .B(_04724_),
    .X(_00491_));
 sky130_fd_sc_hd__nor2_1 _10202_ (.A(_02604_),
    .B(net497),
    .Y(_04725_));
 sky130_fd_sc_hd__a22o_1 _10203_ (.A1(\reg_module.gprf[390] ),
    .A2(net340),
    .B1(_04725_),
    .B2(net513),
    .X(_04726_));
 sky130_fd_sc_hd__and2_1 _10204_ (.A(net1081),
    .B(_04726_),
    .X(_00492_));
 sky130_fd_sc_hd__nor2_1 _10205_ (.A(net724),
    .B(net497),
    .Y(_04727_));
 sky130_fd_sc_hd__a22o_1 _10206_ (.A1(\reg_module.gprf[391] ),
    .A2(net340),
    .B1(_04727_),
    .B2(net514),
    .X(_04728_));
 sky130_fd_sc_hd__and2_1 _10207_ (.A(net1086),
    .B(_04728_),
    .X(_00493_));
 sky130_fd_sc_hd__nor2_1 _10208_ (.A(net689),
    .B(net498),
    .Y(_04729_));
 sky130_fd_sc_hd__a22o_1 _10209_ (.A1(\reg_module.gprf[392] ),
    .A2(net341),
    .B1(_04729_),
    .B2(net530),
    .X(_04730_));
 sky130_fd_sc_hd__and2_1 _10210_ (.A(net1122),
    .B(_04730_),
    .X(_00494_));
 sky130_fd_sc_hd__nor2_1 _10211_ (.A(_03061_),
    .B(net497),
    .Y(_04731_));
 sky130_fd_sc_hd__a22o_1 _10212_ (.A1(\reg_module.gprf[393] ),
    .A2(net340),
    .B1(_04731_),
    .B2(net511),
    .X(_04732_));
 sky130_fd_sc_hd__and2_1 _10213_ (.A(net1075),
    .B(_04732_),
    .X(_00495_));
 sky130_fd_sc_hd__nor2_1 _10214_ (.A(net692),
    .B(net497),
    .Y(_04733_));
 sky130_fd_sc_hd__a22o_1 _10215_ (.A1(\reg_module.gprf[394] ),
    .A2(net340),
    .B1(_04733_),
    .B2(net510),
    .X(_04734_));
 sky130_fd_sc_hd__and2_1 _10216_ (.A(net1073),
    .B(_04734_),
    .X(_00496_));
 sky130_fd_sc_hd__nor2_1 _10217_ (.A(net691),
    .B(net497),
    .Y(_04735_));
 sky130_fd_sc_hd__a22o_1 _10218_ (.A1(\reg_module.gprf[395] ),
    .A2(net340),
    .B1(_04735_),
    .B2(net519),
    .X(_04736_));
 sky130_fd_sc_hd__and2_1 _10219_ (.A(net1095),
    .B(_04736_),
    .X(_00497_));
 sky130_fd_sc_hd__nor2_1 _10220_ (.A(net693),
    .B(net499),
    .Y(_04737_));
 sky130_fd_sc_hd__a22o_1 _10221_ (.A1(\reg_module.gprf[396] ),
    .A2(net340),
    .B1(_04737_),
    .B2(net543),
    .X(_04738_));
 sky130_fd_sc_hd__and2_1 _10222_ (.A(net1152),
    .B(_04738_),
    .X(_00498_));
 sky130_fd_sc_hd__nor2_1 _10223_ (.A(net694),
    .B(net497),
    .Y(_04739_));
 sky130_fd_sc_hd__a22o_1 _10224_ (.A1(\reg_module.gprf[397] ),
    .A2(net340),
    .B1(_04739_),
    .B2(net523),
    .X(_04740_));
 sky130_fd_sc_hd__and2_1 _10225_ (.A(net1097),
    .B(_04740_),
    .X(_00499_));
 sky130_fd_sc_hd__nor2_1 _10226_ (.A(net696),
    .B(net498),
    .Y(_04741_));
 sky130_fd_sc_hd__a22o_1 _10227_ (.A1(\reg_module.gprf[398] ),
    .A2(net341),
    .B1(_04741_),
    .B2(net537),
    .X(_04742_));
 sky130_fd_sc_hd__and2_1 _10228_ (.A(net1135),
    .B(_04742_),
    .X(_00500_));
 sky130_fd_sc_hd__nor2_1 _10229_ (.A(_02984_),
    .B(net499),
    .Y(_04743_));
 sky130_fd_sc_hd__a22o_1 _10230_ (.A1(\reg_module.gprf[399] ),
    .A2(net342),
    .B1(_04743_),
    .B2(net544),
    .X(_04744_));
 sky130_fd_sc_hd__and2_1 _10231_ (.A(net1156),
    .B(_04744_),
    .X(_00501_));
 sky130_fd_sc_hd__nor2_1 _10232_ (.A(net698),
    .B(net500),
    .Y(_04745_));
 sky130_fd_sc_hd__a22o_1 _10233_ (.A1(\reg_module.gprf[400] ),
    .A2(net343),
    .B1(_04745_),
    .B2(net565),
    .X(_04746_));
 sky130_fd_sc_hd__and2_1 _10234_ (.A(net1189),
    .B(_04746_),
    .X(_00502_));
 sky130_fd_sc_hd__nor2_1 _10235_ (.A(net697),
    .B(net499),
    .Y(_04747_));
 sky130_fd_sc_hd__a22o_1 _10236_ (.A1(\reg_module.gprf[401] ),
    .A2(net342),
    .B1(_04747_),
    .B2(net539),
    .X(_04748_));
 sky130_fd_sc_hd__and2_1 _10237_ (.A(net1141),
    .B(_04748_),
    .X(_00503_));
 sky130_fd_sc_hd__nor2_1 _10238_ (.A(net700),
    .B(net497),
    .Y(_04749_));
 sky130_fd_sc_hd__a22o_1 _10239_ (.A1(\reg_module.gprf[402] ),
    .A2(net340),
    .B1(_04749_),
    .B2(net522),
    .X(_04750_));
 sky130_fd_sc_hd__and2_1 _10240_ (.A(net1100),
    .B(_04750_),
    .X(_00504_));
 sky130_fd_sc_hd__nor2_1 _10241_ (.A(net699),
    .B(net499),
    .Y(_04751_));
 sky130_fd_sc_hd__a22o_1 _10242_ (.A1(\reg_module.gprf[403] ),
    .A2(net342),
    .B1(_04751_),
    .B2(net546),
    .X(_04752_));
 sky130_fd_sc_hd__and2_1 _10243_ (.A(net1148),
    .B(_04752_),
    .X(_00505_));
 sky130_fd_sc_hd__nor2_1 _10244_ (.A(net702),
    .B(net497),
    .Y(_04753_));
 sky130_fd_sc_hd__a22o_1 _10245_ (.A1(\reg_module.gprf[404] ),
    .A2(net340),
    .B1(_04753_),
    .B2(net543),
    .X(_04754_));
 sky130_fd_sc_hd__and2_1 _10246_ (.A(net1152),
    .B(_04754_),
    .X(_00506_));
 sky130_fd_sc_hd__nor2_1 _10247_ (.A(net701),
    .B(net500),
    .Y(_04755_));
 sky130_fd_sc_hd__a22o_1 _10248_ (.A1(\reg_module.gprf[405] ),
    .A2(net343),
    .B1(_04755_),
    .B2(net559),
    .X(_04756_));
 sky130_fd_sc_hd__and2_1 _10249_ (.A(net1201),
    .B(_04756_),
    .X(_00507_));
 sky130_fd_sc_hd__nor2_1 _10250_ (.A(net704),
    .B(net500),
    .Y(_04757_));
 sky130_fd_sc_hd__a22o_1 _10251_ (.A1(\reg_module.gprf[406] ),
    .A2(net343),
    .B1(_04757_),
    .B2(net560),
    .X(_04758_));
 sky130_fd_sc_hd__and2_1 _10252_ (.A(net1196),
    .B(_04758_),
    .X(_00508_));
 sky130_fd_sc_hd__nor2_1 _10253_ (.A(net703),
    .B(net499),
    .Y(_04759_));
 sky130_fd_sc_hd__a22o_1 _10254_ (.A1(\reg_module.gprf[407] ),
    .A2(net342),
    .B1(_04759_),
    .B2(net547),
    .X(_04760_));
 sky130_fd_sc_hd__and2_1 _10255_ (.A(net1165),
    .B(_04760_),
    .X(_00509_));
 sky130_fd_sc_hd__nor2_1 _10256_ (.A(net705),
    .B(net499),
    .Y(_04761_));
 sky130_fd_sc_hd__a22o_1 _10257_ (.A1(\reg_module.gprf[408] ),
    .A2(net342),
    .B1(_04761_),
    .B2(net554),
    .X(_04762_));
 sky130_fd_sc_hd__and2_1 _10258_ (.A(net1182),
    .B(_04762_),
    .X(_00510_));
 sky130_fd_sc_hd__nor2_1 _10259_ (.A(net706),
    .B(net499),
    .Y(_04763_));
 sky130_fd_sc_hd__a22o_1 _10260_ (.A1(\reg_module.gprf[409] ),
    .A2(net342),
    .B1(_04763_),
    .B2(net552),
    .X(_04764_));
 sky130_fd_sc_hd__and2_1 _10261_ (.A(net1185),
    .B(_04764_),
    .X(_00511_));
 sky130_fd_sc_hd__nor2_1 _10262_ (.A(net708),
    .B(net499),
    .Y(_04765_));
 sky130_fd_sc_hd__a22o_1 _10263_ (.A1(\reg_module.gprf[410] ),
    .A2(net342),
    .B1(_04765_),
    .B2(net545),
    .X(_04766_));
 sky130_fd_sc_hd__and2_1 _10264_ (.A(net1162),
    .B(_04766_),
    .X(_00512_));
 sky130_fd_sc_hd__nor2_1 _10265_ (.A(net707),
    .B(net499),
    .Y(_04767_));
 sky130_fd_sc_hd__a22o_1 _10266_ (.A1(\reg_module.gprf[411] ),
    .A2(net342),
    .B1(_04767_),
    .B2(net540),
    .X(_04768_));
 sky130_fd_sc_hd__and2_1 _10267_ (.A(net1146),
    .B(_04768_),
    .X(_00513_));
 sky130_fd_sc_hd__nor2_1 _10268_ (.A(_02756_),
    .B(net499),
    .Y(_04769_));
 sky130_fd_sc_hd__a22o_1 _10269_ (.A1(\reg_module.gprf[412] ),
    .A2(net342),
    .B1(_04769_),
    .B2(net549),
    .X(_04770_));
 sky130_fd_sc_hd__and2_1 _10270_ (.A(net1172),
    .B(_04770_),
    .X(_00514_));
 sky130_fd_sc_hd__nor2_1 _10271_ (.A(net709),
    .B(net500),
    .Y(_04771_));
 sky130_fd_sc_hd__a22o_1 _10272_ (.A1(\reg_module.gprf[413] ),
    .A2(net342),
    .B1(_04771_),
    .B2(net555),
    .X(_04772_));
 sky130_fd_sc_hd__and2_1 _10273_ (.A(net1175),
    .B(_04772_),
    .X(_00515_));
 sky130_fd_sc_hd__nor2_1 _10274_ (.A(net711),
    .B(net500),
    .Y(_04773_));
 sky130_fd_sc_hd__a22o_1 _10275_ (.A1(\reg_module.gprf[414] ),
    .A2(net343),
    .B1(_04773_),
    .B2(net558),
    .X(_04774_));
 sky130_fd_sc_hd__and2_1 _10276_ (.A(net1193),
    .B(_04774_),
    .X(_00516_));
 sky130_fd_sc_hd__nor2_1 _10277_ (.A(net574),
    .B(net500),
    .Y(_04775_));
 sky130_fd_sc_hd__a22o_1 _10278_ (.A1(\reg_module.gprf[415] ),
    .A2(net343),
    .B1(_04775_),
    .B2(net562),
    .X(_04776_));
 sky130_fd_sc_hd__and2_1 _10279_ (.A(net1205),
    .B(_04776_),
    .X(_00517_));
 sky130_fd_sc_hd__nand2b_4 _10280_ (.A_N(net965),
    .B(net650),
    .Y(_04777_));
 sky130_fd_sc_hd__or2_4 _10281_ (.A(_04175_),
    .B(net494),
    .X(_04778_));
 sky130_fd_sc_hd__nor2_1 _10282_ (.A(_02685_),
    .B(net494),
    .Y(_04779_));
 sky130_fd_sc_hd__a22o_1 _10283_ (.A1(\reg_module.gprf[416] ),
    .A2(net337),
    .B1(_04779_),
    .B2(net532),
    .X(_04780_));
 sky130_fd_sc_hd__and2_1 _10284_ (.A(net1091),
    .B(_04780_),
    .X(_00518_));
 sky130_fd_sc_hd__nor2_1 _10285_ (.A(net721),
    .B(net494),
    .Y(_04781_));
 sky130_fd_sc_hd__a22o_1 _10286_ (.A1(\reg_module.gprf[417] ),
    .A2(net337),
    .B1(_04781_),
    .B2(net536),
    .X(_04782_));
 sky130_fd_sc_hd__and2_1 _10287_ (.A(net1132),
    .B(_04782_),
    .X(_00519_));
 sky130_fd_sc_hd__nor2_1 _10288_ (.A(net713),
    .B(net494),
    .Y(_04783_));
 sky130_fd_sc_hd__a22o_1 _10289_ (.A1(\reg_module.gprf[418] ),
    .A2(net337),
    .B1(_04783_),
    .B2(net525),
    .X(_04784_));
 sky130_fd_sc_hd__and2_1 _10290_ (.A(net1110),
    .B(_04784_),
    .X(_00520_));
 sky130_fd_sc_hd__nor2_1 _10291_ (.A(net712),
    .B(net493),
    .Y(_04785_));
 sky130_fd_sc_hd__a22o_1 _10292_ (.A1(\reg_module.gprf[419] ),
    .A2(net336),
    .B1(_04785_),
    .B2(net516),
    .X(_04786_));
 sky130_fd_sc_hd__and2_1 _10293_ (.A(net1087),
    .B(_04786_),
    .X(_00521_));
 sky130_fd_sc_hd__nor2_1 _10294_ (.A(net723),
    .B(net494),
    .Y(_04787_));
 sky130_fd_sc_hd__a22o_1 _10295_ (.A1(\reg_module.gprf[420] ),
    .A2(net337),
    .B1(_04787_),
    .B2(net533),
    .X(_04788_));
 sky130_fd_sc_hd__and2_1 _10296_ (.A(net1130),
    .B(_04788_),
    .X(_00522_));
 sky130_fd_sc_hd__nor2_1 _10297_ (.A(net722),
    .B(net494),
    .Y(_04789_));
 sky130_fd_sc_hd__a22o_1 _10298_ (.A1(\reg_module.gprf[421] ),
    .A2(net337),
    .B1(_04789_),
    .B2(net529),
    .X(_04790_));
 sky130_fd_sc_hd__and2_1 _10299_ (.A(net1118),
    .B(_04790_),
    .X(_00523_));
 sky130_fd_sc_hd__nor2_1 _10300_ (.A(net725),
    .B(net493),
    .Y(_04791_));
 sky130_fd_sc_hd__a22o_1 _10301_ (.A1(\reg_module.gprf[422] ),
    .A2(net336),
    .B1(_04791_),
    .B2(net513),
    .X(_04792_));
 sky130_fd_sc_hd__and2_1 _10302_ (.A(net1081),
    .B(_04792_),
    .X(_00524_));
 sky130_fd_sc_hd__nor2_1 _10303_ (.A(_02623_),
    .B(net493),
    .Y(_04793_));
 sky130_fd_sc_hd__a22o_1 _10304_ (.A1(\reg_module.gprf[423] ),
    .A2(net336),
    .B1(_04793_),
    .B2(net514),
    .X(_04794_));
 sky130_fd_sc_hd__and2_1 _10305_ (.A(net1086),
    .B(_04794_),
    .X(_00525_));
 sky130_fd_sc_hd__nor2_1 _10306_ (.A(net689),
    .B(net494),
    .Y(_04795_));
 sky130_fd_sc_hd__a22o_1 _10307_ (.A1(\reg_module.gprf[424] ),
    .A2(net337),
    .B1(_04795_),
    .B2(net530),
    .X(_04796_));
 sky130_fd_sc_hd__and2_1 _10308_ (.A(net1122),
    .B(_04796_),
    .X(_00526_));
 sky130_fd_sc_hd__nor2_1 _10309_ (.A(net690),
    .B(net493),
    .Y(_04797_));
 sky130_fd_sc_hd__a22o_1 _10310_ (.A1(\reg_module.gprf[425] ),
    .A2(net336),
    .B1(_04797_),
    .B2(net511),
    .X(_04798_));
 sky130_fd_sc_hd__and2_1 _10311_ (.A(net1076),
    .B(_04798_),
    .X(_00527_));
 sky130_fd_sc_hd__nor2_1 _10312_ (.A(net692),
    .B(net493),
    .Y(_04799_));
 sky130_fd_sc_hd__a22o_1 _10313_ (.A1(\reg_module.gprf[426] ),
    .A2(net336),
    .B1(_04799_),
    .B2(net510),
    .X(_04800_));
 sky130_fd_sc_hd__and2_1 _10314_ (.A(net1074),
    .B(_04800_),
    .X(_00528_));
 sky130_fd_sc_hd__nor2_1 _10315_ (.A(net691),
    .B(net493),
    .Y(_04801_));
 sky130_fd_sc_hd__a22o_1 _10316_ (.A1(\reg_module.gprf[427] ),
    .A2(net336),
    .B1(_04801_),
    .B2(net519),
    .X(_04802_));
 sky130_fd_sc_hd__and2_1 _10317_ (.A(net1095),
    .B(_04802_),
    .X(_00529_));
 sky130_fd_sc_hd__nor2_1 _10318_ (.A(net693),
    .B(net495),
    .Y(_04803_));
 sky130_fd_sc_hd__a22o_1 _10319_ (.A1(\reg_module.gprf[428] ),
    .A2(net336),
    .B1(_04803_),
    .B2(net526),
    .X(_04804_));
 sky130_fd_sc_hd__and2_1 _10320_ (.A(net1114),
    .B(_04804_),
    .X(_00530_));
 sky130_fd_sc_hd__nor2_1 _10321_ (.A(net694),
    .B(net493),
    .Y(_04805_));
 sky130_fd_sc_hd__a22o_1 _10322_ (.A1(\reg_module.gprf[429] ),
    .A2(net336),
    .B1(_04805_),
    .B2(net512),
    .X(_04806_));
 sky130_fd_sc_hd__and2_1 _10323_ (.A(net1078),
    .B(_04806_),
    .X(_00531_));
 sky130_fd_sc_hd__nor2_1 _10324_ (.A(net696),
    .B(net493),
    .Y(_04807_));
 sky130_fd_sc_hd__a22o_1 _10325_ (.A1(\reg_module.gprf[430] ),
    .A2(net336),
    .B1(_04807_),
    .B2(net537),
    .X(_04808_));
 sky130_fd_sc_hd__and2_1 _10326_ (.A(net1116),
    .B(_04808_),
    .X(_00532_));
 sky130_fd_sc_hd__nor2_1 _10327_ (.A(net695),
    .B(net495),
    .Y(_04809_));
 sky130_fd_sc_hd__a22o_1 _10328_ (.A1(\reg_module.gprf[431] ),
    .A2(net338),
    .B1(_04809_),
    .B2(net544),
    .X(_04810_));
 sky130_fd_sc_hd__and2_1 _10329_ (.A(net1156),
    .B(_04810_),
    .X(_00533_));
 sky130_fd_sc_hd__nor2_1 _10330_ (.A(net698),
    .B(net496),
    .Y(_04811_));
 sky130_fd_sc_hd__a22o_1 _10331_ (.A1(\reg_module.gprf[432] ),
    .A2(net339),
    .B1(_04811_),
    .B2(net565),
    .X(_04812_));
 sky130_fd_sc_hd__and2_1 _10332_ (.A(net1189),
    .B(_04812_),
    .X(_00534_));
 sky130_fd_sc_hd__nor2_1 _10333_ (.A(net697),
    .B(net495),
    .Y(_04813_));
 sky130_fd_sc_hd__a22o_1 _10334_ (.A1(\reg_module.gprf[433] ),
    .A2(net338),
    .B1(_04813_),
    .B2(net539),
    .X(_04814_));
 sky130_fd_sc_hd__and2_1 _10335_ (.A(net1141),
    .B(_04814_),
    .X(_00535_));
 sky130_fd_sc_hd__nor2_1 _10336_ (.A(net700),
    .B(net493),
    .Y(_04815_));
 sky130_fd_sc_hd__a22o_1 _10337_ (.A1(\reg_module.gprf[434] ),
    .A2(net336),
    .B1(_04815_),
    .B2(net522),
    .X(_04816_));
 sky130_fd_sc_hd__and2_1 _10338_ (.A(net1101),
    .B(_04816_),
    .X(_00536_));
 sky130_fd_sc_hd__nor2_1 _10339_ (.A(net699),
    .B(net495),
    .Y(_04817_));
 sky130_fd_sc_hd__a22o_1 _10340_ (.A1(\reg_module.gprf[435] ),
    .A2(net338),
    .B1(_04817_),
    .B2(net543),
    .X(_04818_));
 sky130_fd_sc_hd__and2_1 _10341_ (.A(net1153),
    .B(_04818_),
    .X(_00537_));
 sky130_fd_sc_hd__nor2_1 _10342_ (.A(net702),
    .B(net493),
    .Y(_04819_));
 sky130_fd_sc_hd__a22o_1 _10343_ (.A1(\reg_module.gprf[436] ),
    .A2(net337),
    .B1(_04819_),
    .B2(net527),
    .X(_04820_));
 sky130_fd_sc_hd__and2_1 _10344_ (.A(net1114),
    .B(_04820_),
    .X(_00538_));
 sky130_fd_sc_hd__nor2_1 _10345_ (.A(net701),
    .B(net496),
    .Y(_04821_));
 sky130_fd_sc_hd__a22o_1 _10346_ (.A1(\reg_module.gprf[437] ),
    .A2(net339),
    .B1(_04821_),
    .B2(net563),
    .X(_04822_));
 sky130_fd_sc_hd__and2_1 _10347_ (.A(net1201),
    .B(_04822_),
    .X(_00539_));
 sky130_fd_sc_hd__nor2_1 _10348_ (.A(net704),
    .B(net496),
    .Y(_04823_));
 sky130_fd_sc_hd__a22o_1 _10349_ (.A1(\reg_module.gprf[438] ),
    .A2(net339),
    .B1(_04823_),
    .B2(net564),
    .X(_04824_));
 sky130_fd_sc_hd__and2_1 _10350_ (.A(net1195),
    .B(_04824_),
    .X(_00540_));
 sky130_fd_sc_hd__nor2_1 _10351_ (.A(net703),
    .B(net495),
    .Y(_04825_));
 sky130_fd_sc_hd__a22o_1 _10352_ (.A1(\reg_module.gprf[439] ),
    .A2(net338),
    .B1(_04825_),
    .B2(net547),
    .X(_04826_));
 sky130_fd_sc_hd__and2_1 _10353_ (.A(net1166),
    .B(_04826_),
    .X(_00541_));
 sky130_fd_sc_hd__nor2_1 _10354_ (.A(net705),
    .B(net495),
    .Y(_04827_));
 sky130_fd_sc_hd__a22o_1 _10355_ (.A1(\reg_module.gprf[440] ),
    .A2(net338),
    .B1(_04827_),
    .B2(net554),
    .X(_04828_));
 sky130_fd_sc_hd__and2_1 _10356_ (.A(net1182),
    .B(_04828_),
    .X(_00542_));
 sky130_fd_sc_hd__nor2_1 _10357_ (.A(net706),
    .B(net495),
    .Y(_04829_));
 sky130_fd_sc_hd__a22o_1 _10358_ (.A1(\reg_module.gprf[441] ),
    .A2(net338),
    .B1(_04829_),
    .B2(net553),
    .X(_04830_));
 sky130_fd_sc_hd__and2_1 _10359_ (.A(net1180),
    .B(_04830_),
    .X(_00543_));
 sky130_fd_sc_hd__nor2_1 _10360_ (.A(_02786_),
    .B(net496),
    .Y(_04831_));
 sky130_fd_sc_hd__a22o_1 _10361_ (.A1(\reg_module.gprf[442] ),
    .A2(net338),
    .B1(_04831_),
    .B2(net545),
    .X(_04832_));
 sky130_fd_sc_hd__and2_1 _10362_ (.A(net1162),
    .B(_04832_),
    .X(_00544_));
 sky130_fd_sc_hd__nor2_1 _10363_ (.A(net707),
    .B(net495),
    .Y(_04833_));
 sky130_fd_sc_hd__a22o_1 _10364_ (.A1(\reg_module.gprf[443] ),
    .A2(net338),
    .B1(_04833_),
    .B2(net540),
    .X(_04834_));
 sky130_fd_sc_hd__and2_1 _10365_ (.A(net1145),
    .B(_04834_),
    .X(_00545_));
 sky130_fd_sc_hd__nor2_1 _10366_ (.A(net710),
    .B(net495),
    .Y(_04835_));
 sky130_fd_sc_hd__a22o_1 _10367_ (.A1(\reg_module.gprf[444] ),
    .A2(net338),
    .B1(_04835_),
    .B2(net550),
    .X(_04836_));
 sky130_fd_sc_hd__and2_1 _10368_ (.A(net1172),
    .B(_04836_),
    .X(_00546_));
 sky130_fd_sc_hd__nor2_1 _10369_ (.A(net709),
    .B(net495),
    .Y(_04837_));
 sky130_fd_sc_hd__a22o_1 _10370_ (.A1(\reg_module.gprf[445] ),
    .A2(net338),
    .B1(_04837_),
    .B2(net551),
    .X(_04838_));
 sky130_fd_sc_hd__and2_1 _10371_ (.A(net1175),
    .B(_04838_),
    .X(_00547_));
 sky130_fd_sc_hd__nor2_1 _10372_ (.A(net711),
    .B(net496),
    .Y(_04839_));
 sky130_fd_sc_hd__a22o_1 _10373_ (.A1(\reg_module.gprf[446] ),
    .A2(net339),
    .B1(_04839_),
    .B2(net558),
    .X(_04840_));
 sky130_fd_sc_hd__and2_1 _10374_ (.A(net1194),
    .B(_04840_),
    .X(_00548_));
 sky130_fd_sc_hd__nor2_1 _10375_ (.A(net574),
    .B(net496),
    .Y(_04841_));
 sky130_fd_sc_hd__a22o_1 _10376_ (.A1(\reg_module.gprf[447] ),
    .A2(net339),
    .B1(_04841_),
    .B2(net561),
    .X(_04842_));
 sky130_fd_sc_hd__and2_1 _10377_ (.A(net1205),
    .B(_04842_),
    .X(_00549_));
 sky130_fd_sc_hd__or4_4 _10378_ (.A(_01213_),
    .B(net970),
    .C(net968),
    .D(net967),
    .X(_04843_));
 sky130_fd_sc_hd__or2_4 _10379_ (.A(_04175_),
    .B(net632),
    .X(_04844_));
 sky130_fd_sc_hd__nor2_1 _10380_ (.A(_02685_),
    .B(net632),
    .Y(_04845_));
 sky130_fd_sc_hd__a22o_1 _10381_ (.A1(\reg_module.gprf[448] ),
    .A2(net333),
    .B1(_04845_),
    .B2(net532),
    .X(_04846_));
 sky130_fd_sc_hd__and2_1 _10382_ (.A(net1125),
    .B(_04846_),
    .X(_00550_));
 sky130_fd_sc_hd__nor2_1 _10383_ (.A(net721),
    .B(net632),
    .Y(_04847_));
 sky130_fd_sc_hd__a22o_1 _10384_ (.A1(\reg_module.gprf[449] ),
    .A2(net333),
    .B1(_04847_),
    .B2(net536),
    .X(_04848_));
 sky130_fd_sc_hd__and2_1 _10385_ (.A(net1132),
    .B(_04848_),
    .X(_00551_));
 sky130_fd_sc_hd__nor2_1 _10386_ (.A(_02703_),
    .B(net631),
    .Y(_04849_));
 sky130_fd_sc_hd__a22o_1 _10387_ (.A1(\reg_module.gprf[450] ),
    .A2(net333),
    .B1(_04849_),
    .B2(net525),
    .X(_04850_));
 sky130_fd_sc_hd__and2_1 _10388_ (.A(net1112),
    .B(_04850_),
    .X(_00552_));
 sky130_fd_sc_hd__nor2_1 _10389_ (.A(net712),
    .B(net631),
    .Y(_04851_));
 sky130_fd_sc_hd__a22o_1 _10390_ (.A1(\reg_module.gprf[451] ),
    .A2(net332),
    .B1(_04851_),
    .B2(net516),
    .X(_04852_));
 sky130_fd_sc_hd__and2_1 _10391_ (.A(net1088),
    .B(_04852_),
    .X(_00553_));
 sky130_fd_sc_hd__nor2_1 _10392_ (.A(_02642_),
    .B(net632),
    .Y(_04853_));
 sky130_fd_sc_hd__a22o_1 _10393_ (.A1(\reg_module.gprf[452] ),
    .A2(net333),
    .B1(_04853_),
    .B2(net533),
    .X(_04854_));
 sky130_fd_sc_hd__and2_1 _10394_ (.A(net1130),
    .B(_04854_),
    .X(_00554_));
 sky130_fd_sc_hd__nor2_1 _10395_ (.A(_02654_),
    .B(net632),
    .Y(_04855_));
 sky130_fd_sc_hd__a22o_1 _10396_ (.A1(\reg_module.gprf[453] ),
    .A2(net333),
    .B1(_04855_),
    .B2(net529),
    .X(_04856_));
 sky130_fd_sc_hd__and2_1 _10397_ (.A(net1120),
    .B(_04856_),
    .X(_00555_));
 sky130_fd_sc_hd__nor2_1 _10398_ (.A(net725),
    .B(net631),
    .Y(_04857_));
 sky130_fd_sc_hd__a22o_1 _10399_ (.A1(\reg_module.gprf[454] ),
    .A2(net332),
    .B1(_04857_),
    .B2(net513),
    .X(_04858_));
 sky130_fd_sc_hd__and2_1 _10400_ (.A(net1082),
    .B(_04858_),
    .X(_00556_));
 sky130_fd_sc_hd__nor2_1 _10401_ (.A(net724),
    .B(net631),
    .Y(_04859_));
 sky130_fd_sc_hd__a22o_1 _10402_ (.A1(\reg_module.gprf[455] ),
    .A2(net332),
    .B1(_04859_),
    .B2(net514),
    .X(_04860_));
 sky130_fd_sc_hd__and2_1 _10403_ (.A(net1086),
    .B(_04860_),
    .X(_00557_));
 sky130_fd_sc_hd__nor2_1 _10404_ (.A(net689),
    .B(net632),
    .Y(_04861_));
 sky130_fd_sc_hd__a22o_1 _10405_ (.A1(\reg_module.gprf[456] ),
    .A2(net333),
    .B1(_04861_),
    .B2(net531),
    .X(_04862_));
 sky130_fd_sc_hd__and2_1 _10406_ (.A(net1122),
    .B(_04862_),
    .X(_00558_));
 sky130_fd_sc_hd__nor2_1 _10407_ (.A(net690),
    .B(net631),
    .Y(_04863_));
 sky130_fd_sc_hd__a22o_1 _10408_ (.A1(\reg_module.gprf[457] ),
    .A2(net332),
    .B1(_04863_),
    .B2(net518),
    .X(_04864_));
 sky130_fd_sc_hd__and2_1 _10409_ (.A(net1094),
    .B(_04864_),
    .X(_00559_));
 sky130_fd_sc_hd__nor2_1 _10410_ (.A(net692),
    .B(net631),
    .Y(_04865_));
 sky130_fd_sc_hd__a22o_1 _10411_ (.A1(\reg_module.gprf[458] ),
    .A2(net332),
    .B1(_04865_),
    .B2(net511),
    .X(_04866_));
 sky130_fd_sc_hd__and2_1 _10412_ (.A(net1074),
    .B(_04866_),
    .X(_00560_));
 sky130_fd_sc_hd__nor2_1 _10413_ (.A(net691),
    .B(net631),
    .Y(_04867_));
 sky130_fd_sc_hd__a22o_1 _10414_ (.A1(\reg_module.gprf[459] ),
    .A2(net332),
    .B1(_04867_),
    .B2(net520),
    .X(_04868_));
 sky130_fd_sc_hd__and2_1 _10415_ (.A(net1099),
    .B(_04868_),
    .X(_00561_));
 sky130_fd_sc_hd__nor2_1 _10416_ (.A(_03014_),
    .B(net633),
    .Y(_04869_));
 sky130_fd_sc_hd__a22o_1 _10417_ (.A1(\reg_module.gprf[460] ),
    .A2(net332),
    .B1(_04869_),
    .B2(net543),
    .X(_04870_));
 sky130_fd_sc_hd__and2_1 _10418_ (.A(net1152),
    .B(_04870_),
    .X(_00562_));
 sky130_fd_sc_hd__nor2_1 _10419_ (.A(net694),
    .B(net631),
    .Y(_04871_));
 sky130_fd_sc_hd__a22o_1 _10420_ (.A1(\reg_module.gprf[461] ),
    .A2(net332),
    .B1(_04871_),
    .B2(net523),
    .X(_04872_));
 sky130_fd_sc_hd__and2_1 _10421_ (.A(net1097),
    .B(_04872_),
    .X(_00563_));
 sky130_fd_sc_hd__nor2_1 _10422_ (.A(net696),
    .B(net631),
    .Y(_04873_));
 sky130_fd_sc_hd__a22o_1 _10423_ (.A1(\reg_module.gprf[462] ),
    .A2(net332),
    .B1(_04873_),
    .B2(net565),
    .X(_04874_));
 sky130_fd_sc_hd__and2_1 _10424_ (.A(net1155),
    .B(_04874_),
    .X(_00564_));
 sky130_fd_sc_hd__nor2_1 _10425_ (.A(net695),
    .B(net633),
    .Y(_04875_));
 sky130_fd_sc_hd__a22o_1 _10426_ (.A1(\reg_module.gprf[463] ),
    .A2(net334),
    .B1(_04875_),
    .B2(net545),
    .X(_04876_));
 sky130_fd_sc_hd__and2_1 _10427_ (.A(net1161),
    .B(_04876_),
    .X(_00565_));
 sky130_fd_sc_hd__nor2_1 _10428_ (.A(net698),
    .B(net634),
    .Y(_04877_));
 sky130_fd_sc_hd__a22o_1 _10429_ (.A1(\reg_module.gprf[464] ),
    .A2(net335),
    .B1(_04877_),
    .B2(net559),
    .X(_04878_));
 sky130_fd_sc_hd__and2_1 _10430_ (.A(net1202),
    .B(_04878_),
    .X(_00566_));
 sky130_fd_sc_hd__nor2_1 _10431_ (.A(_02951_),
    .B(net633),
    .Y(_04879_));
 sky130_fd_sc_hd__a22o_1 _10432_ (.A1(\reg_module.gprf[465] ),
    .A2(net334),
    .B1(_04879_),
    .B2(net540),
    .X(_04880_));
 sky130_fd_sc_hd__and2_1 _10433_ (.A(net1147),
    .B(_04880_),
    .X(_00567_));
 sky130_fd_sc_hd__nor2_1 _10434_ (.A(net700),
    .B(net632),
    .Y(_04881_));
 sky130_fd_sc_hd__a22o_1 _10435_ (.A1(\reg_module.gprf[466] ),
    .A2(net332),
    .B1(_04881_),
    .B2(net538),
    .X(_04882_));
 sky130_fd_sc_hd__and2_1 _10436_ (.A(net1139),
    .B(_04882_),
    .X(_00568_));
 sky130_fd_sc_hd__nor2_1 _10437_ (.A(net699),
    .B(net633),
    .Y(_04883_));
 sky130_fd_sc_hd__a22o_1 _10438_ (.A1(\reg_module.gprf[467] ),
    .A2(net334),
    .B1(_04883_),
    .B2(net546),
    .X(_04884_));
 sky130_fd_sc_hd__and2_1 _10439_ (.A(net1158),
    .B(_04884_),
    .X(_00569_));
 sky130_fd_sc_hd__nor2_1 _10440_ (.A(_02881_),
    .B(net631),
    .Y(_04885_));
 sky130_fd_sc_hd__a22o_1 _10441_ (.A1(\reg_module.gprf[468] ),
    .A2(net333),
    .B1(_04885_),
    .B2(net543),
    .X(_04886_));
 sky130_fd_sc_hd__and2_1 _10442_ (.A(net1152),
    .B(_04886_),
    .X(_00570_));
 sky130_fd_sc_hd__nor2_1 _10443_ (.A(_02894_),
    .B(net634),
    .Y(_04887_));
 sky130_fd_sc_hd__a22o_1 _10444_ (.A1(\reg_module.gprf[469] ),
    .A2(net335),
    .B1(_04887_),
    .B2(net561),
    .X(_04888_));
 sky130_fd_sc_hd__and2_1 _10445_ (.A(net1207),
    .B(_04888_),
    .X(_00571_));
 sky130_fd_sc_hd__nor2_1 _10446_ (.A(_02850_),
    .B(net634),
    .Y(_04889_));
 sky130_fd_sc_hd__a22o_1 _10447_ (.A1(\reg_module.gprf[470] ),
    .A2(net335),
    .B1(_04889_),
    .B2(net557),
    .X(_04890_));
 sky130_fd_sc_hd__and2_1 _10448_ (.A(net1196),
    .B(_04890_),
    .X(_00572_));
 sky130_fd_sc_hd__nor2_1 _10449_ (.A(net703),
    .B(net633),
    .Y(_04891_));
 sky130_fd_sc_hd__a22o_1 _10450_ (.A1(\reg_module.gprf[471] ),
    .A2(net334),
    .B1(_04891_),
    .B2(net548),
    .X(_04892_));
 sky130_fd_sc_hd__and2_1 _10451_ (.A(net1165),
    .B(_04892_),
    .X(_00573_));
 sky130_fd_sc_hd__nor2_1 _10452_ (.A(_02832_),
    .B(net633),
    .Y(_04893_));
 sky130_fd_sc_hd__a22o_1 _10453_ (.A1(\reg_module.gprf[472] ),
    .A2(net334),
    .B1(_04893_),
    .B2(net554),
    .X(_04894_));
 sky130_fd_sc_hd__and2_1 _10454_ (.A(net1183),
    .B(_04894_),
    .X(_00574_));
 sky130_fd_sc_hd__nor2_1 _10455_ (.A(net706),
    .B(net633),
    .Y(_04895_));
 sky130_fd_sc_hd__a22o_1 _10456_ (.A1(\reg_module.gprf[473] ),
    .A2(net334),
    .B1(_04895_),
    .B2(net553),
    .X(_04896_));
 sky130_fd_sc_hd__and2_1 _10457_ (.A(net1180),
    .B(_04896_),
    .X(_00575_));
 sky130_fd_sc_hd__nor2_1 _10458_ (.A(_02786_),
    .B(net633),
    .Y(_04897_));
 sky130_fd_sc_hd__a22o_1 _10459_ (.A1(\reg_module.gprf[474] ),
    .A2(net334),
    .B1(_04897_),
    .B2(net565),
    .X(_04898_));
 sky130_fd_sc_hd__and2_1 _10460_ (.A(net1162),
    .B(_04898_),
    .X(_00576_));
 sky130_fd_sc_hd__nor2_1 _10461_ (.A(net707),
    .B(net633),
    .Y(_04899_));
 sky130_fd_sc_hd__a22o_1 _10462_ (.A1(\reg_module.gprf[475] ),
    .A2(net334),
    .B1(_04899_),
    .B2(net540),
    .X(_04900_));
 sky130_fd_sc_hd__and2_1 _10463_ (.A(net1146),
    .B(_04900_),
    .X(_00577_));
 sky130_fd_sc_hd__nor2_1 _10464_ (.A(net710),
    .B(net633),
    .Y(_04901_));
 sky130_fd_sc_hd__a22o_1 _10465_ (.A1(\reg_module.gprf[476] ),
    .A2(net334),
    .B1(_04901_),
    .B2(net550),
    .X(_04902_));
 sky130_fd_sc_hd__and2_1 _10466_ (.A(net1172),
    .B(_04902_),
    .X(_00578_));
 sky130_fd_sc_hd__nor2_1 _10467_ (.A(net709),
    .B(net634),
    .Y(_04903_));
 sky130_fd_sc_hd__a22o_1 _10468_ (.A1(\reg_module.gprf[477] ),
    .A2(net334),
    .B1(_04903_),
    .B2(net551),
    .X(_04904_));
 sky130_fd_sc_hd__and2_1 _10469_ (.A(net1175),
    .B(_04904_),
    .X(_00579_));
 sky130_fd_sc_hd__nor2_1 _10470_ (.A(net711),
    .B(net634),
    .Y(_04905_));
 sky130_fd_sc_hd__a22o_1 _10471_ (.A1(\reg_module.gprf[478] ),
    .A2(net335),
    .B1(_04905_),
    .B2(net558),
    .X(_04906_));
 sky130_fd_sc_hd__and2_1 _10472_ (.A(net1193),
    .B(_04906_),
    .X(_00580_));
 sky130_fd_sc_hd__nor2_1 _10473_ (.A(_02585_),
    .B(net634),
    .Y(_04907_));
 sky130_fd_sc_hd__a22o_1 _10474_ (.A1(\reg_module.gprf[479] ),
    .A2(net335),
    .B1(_04907_),
    .B2(net562),
    .X(_04908_));
 sky130_fd_sc_hd__and2_1 _10475_ (.A(net1205),
    .B(_04908_),
    .X(_00581_));
 sky130_fd_sc_hd__nor2_4 _10476_ (.A(_01254_),
    .B(_04175_),
    .Y(_04909_));
 sky130_fd_sc_hd__mux2_1 _10477_ (.A0(\reg_module.gprf[480] ),
    .A1(_02686_),
    .S(net328),
    .X(_04910_));
 sky130_fd_sc_hd__and2_1 _10478_ (.A(net1091),
    .B(_04910_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _10479_ (.A0(\reg_module.gprf[481] ),
    .A1(_02672_),
    .S(net329),
    .X(_04911_));
 sky130_fd_sc_hd__and2_1 _10480_ (.A(net1132),
    .B(_04911_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _10481_ (.A0(\reg_module.gprf[482] ),
    .A1(_02702_),
    .S(net328),
    .X(_04912_));
 sky130_fd_sc_hd__and2_1 _10482_ (.A(net1110),
    .B(_04912_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _10483_ (.A0(\reg_module.gprf[483] ),
    .A1(_02716_),
    .S(net328),
    .X(_04913_));
 sky130_fd_sc_hd__and2_1 _10484_ (.A(net1088),
    .B(_04913_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _10485_ (.A0(\reg_module.gprf[484] ),
    .A1(_02641_),
    .S(net329),
    .X(_04914_));
 sky130_fd_sc_hd__and2_1 _10486_ (.A(net1130),
    .B(_04914_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _10487_ (.A0(\reg_module.gprf[485] ),
    .A1(_02655_),
    .S(net329),
    .X(_04915_));
 sky130_fd_sc_hd__and2_1 _10488_ (.A(net1120),
    .B(_04915_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _10489_ (.A0(\reg_module.gprf[486] ),
    .A1(_02605_),
    .S(net328),
    .X(_04916_));
 sky130_fd_sc_hd__and2_1 _10490_ (.A(net1082),
    .B(_04916_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _10491_ (.A0(\reg_module.gprf[487] ),
    .A1(_02624_),
    .S(net328),
    .X(_04917_));
 sky130_fd_sc_hd__and2_1 _10492_ (.A(net1089),
    .B(_04917_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _10493_ (.A0(\reg_module.gprf[488] ),
    .A1(_03078_),
    .S(net329),
    .X(_04918_));
 sky130_fd_sc_hd__and2_1 _10494_ (.A(net1122),
    .B(_04918_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _10495_ (.A0(\reg_module.gprf[489] ),
    .A1(_03062_),
    .S(net328),
    .X(_04919_));
 sky130_fd_sc_hd__and2_1 _10496_ (.A(net1096),
    .B(_04919_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _10497_ (.A0(\reg_module.gprf[490] ),
    .A1(_03031_),
    .S(net328),
    .X(_04920_));
 sky130_fd_sc_hd__and2_1 _10498_ (.A(net1074),
    .B(_04920_),
    .X(_00592_));
 sky130_fd_sc_hd__mux2_1 _10499_ (.A0(\reg_module.gprf[491] ),
    .A1(_03045_),
    .S(net328),
    .X(_04921_));
 sky130_fd_sc_hd__and2_1 _10500_ (.A(net1100),
    .B(_04921_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _10501_ (.A0(\reg_module.gprf[492] ),
    .A1(_03015_),
    .S(net328),
    .X(_04922_));
 sky130_fd_sc_hd__and2_1 _10502_ (.A(net1114),
    .B(_04922_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _10503_ (.A0(\reg_module.gprf[493] ),
    .A1(_03001_),
    .S(net328),
    .X(_04923_));
 sky130_fd_sc_hd__and2_1 _10504_ (.A(net1106),
    .B(_04923_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _10505_ (.A0(\reg_module.gprf[494] ),
    .A1(_02970_),
    .S(net329),
    .X(_04924_));
 sky130_fd_sc_hd__and2_1 _10506_ (.A(net1188),
    .B(_04924_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _10507_ (.A0(\reg_module.gprf[495] ),
    .A1(_02985_),
    .S(net330),
    .X(_04925_));
 sky130_fd_sc_hd__and2_1 _10508_ (.A(net1156),
    .B(_04925_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _10509_ (.A0(\reg_module.gprf[496] ),
    .A1(_02939_),
    .S(net331),
    .X(_04926_));
 sky130_fd_sc_hd__and2_1 _10510_ (.A(net1189),
    .B(_04926_),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _10511_ (.A0(\reg_module.gprf[497] ),
    .A1(_02952_),
    .S(net330),
    .X(_04927_));
 sky130_fd_sc_hd__and2_1 _10512_ (.A(net1141),
    .B(_04927_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _10513_ (.A0(\reg_module.gprf[498] ),
    .A1(_02910_),
    .S(net330),
    .X(_04928_));
 sky130_fd_sc_hd__and2_1 _10514_ (.A(net1141),
    .B(_04928_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _10515_ (.A0(\reg_module.gprf[499] ),
    .A1(_02924_),
    .S(net330),
    .X(_04929_));
 sky130_fd_sc_hd__and2_1 _10516_ (.A(net1153),
    .B(_04929_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _10517_ (.A0(\reg_module.gprf[500] ),
    .A1(_02882_),
    .S(net330),
    .X(_04930_));
 sky130_fd_sc_hd__and2_1 _10518_ (.A(net1152),
    .B(_04930_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _10519_ (.A0(\reg_module.gprf[501] ),
    .A1(_02895_),
    .S(net331),
    .X(_04931_));
 sky130_fd_sc_hd__and2_1 _10520_ (.A(net1201),
    .B(_04931_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _10521_ (.A0(\reg_module.gprf[502] ),
    .A1(_02851_),
    .S(net331),
    .X(_04932_));
 sky130_fd_sc_hd__and2_1 _10522_ (.A(net1195),
    .B(_04932_),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _10523_ (.A0(\reg_module.gprf[503] ),
    .A1(_02865_),
    .S(net330),
    .X(_04933_));
 sky130_fd_sc_hd__and2_1 _10524_ (.A(net1166),
    .B(_04933_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _10525_ (.A0(\reg_module.gprf[504] ),
    .A1(_02833_),
    .S(net330),
    .X(_04934_));
 sky130_fd_sc_hd__and2_1 _10526_ (.A(net1182),
    .B(_04934_),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _10527_ (.A0(\reg_module.gprf[505] ),
    .A1(_02817_),
    .S(net330),
    .X(_04935_));
 sky130_fd_sc_hd__and2_1 _10528_ (.A(net1181),
    .B(_04935_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _10529_ (.A0(\reg_module.gprf[506] ),
    .A1(_02787_),
    .S(net330),
    .X(_04936_));
 sky130_fd_sc_hd__and2_1 _10530_ (.A(net1162),
    .B(_04936_),
    .X(_00608_));
 sky130_fd_sc_hd__mux2_1 _10531_ (.A0(\reg_module.gprf[507] ),
    .A1(_02801_),
    .S(net331),
    .X(_04937_));
 sky130_fd_sc_hd__and2_1 _10532_ (.A(net1147),
    .B(_04937_),
    .X(_00609_));
 sky130_fd_sc_hd__mux2_1 _10533_ (.A0(\reg_module.gprf[508] ),
    .A1(_02757_),
    .S(net330),
    .X(_04938_));
 sky130_fd_sc_hd__and2_1 _10534_ (.A(net1171),
    .B(_04938_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _10535_ (.A0(\reg_module.gprf[509] ),
    .A1(_02771_),
    .S(net331),
    .X(_04939_));
 sky130_fd_sc_hd__and2_1 _10536_ (.A(net1178),
    .B(_04939_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _10537_ (.A0(\reg_module.gprf[510] ),
    .A1(_02743_),
    .S(net331),
    .X(_04940_));
 sky130_fd_sc_hd__and2_1 _10538_ (.A(net1190),
    .B(_04940_),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _10539_ (.A0(\reg_module.gprf[511] ),
    .A1(_02586_),
    .S(net331),
    .X(_04941_));
 sky130_fd_sc_hd__and2_1 _10540_ (.A(net1204),
    .B(_04941_),
    .X(_00613_));
 sky130_fd_sc_hd__and3b_2 _10541_ (.A_N(\rReg_d2[4] ),
    .B(_01974_),
    .C(_04139_),
    .X(_04942_));
 sky130_fd_sc_hd__mux2_1 _10542_ (.A0(\reg_module.gprf[512] ),
    .A1(_02686_),
    .S(net489),
    .X(_04943_));
 sky130_fd_sc_hd__and2_1 _10543_ (.A(net1135),
    .B(_04943_),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_1 _10544_ (.A0(\reg_module.gprf[513] ),
    .A1(_02672_),
    .S(net490),
    .X(_04944_));
 sky130_fd_sc_hd__and2_1 _10545_ (.A(net1132),
    .B(_04944_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _10546_ (.A0(\reg_module.gprf[514] ),
    .A1(_02702_),
    .S(net489),
    .X(_04945_));
 sky130_fd_sc_hd__and2_1 _10547_ (.A(net1090),
    .B(_04945_),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _10548_ (.A0(\reg_module.gprf[515] ),
    .A1(_02716_),
    .S(net489),
    .X(_04946_));
 sky130_fd_sc_hd__and2_1 _10549_ (.A(net1087),
    .B(_04946_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _10550_ (.A0(\reg_module.gprf[516] ),
    .A1(_02641_),
    .S(net490),
    .X(_04947_));
 sky130_fd_sc_hd__and2_1 _10551_ (.A(net1128),
    .B(_04947_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _10552_ (.A0(\reg_module.gprf[517] ),
    .A1(_02655_),
    .S(net490),
    .X(_04948_));
 sky130_fd_sc_hd__and2_1 _10553_ (.A(net1120),
    .B(_04948_),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _10554_ (.A0(\reg_module.gprf[518] ),
    .A1(_02605_),
    .S(net489),
    .X(_04949_));
 sky130_fd_sc_hd__and2_1 _10555_ (.A(net1072),
    .B(_04949_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _10556_ (.A0(\reg_module.gprf[519] ),
    .A1(_02624_),
    .S(net489),
    .X(_04950_));
 sky130_fd_sc_hd__and2_1 _10557_ (.A(net1089),
    .B(_04950_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _10558_ (.A0(\reg_module.gprf[520] ),
    .A1(_03078_),
    .S(net490),
    .X(_04951_));
 sky130_fd_sc_hd__and2_1 _10559_ (.A(net1125),
    .B(_04951_),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _10560_ (.A0(\reg_module.gprf[521] ),
    .A1(_03062_),
    .S(net489),
    .X(_04952_));
 sky130_fd_sc_hd__and2_1 _10561_ (.A(net1097),
    .B(_04952_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _10562_ (.A0(\reg_module.gprf[522] ),
    .A1(_03031_),
    .S(net489),
    .X(_04953_));
 sky130_fd_sc_hd__and2_1 _10563_ (.A(net1077),
    .B(_04953_),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _10564_ (.A0(\reg_module.gprf[523] ),
    .A1(_03045_),
    .S(net490),
    .X(_04954_));
 sky130_fd_sc_hd__and2_1 _10565_ (.A(net1102),
    .B(_04954_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _10566_ (.A0(\reg_module.gprf[524] ),
    .A1(_03015_),
    .S(net489),
    .X(_04955_));
 sky130_fd_sc_hd__and2_1 _10567_ (.A(net1114),
    .B(_04955_),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _10568_ (.A0(\reg_module.gprf[525] ),
    .A1(_03001_),
    .S(net490),
    .X(_04956_));
 sky130_fd_sc_hd__and2_1 _10569_ (.A(net1108),
    .B(_04956_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _10570_ (.A0(\reg_module.gprf[526] ),
    .A1(_02970_),
    .S(net489),
    .X(_04957_));
 sky130_fd_sc_hd__and2_1 _10571_ (.A(net1135),
    .B(_04957_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _10572_ (.A0(\reg_module.gprf[527] ),
    .A1(_02985_),
    .S(net491),
    .X(_04958_));
 sky130_fd_sc_hd__and2_1 _10573_ (.A(net1156),
    .B(_04958_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _10574_ (.A0(\reg_module.gprf[528] ),
    .A1(_02939_),
    .S(net492),
    .X(_04959_));
 sky130_fd_sc_hd__and2_1 _10575_ (.A(net1189),
    .B(_04959_),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _10576_ (.A0(\reg_module.gprf[529] ),
    .A1(_02952_),
    .S(net491),
    .X(_04960_));
 sky130_fd_sc_hd__and2_1 _10577_ (.A(net1142),
    .B(_04960_),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _10578_ (.A0(\reg_module.gprf[530] ),
    .A1(_02910_),
    .S(net491),
    .X(_04961_));
 sky130_fd_sc_hd__and2_1 _10579_ (.A(net1143),
    .B(_04961_),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _10580_ (.A0(\reg_module.gprf[531] ),
    .A1(_02924_),
    .S(net491),
    .X(_04962_));
 sky130_fd_sc_hd__and2_1 _10581_ (.A(net1142),
    .B(_04962_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _10582_ (.A0(\reg_module.gprf[532] ),
    .A1(_02882_),
    .S(net489),
    .X(_04963_));
 sky130_fd_sc_hd__and2_1 _10583_ (.A(net1116),
    .B(_04963_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _10584_ (.A0(\reg_module.gprf[533] ),
    .A1(_02895_),
    .S(net492),
    .X(_04964_));
 sky130_fd_sc_hd__and2_1 _10585_ (.A(net1201),
    .B(_04964_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _10586_ (.A0(\reg_module.gprf[534] ),
    .A1(_02851_),
    .S(net492),
    .X(_04965_));
 sky130_fd_sc_hd__and2_1 _10587_ (.A(net1191),
    .B(_04965_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _10588_ (.A0(\reg_module.gprf[535] ),
    .A1(_02865_),
    .S(net491),
    .X(_04966_));
 sky130_fd_sc_hd__and2_1 _10589_ (.A(net1167),
    .B(_04966_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _10590_ (.A0(\reg_module.gprf[536] ),
    .A1(_02833_),
    .S(net491),
    .X(_04967_));
 sky130_fd_sc_hd__and2_1 _10591_ (.A(net1178),
    .B(_04967_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _10592_ (.A0(\reg_module.gprf[537] ),
    .A1(_02817_),
    .S(net491),
    .X(_04968_));
 sky130_fd_sc_hd__and2_1 _10593_ (.A(net1176),
    .B(_04968_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _10594_ (.A0(\reg_module.gprf[538] ),
    .A1(_02787_),
    .S(net491),
    .X(_04969_));
 sky130_fd_sc_hd__and2_1 _10595_ (.A(net1188),
    .B(_04969_),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _10596_ (.A0(\reg_module.gprf[539] ),
    .A1(_02801_),
    .S(net491),
    .X(_04970_));
 sky130_fd_sc_hd__and2_1 _10597_ (.A(net1150),
    .B(_04970_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _10598_ (.A0(\reg_module.gprf[540] ),
    .A1(_02757_),
    .S(net491),
    .X(_04971_));
 sky130_fd_sc_hd__and2_1 _10599_ (.A(net1168),
    .B(_04971_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _10600_ (.A0(\reg_module.gprf[541] ),
    .A1(_02771_),
    .S(net492),
    .X(_04972_));
 sky130_fd_sc_hd__and2_1 _10601_ (.A(net1175),
    .B(_04972_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _10602_ (.A0(\reg_module.gprf[542] ),
    .A1(_02743_),
    .S(net492),
    .X(_04973_));
 sky130_fd_sc_hd__and2_1 _10603_ (.A(net1190),
    .B(_04973_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _10604_ (.A0(\reg_module.gprf[543] ),
    .A1(_02586_),
    .S(net492),
    .X(_04974_));
 sky130_fd_sc_hd__and2_1 _10605_ (.A(net1199),
    .B(_04974_),
    .X(_00645_));
 sky130_fd_sc_hd__and2_1 _10606_ (.A(_01974_),
    .B(_04173_),
    .X(_04975_));
 sky130_fd_sc_hd__nand2_2 _10607_ (.A(_01974_),
    .B(_04173_),
    .Y(_04976_));
 sky130_fd_sc_hd__nand3_4 _10608_ (.A(net966),
    .B(net674),
    .C(net454),
    .Y(_04977_));
 sky130_fd_sc_hd__a32o_1 _10609_ (.A1(net673),
    .A2(_04181_),
    .A3(net453),
    .B1(net324),
    .B2(\reg_module.gprf[544] ),
    .X(_04978_));
 sky130_fd_sc_hd__and2_1 _10610_ (.A(net1091),
    .B(_04978_),
    .X(_00646_));
 sky130_fd_sc_hd__a32o_1 _10611_ (.A1(net674),
    .A2(net417),
    .A3(net455),
    .B1(net325),
    .B2(\reg_module.gprf[545] ),
    .X(_04979_));
 sky130_fd_sc_hd__and2_1 _10612_ (.A(net1130),
    .B(_04979_),
    .X(_00647_));
 sky130_fd_sc_hd__a32o_1 _10613_ (.A1(net673),
    .A2(net416),
    .A3(net441),
    .B1(net324),
    .B2(\reg_module.gprf[546] ),
    .X(_04980_));
 sky130_fd_sc_hd__and2_1 _10614_ (.A(net1090),
    .B(_04980_),
    .X(_00648_));
 sky130_fd_sc_hd__a32o_1 _10615_ (.A1(net672),
    .A2(net415),
    .A3(net439),
    .B1(net324),
    .B2(\reg_module.gprf[547] ),
    .X(_04981_));
 sky130_fd_sc_hd__and2_1 _10616_ (.A(net1082),
    .B(_04981_),
    .X(_00649_));
 sky130_fd_sc_hd__a32o_1 _10617_ (.A1(net674),
    .A2(_04189_),
    .A3(net456),
    .B1(net325),
    .B2(\reg_module.gprf[548] ),
    .X(_04982_));
 sky130_fd_sc_hd__and2_1 _10618_ (.A(net1128),
    .B(_04982_),
    .X(_00650_));
 sky130_fd_sc_hd__a32o_1 _10619_ (.A1(net674),
    .A2(_04191_),
    .A3(net452),
    .B1(net324),
    .B2(\reg_module.gprf[549] ),
    .X(_04983_));
 sky130_fd_sc_hd__and2_1 _10620_ (.A(net1120),
    .B(_04983_),
    .X(_00651_));
 sky130_fd_sc_hd__a32o_1 _10621_ (.A1(net672),
    .A2(net412),
    .A3(net433),
    .B1(net324),
    .B2(\reg_module.gprf[550] ),
    .X(_04984_));
 sky130_fd_sc_hd__and2_1 _10622_ (.A(net1072),
    .B(_04984_),
    .X(_00652_));
 sky130_fd_sc_hd__a32o_1 _10623_ (.A1(net672),
    .A2(net411),
    .A3(net438),
    .B1(net324),
    .B2(\reg_module.gprf[551] ),
    .X(_04985_));
 sky130_fd_sc_hd__and2_1 _10624_ (.A(net1082),
    .B(_04985_),
    .X(_00653_));
 sky130_fd_sc_hd__a32o_1 _10625_ (.A1(net674),
    .A2(_04197_),
    .A3(net453),
    .B1(net325),
    .B2(\reg_module.gprf[552] ),
    .X(_04986_));
 sky130_fd_sc_hd__and2_1 _10626_ (.A(net1125),
    .B(_04986_),
    .X(_00654_));
 sky130_fd_sc_hd__a32o_1 _10627_ (.A1(net672),
    .A2(net409),
    .A3(net436),
    .B1(net324),
    .B2(\reg_module.gprf[553] ),
    .X(_04987_));
 sky130_fd_sc_hd__and2_1 _10628_ (.A(net1078),
    .B(_04987_),
    .X(_00655_));
 sky130_fd_sc_hd__a32o_1 _10629_ (.A1(net672),
    .A2(net408),
    .A3(net434),
    .B1(net324),
    .B2(\reg_module.gprf[554] ),
    .X(_04988_));
 sky130_fd_sc_hd__and2_1 _10630_ (.A(net1077),
    .B(_04988_),
    .X(_00656_));
 sky130_fd_sc_hd__a32o_1 _10631_ (.A1(net671),
    .A2(net407),
    .A3(net444),
    .B1(net325),
    .B2(\reg_module.gprf[555] ),
    .X(_04989_));
 sky130_fd_sc_hd__and2_1 _10632_ (.A(net1098),
    .B(_04989_),
    .X(_00657_));
 sky130_fd_sc_hd__a32o_1 _10633_ (.A1(net671),
    .A2(_04205_),
    .A3(net449),
    .B1(net325),
    .B2(\reg_module.gprf[556] ),
    .X(_04990_));
 sky130_fd_sc_hd__and2_1 _10634_ (.A(net1113),
    .B(_04990_),
    .X(_00658_));
 sky130_fd_sc_hd__a32o_1 _10635_ (.A1(net671),
    .A2(net405),
    .A3(net448),
    .B1(net324),
    .B2(\reg_module.gprf[557] ),
    .X(_04991_));
 sky130_fd_sc_hd__and2_1 _10636_ (.A(net1108),
    .B(_04991_),
    .X(_00659_));
 sky130_fd_sc_hd__a32o_1 _10637_ (.A1(net673),
    .A2(net404),
    .A3(net450),
    .B1(net324),
    .B2(\reg_module.gprf[558] ),
    .X(_04992_));
 sky130_fd_sc_hd__and2_1 _10638_ (.A(net1115),
    .B(_04992_),
    .X(_00660_));
 sky130_fd_sc_hd__a32o_1 _10639_ (.A1(net676),
    .A2(net403),
    .A3(net465),
    .B1(net326),
    .B2(\reg_module.gprf[559] ),
    .X(_04993_));
 sky130_fd_sc_hd__and2_1 _10640_ (.A(net1155),
    .B(_04993_),
    .X(_00661_));
 sky130_fd_sc_hd__a32o_1 _10641_ (.A1(net677),
    .A2(net402),
    .A3(net487),
    .B1(net327),
    .B2(\reg_module.gprf[560] ),
    .X(_04994_));
 sky130_fd_sc_hd__and2_1 _10642_ (.A(net1189),
    .B(_04994_),
    .X(_00662_));
 sky130_fd_sc_hd__a32o_1 _10643_ (.A1(net676),
    .A2(net401),
    .A3(net460),
    .B1(net326),
    .B2(\reg_module.gprf[561] ),
    .X(_04995_));
 sky130_fd_sc_hd__and2_1 _10644_ (.A(net1142),
    .B(_04995_),
    .X(_00663_));
 sky130_fd_sc_hd__a32o_1 _10645_ (.A1(net676),
    .A2(net400),
    .A3(net460),
    .B1(net326),
    .B2(\reg_module.gprf[562] ),
    .X(_04996_));
 sky130_fd_sc_hd__and2_1 _10646_ (.A(net1143),
    .B(_04996_),
    .X(_00664_));
 sky130_fd_sc_hd__a32o_1 _10647_ (.A1(net676),
    .A2(net399),
    .A3(net460),
    .B1(net326),
    .B2(\reg_module.gprf[563] ),
    .X(_04997_));
 sky130_fd_sc_hd__and2_1 _10648_ (.A(net1142),
    .B(_04997_),
    .X(_00665_));
 sky130_fd_sc_hd__a32o_1 _10649_ (.A1(net671),
    .A2(net398),
    .A3(net449),
    .B1(net325),
    .B2(\reg_module.gprf[564] ),
    .X(_04998_));
 sky130_fd_sc_hd__and2_1 _10650_ (.A(net1113),
    .B(_04998_),
    .X(_00666_));
 sky130_fd_sc_hd__a32o_1 _10651_ (.A1(net677),
    .A2(net397),
    .A3(net484),
    .B1(net327),
    .B2(\reg_module.gprf[565] ),
    .X(_04999_));
 sky130_fd_sc_hd__and2_1 _10652_ (.A(net1199),
    .B(_04999_),
    .X(_00667_));
 sky130_fd_sc_hd__a32o_1 _10653_ (.A1(net677),
    .A2(net396),
    .A3(net482),
    .B1(net327),
    .B2(\reg_module.gprf[566] ),
    .X(_05000_));
 sky130_fd_sc_hd__and2_1 _10654_ (.A(net1191),
    .B(_05000_),
    .X(_00668_));
 sky130_fd_sc_hd__a32o_1 _10655_ (.A1(net675),
    .A2(net395),
    .A3(net470),
    .B1(net326),
    .B2(\reg_module.gprf[567] ),
    .X(_05001_));
 sky130_fd_sc_hd__and2_1 _10656_ (.A(net1169),
    .B(_05001_),
    .X(_00669_));
 sky130_fd_sc_hd__a32o_1 _10657_ (.A1(net676),
    .A2(net394),
    .A3(net476),
    .B1(net326),
    .B2(\reg_module.gprf[568] ),
    .X(_05002_));
 sky130_fd_sc_hd__and2_1 _10658_ (.A(net1179),
    .B(_05002_),
    .X(_00670_));
 sky130_fd_sc_hd__a32o_1 _10659_ (.A1(net675),
    .A2(_04231_),
    .A3(net475),
    .B1(net326),
    .B2(\reg_module.gprf[569] ),
    .X(_05003_));
 sky130_fd_sc_hd__and2_1 _10660_ (.A(net1176),
    .B(_05003_),
    .X(_00671_));
 sky130_fd_sc_hd__a32o_1 _10661_ (.A1(net677),
    .A2(net392),
    .A3(net487),
    .B1(net326),
    .B2(\reg_module.gprf[570] ),
    .X(_05004_));
 sky130_fd_sc_hd__and2_1 _10662_ (.A(net1161),
    .B(_05004_),
    .X(_00672_));
 sky130_fd_sc_hd__a32o_1 _10663_ (.A1(net675),
    .A2(_04235_),
    .A3(net463),
    .B1(net326),
    .B2(\reg_module.gprf[571] ),
    .X(_05005_));
 sky130_fd_sc_hd__and2_1 _10664_ (.A(net1149),
    .B(_05005_),
    .X(_00673_));
 sky130_fd_sc_hd__a32o_1 _10665_ (.A1(net678),
    .A2(_04237_),
    .A3(net471),
    .B1(net326),
    .B2(\reg_module.gprf[572] ),
    .X(_05006_));
 sky130_fd_sc_hd__and2_1 _10666_ (.A(net1168),
    .B(_05006_),
    .X(_00674_));
 sky130_fd_sc_hd__a32o_1 _10667_ (.A1(net675),
    .A2(net389),
    .A3(net470),
    .B1(net327),
    .B2(\reg_module.gprf[573] ),
    .X(_05007_));
 sky130_fd_sc_hd__and2_1 _10668_ (.A(net1168),
    .B(_05007_),
    .X(_00675_));
 sky130_fd_sc_hd__a32o_1 _10669_ (.A1(net677),
    .A2(net388),
    .A3(net482),
    .B1(net327),
    .B2(\reg_module.gprf[574] ),
    .X(_05008_));
 sky130_fd_sc_hd__and2_1 _10670_ (.A(net1190),
    .B(_05008_),
    .X(_00676_));
 sky130_fd_sc_hd__a32o_1 _10671_ (.A1(net678),
    .A2(net387),
    .A3(net483),
    .B1(net327),
    .B2(\reg_module.gprf[575] ),
    .X(_05009_));
 sky130_fd_sc_hd__and2_1 _10672_ (.A(net1199),
    .B(_05009_),
    .X(_00677_));
 sky130_fd_sc_hd__nand3_4 _10673_ (.A(net965),
    .B(net748),
    .C(net454),
    .Y(_05010_));
 sky130_fd_sc_hd__a32o_1 _10674_ (.A1(_04181_),
    .A2(net747),
    .A3(net447),
    .B1(net320),
    .B2(\reg_module.gprf[576] ),
    .X(_05011_));
 sky130_fd_sc_hd__and2_1 _10675_ (.A(net1111),
    .B(_05011_),
    .X(_00678_));
 sky130_fd_sc_hd__a32o_1 _10676_ (.A1(net417),
    .A2(net748),
    .A3(net457),
    .B1(net321),
    .B2(\reg_module.gprf[577] ),
    .X(_05012_));
 sky130_fd_sc_hd__and2_1 _10677_ (.A(net1132),
    .B(_05012_),
    .X(_00679_));
 sky130_fd_sc_hd__a32o_1 _10678_ (.A1(net416),
    .A2(net745),
    .A3(net441),
    .B1(net320),
    .B2(\reg_module.gprf[578] ),
    .X(_05013_));
 sky130_fd_sc_hd__and2_1 _10679_ (.A(net1090),
    .B(_05013_),
    .X(_00680_));
 sky130_fd_sc_hd__a32o_1 _10680_ (.A1(net415),
    .A2(net747),
    .A3(net440),
    .B1(net320),
    .B2(\reg_module.gprf[579] ),
    .X(_05014_));
 sky130_fd_sc_hd__and2_1 _10681_ (.A(net1083),
    .B(_05014_),
    .X(_00681_));
 sky130_fd_sc_hd__a32o_1 _10682_ (.A1(net414),
    .A2(net748),
    .A3(net457),
    .B1(net321),
    .B2(\reg_module.gprf[580] ),
    .X(_05015_));
 sky130_fd_sc_hd__and2_1 _10683_ (.A(net1125),
    .B(_05015_),
    .X(_00682_));
 sky130_fd_sc_hd__a32o_1 _10684_ (.A1(_04191_),
    .A2(net745),
    .A3(net437),
    .B1(net320),
    .B2(\reg_module.gprf[581] ),
    .X(_05016_));
 sky130_fd_sc_hd__and2_1 _10685_ (.A(net1086),
    .B(_05016_),
    .X(_00683_));
 sky130_fd_sc_hd__a32o_1 _10686_ (.A1(net412),
    .A2(net745),
    .A3(net433),
    .B1(net320),
    .B2(\reg_module.gprf[582] ),
    .X(_05017_));
 sky130_fd_sc_hd__and2_1 _10687_ (.A(net1079),
    .B(_05017_),
    .X(_00684_));
 sky130_fd_sc_hd__a32o_1 _10688_ (.A1(net411),
    .A2(net747),
    .A3(net440),
    .B1(net320),
    .B2(\reg_module.gprf[583] ),
    .X(_05018_));
 sky130_fd_sc_hd__and2_1 _10689_ (.A(net1087),
    .B(_05018_),
    .X(_00685_));
 sky130_fd_sc_hd__a32o_1 _10690_ (.A1(net410),
    .A2(net748),
    .A3(net454),
    .B1(net321),
    .B2(\reg_module.gprf[584] ),
    .X(_05019_));
 sky130_fd_sc_hd__and2_1 _10691_ (.A(net1125),
    .B(_05019_),
    .X(_00686_));
 sky130_fd_sc_hd__a32o_1 _10692_ (.A1(net409),
    .A2(net745),
    .A3(net434),
    .B1(net320),
    .B2(\reg_module.gprf[585] ),
    .X(_05020_));
 sky130_fd_sc_hd__and2_1 _10693_ (.A(net1078),
    .B(_05020_),
    .X(_00687_));
 sky130_fd_sc_hd__a32o_1 _10694_ (.A1(net408),
    .A2(net745),
    .A3(net434),
    .B1(net320),
    .B2(\reg_module.gprf[586] ),
    .X(_05021_));
 sky130_fd_sc_hd__and2_1 _10695_ (.A(net1077),
    .B(_05021_),
    .X(_00688_));
 sky130_fd_sc_hd__a32o_1 _10696_ (.A1(net407),
    .A2(net746),
    .A3(net444),
    .B1(net321),
    .B2(\reg_module.gprf[587] ),
    .X(_05022_));
 sky130_fd_sc_hd__and2_1 _10697_ (.A(net1098),
    .B(_05022_),
    .X(_00689_));
 sky130_fd_sc_hd__a32o_1 _10698_ (.A1(net406),
    .A2(net746),
    .A3(net446),
    .B1(net320),
    .B2(\reg_module.gprf[588] ),
    .X(_05023_));
 sky130_fd_sc_hd__and2_1 _10699_ (.A(net1104),
    .B(_05023_),
    .X(_00690_));
 sky130_fd_sc_hd__a32o_1 _10700_ (.A1(_04207_),
    .A2(net746),
    .A3(net448),
    .B1(net320),
    .B2(\reg_module.gprf[589] ),
    .X(_05024_));
 sky130_fd_sc_hd__and2_1 _10701_ (.A(net1108),
    .B(_05024_),
    .X(_00691_));
 sky130_fd_sc_hd__a32o_1 _10702_ (.A1(net404),
    .A2(_04245_),
    .A3(net459),
    .B1(net321),
    .B2(\reg_module.gprf[590] ),
    .X(_05025_));
 sky130_fd_sc_hd__and2_1 _10703_ (.A(net1115),
    .B(_05025_),
    .X(_00692_));
 sky130_fd_sc_hd__a32o_1 _10704_ (.A1(net403),
    .A2(net750),
    .A3(net465),
    .B1(net322),
    .B2(\reg_module.gprf[591] ),
    .X(_05026_));
 sky130_fd_sc_hd__and2_1 _10705_ (.A(net1156),
    .B(_05026_),
    .X(_00693_));
 sky130_fd_sc_hd__a32o_1 _10706_ (.A1(net402),
    .A2(net751),
    .A3(net487),
    .B1(net323),
    .B2(\reg_module.gprf[592] ),
    .X(_05027_));
 sky130_fd_sc_hd__and2_1 _10707_ (.A(net1189),
    .B(_05027_),
    .X(_00694_));
 sky130_fd_sc_hd__a32o_1 _10708_ (.A1(net401),
    .A2(net750),
    .A3(net463),
    .B1(net322),
    .B2(\reg_module.gprf[593] ),
    .X(_05028_));
 sky130_fd_sc_hd__and2_1 _10709_ (.A(net1148),
    .B(_05028_),
    .X(_00695_));
 sky130_fd_sc_hd__a32o_1 _10710_ (.A1(net400),
    .A2(net750),
    .A3(net460),
    .B1(net322),
    .B2(\reg_module.gprf[594] ),
    .X(_05029_));
 sky130_fd_sc_hd__and2_1 _10711_ (.A(net1143),
    .B(_05029_),
    .X(_00696_));
 sky130_fd_sc_hd__a32o_1 _10712_ (.A1(net399),
    .A2(net750),
    .A3(net460),
    .B1(net322),
    .B2(\reg_module.gprf[595] ),
    .X(_05030_));
 sky130_fd_sc_hd__and2_1 _10713_ (.A(net1144),
    .B(_05030_),
    .X(_00697_));
 sky130_fd_sc_hd__a32o_1 _10714_ (.A1(net398),
    .A2(net746),
    .A3(net450),
    .B1(net321),
    .B2(\reg_module.gprf[596] ),
    .X(_05031_));
 sky130_fd_sc_hd__and2_1 _10715_ (.A(net1115),
    .B(_05031_),
    .X(_00698_));
 sky130_fd_sc_hd__a32o_1 _10716_ (.A1(net397),
    .A2(net751),
    .A3(net484),
    .B1(net323),
    .B2(\reg_module.gprf[597] ),
    .X(_05032_));
 sky130_fd_sc_hd__and2_1 _10717_ (.A(net1201),
    .B(_05032_),
    .X(_00699_));
 sky130_fd_sc_hd__a32o_1 _10718_ (.A1(net396),
    .A2(net751),
    .A3(net482),
    .B1(net323),
    .B2(\reg_module.gprf[598] ),
    .X(_05033_));
 sky130_fd_sc_hd__and2_1 _10719_ (.A(net1191),
    .B(_05033_),
    .X(_00700_));
 sky130_fd_sc_hd__a32o_1 _10720_ (.A1(net395),
    .A2(net749),
    .A3(net470),
    .B1(net322),
    .B2(\reg_module.gprf[599] ),
    .X(_05034_));
 sky130_fd_sc_hd__and2_1 _10721_ (.A(net1169),
    .B(_05034_),
    .X(_00701_));
 sky130_fd_sc_hd__a32o_1 _10722_ (.A1(net394),
    .A2(net752),
    .A3(net476),
    .B1(net322),
    .B2(\reg_module.gprf[600] ),
    .X(_05035_));
 sky130_fd_sc_hd__and2_1 _10723_ (.A(net1176),
    .B(_05035_),
    .X(_00702_));
 sky130_fd_sc_hd__a32o_1 _10724_ (.A1(net393),
    .A2(net749),
    .A3(net475),
    .B1(net322),
    .B2(\reg_module.gprf[601] ),
    .X(_05036_));
 sky130_fd_sc_hd__and2_1 _10725_ (.A(net1176),
    .B(_05036_),
    .X(_00703_));
 sky130_fd_sc_hd__a32o_1 _10726_ (.A1(net392),
    .A2(net751),
    .A3(net487),
    .B1(net322),
    .B2(\reg_module.gprf[602] ),
    .X(_05037_));
 sky130_fd_sc_hd__and2_1 _10727_ (.A(net1161),
    .B(_05037_),
    .X(_00704_));
 sky130_fd_sc_hd__a32o_1 _10728_ (.A1(net391),
    .A2(net749),
    .A3(net470),
    .B1(net322),
    .B2(\reg_module.gprf[603] ),
    .X(_05038_));
 sky130_fd_sc_hd__and2_1 _10729_ (.A(net1149),
    .B(_05038_),
    .X(_00705_));
 sky130_fd_sc_hd__a32o_1 _10730_ (.A1(net390),
    .A2(net749),
    .A3(net471),
    .B1(net322),
    .B2(\reg_module.gprf[604] ),
    .X(_05039_));
 sky130_fd_sc_hd__and2_1 _10731_ (.A(net1168),
    .B(_05039_),
    .X(_00706_));
 sky130_fd_sc_hd__a32o_1 _10732_ (.A1(_04239_),
    .A2(net752),
    .A3(net475),
    .B1(net323),
    .B2(\reg_module.gprf[605] ),
    .X(_05040_));
 sky130_fd_sc_hd__and2_1 _10733_ (.A(net1176),
    .B(_05040_),
    .X(_00707_));
 sky130_fd_sc_hd__a32o_1 _10734_ (.A1(net388),
    .A2(net751),
    .A3(net482),
    .B1(net323),
    .B2(\reg_module.gprf[606] ),
    .X(_05041_));
 sky130_fd_sc_hd__and2_1 _10735_ (.A(net1190),
    .B(_05041_),
    .X(_00708_));
 sky130_fd_sc_hd__a32o_1 _10736_ (.A1(_04243_),
    .A2(net752),
    .A3(net483),
    .B1(net323),
    .B2(\reg_module.gprf[607] ),
    .X(_05042_));
 sky130_fd_sc_hd__and2_1 _10737_ (.A(net1199),
    .B(_05042_),
    .X(_00709_));
 sky130_fd_sc_hd__nand3_4 _10738_ (.A(net965),
    .B(net666),
    .C(net453),
    .Y(_05043_));
 sky130_fd_sc_hd__a32o_1 _10739_ (.A1(net418),
    .A2(net665),
    .A3(net459),
    .B1(net316),
    .B2(\reg_module.gprf[608] ),
    .X(_05044_));
 sky130_fd_sc_hd__and2_1 _10740_ (.A(net1111),
    .B(_05044_),
    .X(_00710_));
 sky130_fd_sc_hd__a32o_1 _10741_ (.A1(_04183_),
    .A2(net666),
    .A3(net458),
    .B1(net317),
    .B2(\reg_module.gprf[609] ),
    .X(_05045_));
 sky130_fd_sc_hd__and2_1 _10742_ (.A(net1132),
    .B(_05045_),
    .X(_00711_));
 sky130_fd_sc_hd__a32o_1 _10743_ (.A1(net416),
    .A2(net663),
    .A3(net447),
    .B1(net316),
    .B2(\reg_module.gprf[610] ),
    .X(_05046_));
 sky130_fd_sc_hd__and2_1 _10744_ (.A(net1107),
    .B(_05046_),
    .X(_00712_));
 sky130_fd_sc_hd__a32o_1 _10745_ (.A1(_04187_),
    .A2(net665),
    .A3(net440),
    .B1(net316),
    .B2(\reg_module.gprf[611] ),
    .X(_05047_));
 sky130_fd_sc_hd__and2_1 _10746_ (.A(net1092),
    .B(_05047_),
    .X(_00713_));
 sky130_fd_sc_hd__a32o_1 _10747_ (.A1(net414),
    .A2(net666),
    .A3(net457),
    .B1(net317),
    .B2(\reg_module.gprf[612] ),
    .X(_05048_));
 sky130_fd_sc_hd__and2_1 _10748_ (.A(net1133),
    .B(_05048_),
    .X(_00714_));
 sky130_fd_sc_hd__a32o_1 _10749_ (.A1(net413),
    .A2(net665),
    .A3(net438),
    .B1(net316),
    .B2(\reg_module.gprf[613] ),
    .X(_05049_));
 sky130_fd_sc_hd__and2_1 _10750_ (.A(net1091),
    .B(_05049_),
    .X(_00715_));
 sky130_fd_sc_hd__a32o_1 _10751_ (.A1(_04193_),
    .A2(net663),
    .A3(net434),
    .B1(net316),
    .B2(\reg_module.gprf[614] ),
    .X(_05050_));
 sky130_fd_sc_hd__and2_1 _10752_ (.A(net1079),
    .B(_05050_),
    .X(_00716_));
 sky130_fd_sc_hd__a32o_1 _10753_ (.A1(net411),
    .A2(net663),
    .A3(net441),
    .B1(net316),
    .B2(\reg_module.gprf[615] ),
    .X(_05051_));
 sky130_fd_sc_hd__and2_1 _10754_ (.A(net1089),
    .B(_05051_),
    .X(_00717_));
 sky130_fd_sc_hd__a32o_1 _10755_ (.A1(net410),
    .A2(net666),
    .A3(net453),
    .B1(net317),
    .B2(\reg_module.gprf[616] ),
    .X(_05052_));
 sky130_fd_sc_hd__and2_1 _10756_ (.A(net1124),
    .B(_05052_),
    .X(_00718_));
 sky130_fd_sc_hd__a32o_1 _10757_ (.A1(net409),
    .A2(net663),
    .A3(net436),
    .B1(net316),
    .B2(\reg_module.gprf[617] ),
    .X(_05053_));
 sky130_fd_sc_hd__and2_1 _10758_ (.A(net1078),
    .B(_05053_),
    .X(_00719_));
 sky130_fd_sc_hd__a32o_1 _10759_ (.A1(net408),
    .A2(net663),
    .A3(net434),
    .B1(net316),
    .B2(\reg_module.gprf[618] ),
    .X(_05054_));
 sky130_fd_sc_hd__and2_1 _10760_ (.A(net1077),
    .B(_05054_),
    .X(_00720_));
 sky130_fd_sc_hd__a32o_1 _10761_ (.A1(net407),
    .A2(net664),
    .A3(net446),
    .B1(net317),
    .B2(\reg_module.gprf[619] ),
    .X(_05055_));
 sky130_fd_sc_hd__and2_1 _10762_ (.A(net1102),
    .B(_05055_),
    .X(_00721_));
 sky130_fd_sc_hd__a32o_1 _10763_ (.A1(net406),
    .A2(net664),
    .A3(net446),
    .B1(net316),
    .B2(\reg_module.gprf[620] ),
    .X(_05056_));
 sky130_fd_sc_hd__and2_1 _10764_ (.A(net1104),
    .B(_05056_),
    .X(_00722_));
 sky130_fd_sc_hd__a32o_1 _10765_ (.A1(net405),
    .A2(net664),
    .A3(net448),
    .B1(net316),
    .B2(\reg_module.gprf[621] ),
    .X(_05057_));
 sky130_fd_sc_hd__and2_1 _10766_ (.A(net1108),
    .B(_05057_),
    .X(_00723_));
 sky130_fd_sc_hd__a32o_1 _10767_ (.A1(net404),
    .A2(net665),
    .A3(net450),
    .B1(net317),
    .B2(\reg_module.gprf[622] ),
    .X(_05058_));
 sky130_fd_sc_hd__and2_1 _10768_ (.A(net1115),
    .B(_05058_),
    .X(_00724_));
 sky130_fd_sc_hd__a32o_1 _10769_ (.A1(net403),
    .A2(net668),
    .A3(net465),
    .B1(net318),
    .B2(\reg_module.gprf[623] ),
    .X(_05059_));
 sky130_fd_sc_hd__and2_1 _10770_ (.A(net1156),
    .B(_05059_),
    .X(_00725_));
 sky130_fd_sc_hd__a32o_1 _10771_ (.A1(net402),
    .A2(net669),
    .A3(net484),
    .B1(net319),
    .B2(\reg_module.gprf[624] ),
    .X(_05060_));
 sky130_fd_sc_hd__and2_1 _10772_ (.A(net1202),
    .B(_05060_),
    .X(_00726_));
 sky130_fd_sc_hd__a32o_1 _10773_ (.A1(_04215_),
    .A2(net668),
    .A3(net463),
    .B1(net318),
    .B2(\reg_module.gprf[625] ),
    .X(_05061_));
 sky130_fd_sc_hd__and2_1 _10774_ (.A(net1148),
    .B(_05061_),
    .X(_00727_));
 sky130_fd_sc_hd__a32o_1 _10775_ (.A1(_04217_),
    .A2(net668),
    .A3(net460),
    .B1(net318),
    .B2(\reg_module.gprf[626] ),
    .X(_05062_));
 sky130_fd_sc_hd__and2_1 _10776_ (.A(net1143),
    .B(_05062_),
    .X(_00728_));
 sky130_fd_sc_hd__a32o_1 _10777_ (.A1(net399),
    .A2(net668),
    .A3(net463),
    .B1(net318),
    .B2(\reg_module.gprf[627] ),
    .X(_05063_));
 sky130_fd_sc_hd__and2_1 _10778_ (.A(net1148),
    .B(_05063_),
    .X(_00729_));
 sky130_fd_sc_hd__a32o_1 _10779_ (.A1(net398),
    .A2(net664),
    .A3(net449),
    .B1(net317),
    .B2(\reg_module.gprf[628] ),
    .X(_05064_));
 sky130_fd_sc_hd__and2_1 _10780_ (.A(net1113),
    .B(_05064_),
    .X(_00730_));
 sky130_fd_sc_hd__a32o_1 _10781_ (.A1(net397),
    .A2(net669),
    .A3(net486),
    .B1(net319),
    .B2(\reg_module.gprf[629] ),
    .X(_05065_));
 sky130_fd_sc_hd__and2_1 _10782_ (.A(net1207),
    .B(_05065_),
    .X(_00731_));
 sky130_fd_sc_hd__a32o_1 _10783_ (.A1(net396),
    .A2(net669),
    .A3(net481),
    .B1(net319),
    .B2(\reg_module.gprf[630] ),
    .X(_05066_));
 sky130_fd_sc_hd__and2_1 _10784_ (.A(net1191),
    .B(_05066_),
    .X(_00732_));
 sky130_fd_sc_hd__a32o_1 _10785_ (.A1(net395),
    .A2(net667),
    .A3(net470),
    .B1(net318),
    .B2(\reg_module.gprf[631] ),
    .X(_05067_));
 sky130_fd_sc_hd__and2_1 _10786_ (.A(net1169),
    .B(_05067_),
    .X(_00733_));
 sky130_fd_sc_hd__a32o_1 _10787_ (.A1(net394),
    .A2(net670),
    .A3(net477),
    .B1(net318),
    .B2(\reg_module.gprf[632] ),
    .X(_05068_));
 sky130_fd_sc_hd__and2_1 _10788_ (.A(net1179),
    .B(_05068_),
    .X(_00734_));
 sky130_fd_sc_hd__a32o_1 _10789_ (.A1(_04231_),
    .A2(net670),
    .A3(net477),
    .B1(net318),
    .B2(\reg_module.gprf[633] ),
    .X(_05069_));
 sky130_fd_sc_hd__and2_1 _10790_ (.A(net1176),
    .B(_05069_),
    .X(_00735_));
 sky130_fd_sc_hd__a32o_1 _10791_ (.A1(net392),
    .A2(net669),
    .A3(net487),
    .B1(net318),
    .B2(\reg_module.gprf[634] ),
    .X(_05070_));
 sky130_fd_sc_hd__and2_1 _10792_ (.A(net1161),
    .B(_05070_),
    .X(_00736_));
 sky130_fd_sc_hd__a32o_1 _10793_ (.A1(_04235_),
    .A2(net667),
    .A3(net470),
    .B1(net318),
    .B2(\reg_module.gprf[635] ),
    .X(_05071_));
 sky130_fd_sc_hd__and2_1 _10794_ (.A(net1167),
    .B(_05071_),
    .X(_00737_));
 sky130_fd_sc_hd__a32o_1 _10795_ (.A1(net390),
    .A2(net667),
    .A3(net473),
    .B1(net319),
    .B2(\reg_module.gprf[636] ),
    .X(_05072_));
 sky130_fd_sc_hd__and2_1 _10796_ (.A(net1171),
    .B(_05072_),
    .X(_00738_));
 sky130_fd_sc_hd__a32o_1 _10797_ (.A1(net389),
    .A2(net667),
    .A3(net475),
    .B1(net319),
    .B2(\reg_module.gprf[637] ),
    .X(_05073_));
 sky130_fd_sc_hd__and2_1 _10798_ (.A(net1176),
    .B(_05073_),
    .X(_00739_));
 sky130_fd_sc_hd__a32o_1 _10799_ (.A1(net388),
    .A2(net669),
    .A3(net482),
    .B1(net318),
    .B2(\reg_module.gprf[638] ),
    .X(_05074_));
 sky130_fd_sc_hd__and2_1 _10800_ (.A(net1190),
    .B(_05074_),
    .X(_00740_));
 sky130_fd_sc_hd__a32o_1 _10801_ (.A1(_04243_),
    .A2(net670),
    .A3(net485),
    .B1(net319),
    .B2(\reg_module.gprf[639] ),
    .X(_05075_));
 sky130_fd_sc_hd__and2_1 _10802_ (.A(net1199),
    .B(_05075_),
    .X(_00741_));
 sky130_fd_sc_hd__nand3_4 _10803_ (.A(net967),
    .B(net658),
    .C(net457),
    .Y(_05076_));
 sky130_fd_sc_hd__a32o_1 _10804_ (.A1(net418),
    .A2(net657),
    .A3(net441),
    .B1(net312),
    .B2(\reg_module.gprf[640] ),
    .X(_05077_));
 sky130_fd_sc_hd__and2_1 _10805_ (.A(net1091),
    .B(_05077_),
    .X(_00742_));
 sky130_fd_sc_hd__a32o_1 _10806_ (.A1(_04183_),
    .A2(net658),
    .A3(net457),
    .B1(net313),
    .B2(\reg_module.gprf[641] ),
    .X(_05078_));
 sky130_fd_sc_hd__and2_1 _10807_ (.A(net1133),
    .B(_05078_),
    .X(_00743_));
 sky130_fd_sc_hd__a32o_1 _10808_ (.A1(net416),
    .A2(net657),
    .A3(net440),
    .B1(net312),
    .B2(\reg_module.gprf[642] ),
    .X(_05079_));
 sky130_fd_sc_hd__and2_1 _10809_ (.A(net1088),
    .B(_05079_),
    .X(_00744_));
 sky130_fd_sc_hd__a32o_1 _10810_ (.A1(net415),
    .A2(net655),
    .A3(net439),
    .B1(net312),
    .B2(\reg_module.gprf[643] ),
    .X(_05080_));
 sky130_fd_sc_hd__and2_1 _10811_ (.A(net1082),
    .B(_05080_),
    .X(_00745_));
 sky130_fd_sc_hd__a32o_1 _10812_ (.A1(net414),
    .A2(net658),
    .A3(net456),
    .B1(net313),
    .B2(\reg_module.gprf[644] ),
    .X(_05081_));
 sky130_fd_sc_hd__and2_1 _10813_ (.A(net1126),
    .B(_05081_),
    .X(_00746_));
 sky130_fd_sc_hd__a32o_1 _10814_ (.A1(net413),
    .A2(net655),
    .A3(net437),
    .B1(net312),
    .B2(\reg_module.gprf[645] ),
    .X(_05082_));
 sky130_fd_sc_hd__and2_1 _10815_ (.A(net1085),
    .B(_05082_),
    .X(_00747_));
 sky130_fd_sc_hd__a32o_1 _10816_ (.A1(net412),
    .A2(net655),
    .A3(net433),
    .B1(net312),
    .B2(\reg_module.gprf[646] ),
    .X(_05083_));
 sky130_fd_sc_hd__and2_1 _10817_ (.A(net1071),
    .B(_05083_),
    .X(_00748_));
 sky130_fd_sc_hd__a32o_1 _10818_ (.A1(net411),
    .A2(net655),
    .A3(net437),
    .B1(net312),
    .B2(\reg_module.gprf[647] ),
    .X(_05084_));
 sky130_fd_sc_hd__and2_1 _10819_ (.A(net1084),
    .B(_05084_),
    .X(_00749_));
 sky130_fd_sc_hd__a32o_1 _10820_ (.A1(net410),
    .A2(net658),
    .A3(net454),
    .B1(net313),
    .B2(\reg_module.gprf[648] ),
    .X(_05085_));
 sky130_fd_sc_hd__and2_1 _10821_ (.A(net1120),
    .B(_05085_),
    .X(_00750_));
 sky130_fd_sc_hd__a32o_1 _10822_ (.A1(net409),
    .A2(net655),
    .A3(net434),
    .B1(net312),
    .B2(\reg_module.gprf[649] ),
    .X(_05086_));
 sky130_fd_sc_hd__and2_1 _10823_ (.A(net1078),
    .B(_05086_),
    .X(_00751_));
 sky130_fd_sc_hd__a32o_1 _10824_ (.A1(net408),
    .A2(net655),
    .A3(net433),
    .B1(net312),
    .B2(\reg_module.gprf[650] ),
    .X(_05087_));
 sky130_fd_sc_hd__and2_1 _10825_ (.A(net1072),
    .B(_05087_),
    .X(_00752_));
 sky130_fd_sc_hd__a32o_1 _10826_ (.A1(net407),
    .A2(net656),
    .A3(net444),
    .B1(net312),
    .B2(\reg_module.gprf[651] ),
    .X(_05088_));
 sky130_fd_sc_hd__and2_1 _10827_ (.A(net1098),
    .B(_05088_),
    .X(_00753_));
 sky130_fd_sc_hd__a32o_1 _10828_ (.A1(net406),
    .A2(net656),
    .A3(net449),
    .B1(net313),
    .B2(\reg_module.gprf[652] ),
    .X(_05089_));
 sky130_fd_sc_hd__and2_1 _10829_ (.A(net1102),
    .B(_05089_),
    .X(_00754_));
 sky130_fd_sc_hd__a32o_1 _10830_ (.A1(net405),
    .A2(net656),
    .A3(net444),
    .B1(net312),
    .B2(\reg_module.gprf[653] ),
    .X(_05090_));
 sky130_fd_sc_hd__and2_1 _10831_ (.A(net1098),
    .B(_05090_),
    .X(_00755_));
 sky130_fd_sc_hd__a32o_1 _10832_ (.A1(net404),
    .A2(net656),
    .A3(net447),
    .B1(net313),
    .B2(\reg_module.gprf[654] ),
    .X(_05091_));
 sky130_fd_sc_hd__and2_1 _10833_ (.A(net1111),
    .B(_05091_),
    .X(_00756_));
 sky130_fd_sc_hd__a32o_1 _10834_ (.A1(net403),
    .A2(net661),
    .A3(net465),
    .B1(net314),
    .B2(\reg_module.gprf[655] ),
    .X(_05092_));
 sky130_fd_sc_hd__and2_1 _10835_ (.A(net1155),
    .B(_05092_),
    .X(_00757_));
 sky130_fd_sc_hd__a32o_1 _10836_ (.A1(net402),
    .A2(net662),
    .A3(net483),
    .B1(net315),
    .B2(\reg_module.gprf[656] ),
    .X(_05093_));
 sky130_fd_sc_hd__and2_1 _10837_ (.A(net1200),
    .B(_05093_),
    .X(_00758_));
 sky130_fd_sc_hd__a32o_1 _10838_ (.A1(net401),
    .A2(net659),
    .A3(net463),
    .B1(net315),
    .B2(\reg_module.gprf[657] ),
    .X(_05094_));
 sky130_fd_sc_hd__and2_1 _10839_ (.A(net1148),
    .B(_05094_),
    .X(_00759_));
 sky130_fd_sc_hd__a32o_1 _10840_ (.A1(net400),
    .A2(net659),
    .A3(net446),
    .B1(net314),
    .B2(\reg_module.gprf[658] ),
    .X(_05095_));
 sky130_fd_sc_hd__and2_1 _10841_ (.A(net1103),
    .B(_05095_),
    .X(_00760_));
 sky130_fd_sc_hd__a32o_1 _10842_ (.A1(net399),
    .A2(net659),
    .A3(net463),
    .B1(net314),
    .B2(\reg_module.gprf[659] ),
    .X(_05096_));
 sky130_fd_sc_hd__and2_1 _10843_ (.A(net1144),
    .B(_05096_),
    .X(_00761_));
 sky130_fd_sc_hd__a32o_1 _10844_ (.A1(net398),
    .A2(net657),
    .A3(net447),
    .B1(net313),
    .B2(\reg_module.gprf[660] ),
    .X(_05097_));
 sky130_fd_sc_hd__and2_1 _10845_ (.A(net1110),
    .B(_05097_),
    .X(_00762_));
 sky130_fd_sc_hd__a32o_1 _10846_ (.A1(net397),
    .A2(net662),
    .A3(net483),
    .B1(net315),
    .B2(\reg_module.gprf[661] ),
    .X(_05098_));
 sky130_fd_sc_hd__and2_1 _10847_ (.A(net1199),
    .B(_05098_),
    .X(_00763_));
 sky130_fd_sc_hd__a32o_1 _10848_ (.A1(net396),
    .A2(net662),
    .A3(net482),
    .B1(net315),
    .B2(\reg_module.gprf[662] ),
    .X(_05099_));
 sky130_fd_sc_hd__and2_1 _10849_ (.A(net1190),
    .B(_05099_),
    .X(_00764_));
 sky130_fd_sc_hd__a32o_1 _10850_ (.A1(net395),
    .A2(net660),
    .A3(net471),
    .B1(net314),
    .B2(\reg_module.gprf[663] ),
    .X(_05100_));
 sky130_fd_sc_hd__and2_1 _10851_ (.A(net1167),
    .B(_05100_),
    .X(_00765_));
 sky130_fd_sc_hd__a32o_1 _10852_ (.A1(net394),
    .A2(net660),
    .A3(net475),
    .B1(net314),
    .B2(\reg_module.gprf[664] ),
    .X(_05101_));
 sky130_fd_sc_hd__and2_1 _10853_ (.A(net1176),
    .B(_05101_),
    .X(_00766_));
 sky130_fd_sc_hd__a32o_1 _10854_ (.A1(net393),
    .A2(net660),
    .A3(net471),
    .B1(net314),
    .B2(\reg_module.gprf[665] ),
    .X(_05102_));
 sky130_fd_sc_hd__and2_1 _10855_ (.A(net1168),
    .B(_05102_),
    .X(_00767_));
 sky130_fd_sc_hd__a32o_1 _10856_ (.A1(net392),
    .A2(net659),
    .A3(net468),
    .B1(net314),
    .B2(\reg_module.gprf[666] ),
    .X(_05103_));
 sky130_fd_sc_hd__and2_1 _10857_ (.A(net1161),
    .B(_05103_),
    .X(_00768_));
 sky130_fd_sc_hd__a32o_1 _10858_ (.A1(net391),
    .A2(net659),
    .A3(net464),
    .B1(net314),
    .B2(\reg_module.gprf[667] ),
    .X(_05104_));
 sky130_fd_sc_hd__and2_1 _10859_ (.A(net1148),
    .B(_05104_),
    .X(_00769_));
 sky130_fd_sc_hd__a32o_1 _10860_ (.A1(net390),
    .A2(net660),
    .A3(net470),
    .B1(net314),
    .B2(\reg_module.gprf[668] ),
    .X(_05105_));
 sky130_fd_sc_hd__and2_1 _10861_ (.A(net1168),
    .B(_05105_),
    .X(_00770_));
 sky130_fd_sc_hd__a32o_1 _10862_ (.A1(net389),
    .A2(net660),
    .A3(net476),
    .B1(net314),
    .B2(\reg_module.gprf[669] ),
    .X(_05106_));
 sky130_fd_sc_hd__and2_1 _10863_ (.A(net1175),
    .B(_05106_),
    .X(_00771_));
 sky130_fd_sc_hd__a32o_1 _10864_ (.A1(net388),
    .A2(net661),
    .A3(net476),
    .B1(net315),
    .B2(\reg_module.gprf[670] ),
    .X(_05107_));
 sky130_fd_sc_hd__and2_1 _10865_ (.A(net1179),
    .B(_05107_),
    .X(_00772_));
 sky130_fd_sc_hd__a32o_1 _10866_ (.A1(net387),
    .A2(net662),
    .A3(net482),
    .B1(net315),
    .B2(\reg_module.gprf[671] ),
    .X(_05108_));
 sky130_fd_sc_hd__and2_1 _10867_ (.A(net1191),
    .B(_05108_),
    .X(_00773_));
 sky130_fd_sc_hd__nand3_4 _10868_ (.A(net967),
    .B(net650),
    .C(net457),
    .Y(_05109_));
 sky130_fd_sc_hd__a32o_1 _10869_ (.A1(net418),
    .A2(net647),
    .A3(net441),
    .B1(net308),
    .B2(\reg_module.gprf[672] ),
    .X(_05110_));
 sky130_fd_sc_hd__and2_1 _10870_ (.A(net1091),
    .B(_05110_),
    .X(_00774_));
 sky130_fd_sc_hd__a32o_1 _10871_ (.A1(net417),
    .A2(net650),
    .A3(net456),
    .B1(net309),
    .B2(\reg_module.gprf[673] ),
    .X(_05111_));
 sky130_fd_sc_hd__and2_1 _10872_ (.A(net1128),
    .B(_05111_),
    .X(_00775_));
 sky130_fd_sc_hd__a32o_1 _10873_ (.A1(net416),
    .A2(net649),
    .A3(net440),
    .B1(net308),
    .B2(\reg_module.gprf[674] ),
    .X(_05112_));
 sky130_fd_sc_hd__and2_1 _10874_ (.A(net1088),
    .B(_05112_),
    .X(_00776_));
 sky130_fd_sc_hd__a32o_1 _10875_ (.A1(net415),
    .A2(net647),
    .A3(net439),
    .B1(net308),
    .B2(\reg_module.gprf[675] ),
    .X(_05113_));
 sky130_fd_sc_hd__and2_1 _10876_ (.A(net1082),
    .B(_05113_),
    .X(_00777_));
 sky130_fd_sc_hd__a32o_1 _10877_ (.A1(net414),
    .A2(net650),
    .A3(net456),
    .B1(net309),
    .B2(\reg_module.gprf[676] ),
    .X(_05114_));
 sky130_fd_sc_hd__and2_1 _10878_ (.A(net1126),
    .B(_05114_),
    .X(_00778_));
 sky130_fd_sc_hd__a32o_1 _10879_ (.A1(net413),
    .A2(net650),
    .A3(net437),
    .B1(net308),
    .B2(\reg_module.gprf[677] ),
    .X(_05115_));
 sky130_fd_sc_hd__and2_1 _10880_ (.A(net1085),
    .B(_05115_),
    .X(_00779_));
 sky130_fd_sc_hd__a32o_1 _10881_ (.A1(net412),
    .A2(net647),
    .A3(net433),
    .B1(net308),
    .B2(\reg_module.gprf[678] ),
    .X(_05116_));
 sky130_fd_sc_hd__and2_1 _10882_ (.A(net1072),
    .B(_05116_),
    .X(_00780_));
 sky130_fd_sc_hd__a32o_1 _10883_ (.A1(net411),
    .A2(net647),
    .A3(net437),
    .B1(net308),
    .B2(\reg_module.gprf[679] ),
    .X(_05117_));
 sky130_fd_sc_hd__and2_1 _10884_ (.A(net1084),
    .B(_05117_),
    .X(_00781_));
 sky130_fd_sc_hd__a32o_1 _10885_ (.A1(_04197_),
    .A2(net650),
    .A3(net452),
    .B1(net309),
    .B2(\reg_module.gprf[680] ),
    .X(_05118_));
 sky130_fd_sc_hd__and2_1 _10886_ (.A(net1120),
    .B(_05118_),
    .X(_00782_));
 sky130_fd_sc_hd__a32o_1 _10887_ (.A1(net409),
    .A2(net647),
    .A3(net435),
    .B1(net308),
    .B2(\reg_module.gprf[681] ),
    .X(_05119_));
 sky130_fd_sc_hd__and2_1 _10888_ (.A(net1076),
    .B(_05119_),
    .X(_00783_));
 sky130_fd_sc_hd__a32o_1 _10889_ (.A1(net408),
    .A2(net647),
    .A3(net433),
    .B1(net308),
    .B2(\reg_module.gprf[682] ),
    .X(_05120_));
 sky130_fd_sc_hd__and2_1 _10890_ (.A(net1072),
    .B(_05120_),
    .X(_00784_));
 sky130_fd_sc_hd__a32o_1 _10891_ (.A1(net407),
    .A2(net648),
    .A3(net443),
    .B1(net309),
    .B2(\reg_module.gprf[683] ),
    .X(_05121_));
 sky130_fd_sc_hd__and2_1 _10892_ (.A(net1096),
    .B(_05121_),
    .X(_00785_));
 sky130_fd_sc_hd__a32o_1 _10893_ (.A1(net406),
    .A2(net648),
    .A3(net445),
    .B1(net309),
    .B2(\reg_module.gprf[684] ),
    .X(_05122_));
 sky130_fd_sc_hd__and2_1 _10894_ (.A(net1102),
    .B(_05122_),
    .X(_00786_));
 sky130_fd_sc_hd__a32o_1 _10895_ (.A1(net405),
    .A2(net648),
    .A3(net444),
    .B1(net308),
    .B2(\reg_module.gprf[685] ),
    .X(_05123_));
 sky130_fd_sc_hd__and2_1 _10896_ (.A(net1105),
    .B(_05123_),
    .X(_00787_));
 sky130_fd_sc_hd__a32o_1 _10897_ (.A1(net404),
    .A2(net648),
    .A3(net447),
    .B1(net308),
    .B2(\reg_module.gprf[686] ),
    .X(_05124_));
 sky130_fd_sc_hd__and2_1 _10898_ (.A(net1111),
    .B(_05124_),
    .X(_00788_));
 sky130_fd_sc_hd__a32o_1 _10899_ (.A1(_04211_),
    .A2(net652),
    .A3(net465),
    .B1(net310),
    .B2(\reg_module.gprf[687] ),
    .X(_05125_));
 sky130_fd_sc_hd__and2_1 _10900_ (.A(net1157),
    .B(_05125_),
    .X(_00789_));
 sky130_fd_sc_hd__a32o_1 _10901_ (.A1(net402),
    .A2(net653),
    .A3(net483),
    .B1(net311),
    .B2(\reg_module.gprf[688] ),
    .X(_05126_));
 sky130_fd_sc_hd__and2_1 _10902_ (.A(net1189),
    .B(_05126_),
    .X(_00790_));
 sky130_fd_sc_hd__a32o_1 _10903_ (.A1(_04215_),
    .A2(net652),
    .A3(net462),
    .B1(net310),
    .B2(\reg_module.gprf[689] ),
    .X(_05127_));
 sky130_fd_sc_hd__and2_1 _10904_ (.A(net1147),
    .B(_05127_),
    .X(_00791_));
 sky130_fd_sc_hd__a32o_1 _10905_ (.A1(net400),
    .A2(net648),
    .A3(net446),
    .B1(net310),
    .B2(\reg_module.gprf[690] ),
    .X(_05128_));
 sky130_fd_sc_hd__and2_1 _10906_ (.A(net1103),
    .B(_05128_),
    .X(_00792_));
 sky130_fd_sc_hd__a32o_1 _10907_ (.A1(net399),
    .A2(net652),
    .A3(net461),
    .B1(net310),
    .B2(\reg_module.gprf[691] ),
    .X(_05129_));
 sky130_fd_sc_hd__and2_1 _10908_ (.A(net1144),
    .B(_05129_),
    .X(_00793_));
 sky130_fd_sc_hd__a32o_1 _10909_ (.A1(_04221_),
    .A2(net649),
    .A3(net447),
    .B1(net309),
    .B2(\reg_module.gprf[692] ),
    .X(_05130_));
 sky130_fd_sc_hd__and2_1 _10910_ (.A(net1110),
    .B(_05130_),
    .X(_00794_));
 sky130_fd_sc_hd__a32o_1 _10911_ (.A1(net397),
    .A2(net654),
    .A3(net483),
    .B1(net311),
    .B2(\reg_module.gprf[693] ),
    .X(_05131_));
 sky130_fd_sc_hd__and2_1 _10912_ (.A(net1199),
    .B(_05131_),
    .X(_00795_));
 sky130_fd_sc_hd__a32o_1 _10913_ (.A1(net396),
    .A2(net653),
    .A3(net482),
    .B1(net311),
    .B2(\reg_module.gprf[694] ),
    .X(_05132_));
 sky130_fd_sc_hd__and2_1 _10914_ (.A(net1191),
    .B(_05132_),
    .X(_00796_));
 sky130_fd_sc_hd__a32o_1 _10915_ (.A1(_04227_),
    .A2(net651),
    .A3(net470),
    .B1(net310),
    .B2(\reg_module.gprf[695] ),
    .X(_05133_));
 sky130_fd_sc_hd__and2_1 _10916_ (.A(net1167),
    .B(_05133_),
    .X(_00797_));
 sky130_fd_sc_hd__a32o_1 _10917_ (.A1(net394),
    .A2(net651),
    .A3(net475),
    .B1(net310),
    .B2(\reg_module.gprf[696] ),
    .X(_05134_));
 sky130_fd_sc_hd__and2_1 _10918_ (.A(net1176),
    .B(_05134_),
    .X(_00798_));
 sky130_fd_sc_hd__a32o_1 _10919_ (.A1(net393),
    .A2(net651),
    .A3(net471),
    .B1(net310),
    .B2(\reg_module.gprf[697] ),
    .X(_05135_));
 sky130_fd_sc_hd__and2_1 _10920_ (.A(net1168),
    .B(_05135_),
    .X(_00799_));
 sky130_fd_sc_hd__a32o_1 _10921_ (.A1(_04233_),
    .A2(net652),
    .A3(net468),
    .B1(net310),
    .B2(\reg_module.gprf[698] ),
    .X(_05136_));
 sky130_fd_sc_hd__and2_1 _10922_ (.A(net1162),
    .B(_05136_),
    .X(_00800_));
 sky130_fd_sc_hd__a32o_1 _10923_ (.A1(net391),
    .A2(net652),
    .A3(net464),
    .B1(net310),
    .B2(\reg_module.gprf[699] ),
    .X(_05137_));
 sky130_fd_sc_hd__and2_1 _10924_ (.A(net1148),
    .B(_05137_),
    .X(_00801_));
 sky130_fd_sc_hd__a32o_1 _10925_ (.A1(net390),
    .A2(net651),
    .A3(net472),
    .B1(net310),
    .B2(\reg_module.gprf[700] ),
    .X(_05138_));
 sky130_fd_sc_hd__and2_1 _10926_ (.A(net1166),
    .B(_05138_),
    .X(_00802_));
 sky130_fd_sc_hd__a32o_1 _10927_ (.A1(net389),
    .A2(net651),
    .A3(net470),
    .B1(net311),
    .B2(\reg_module.gprf[701] ),
    .X(_05139_));
 sky130_fd_sc_hd__and2_1 _10928_ (.A(net1169),
    .B(_05139_),
    .X(_00803_));
 sky130_fd_sc_hd__a32o_1 _10929_ (.A1(net388),
    .A2(net653),
    .A3(net476),
    .B1(net311),
    .B2(\reg_module.gprf[702] ),
    .X(_05140_));
 sky130_fd_sc_hd__and2_1 _10930_ (.A(net1179),
    .B(_05140_),
    .X(_00804_));
 sky130_fd_sc_hd__a32o_1 _10931_ (.A1(net387),
    .A2(net653),
    .A3(net482),
    .B1(net311),
    .B2(\reg_module.gprf[703] ),
    .X(_05141_));
 sky130_fd_sc_hd__and2_1 _10932_ (.A(net1191),
    .B(_05141_),
    .X(_00805_));
 sky130_fd_sc_hd__or2_2 _10933_ (.A(net644),
    .B(_04976_),
    .X(_05142_));
 sky130_fd_sc_hd__a22o_1 _10934_ (.A1(_04383_),
    .A2(net441),
    .B1(net304),
    .B2(\reg_module.gprf[704] ),
    .X(_05143_));
 sky130_fd_sc_hd__and2_1 _10935_ (.A(net1090),
    .B(_05143_),
    .X(_00806_));
 sky130_fd_sc_hd__a22o_1 _10936_ (.A1(_04385_),
    .A2(net455),
    .B1(net305),
    .B2(\reg_module.gprf[705] ),
    .X(_05144_));
 sky130_fd_sc_hd__and2_1 _10937_ (.A(net1128),
    .B(_05144_),
    .X(_00807_));
 sky130_fd_sc_hd__a22o_1 _10938_ (.A1(_04387_),
    .A2(net448),
    .B1(net304),
    .B2(\reg_module.gprf[706] ),
    .X(_05145_));
 sky130_fd_sc_hd__and2_1 _10939_ (.A(net1107),
    .B(_05145_),
    .X(_00808_));
 sky130_fd_sc_hd__a22o_1 _10940_ (.A1(_04389_),
    .A2(net440),
    .B1(net304),
    .B2(\reg_module.gprf[707] ),
    .X(_05146_));
 sky130_fd_sc_hd__and2_1 _10941_ (.A(net1087),
    .B(_05146_),
    .X(_00809_));
 sky130_fd_sc_hd__a22o_1 _10942_ (.A1(_04391_),
    .A2(net456),
    .B1(net305),
    .B2(\reg_module.gprf[708] ),
    .X(_05147_));
 sky130_fd_sc_hd__and2_1 _10943_ (.A(net1131),
    .B(_05147_),
    .X(_00810_));
 sky130_fd_sc_hd__a22o_1 _10944_ (.A1(_04393_),
    .A2(net452),
    .B1(net305),
    .B2(\reg_module.gprf[709] ),
    .X(_05148_));
 sky130_fd_sc_hd__and2_1 _10945_ (.A(net1086),
    .B(_05148_),
    .X(_00811_));
 sky130_fd_sc_hd__a22o_1 _10946_ (.A1(_04395_),
    .A2(net436),
    .B1(net304),
    .B2(\reg_module.gprf[710] ),
    .X(_05149_));
 sky130_fd_sc_hd__and2_1 _10947_ (.A(net1072),
    .B(_05149_),
    .X(_00812_));
 sky130_fd_sc_hd__a22o_1 _10948_ (.A1(_04397_),
    .A2(net437),
    .B1(net304),
    .B2(\reg_module.gprf[711] ),
    .X(_05150_));
 sky130_fd_sc_hd__and2_1 _10949_ (.A(net1083),
    .B(_05150_),
    .X(_00813_));
 sky130_fd_sc_hd__a22o_1 _10950_ (.A1(_04399_),
    .A2(net454),
    .B1(net305),
    .B2(\reg_module.gprf[712] ),
    .X(_05151_));
 sky130_fd_sc_hd__and2_1 _10951_ (.A(net1123),
    .B(_05151_),
    .X(_00814_));
 sky130_fd_sc_hd__a22o_1 _10952_ (.A1(_04401_),
    .A2(net435),
    .B1(net304),
    .B2(\reg_module.gprf[713] ),
    .X(_05152_));
 sky130_fd_sc_hd__and2_1 _10953_ (.A(net1076),
    .B(_05152_),
    .X(_00815_));
 sky130_fd_sc_hd__a22o_1 _10954_ (.A1(_04403_),
    .A2(net433),
    .B1(net304),
    .B2(\reg_module.gprf[714] ),
    .X(_05153_));
 sky130_fd_sc_hd__and2_1 _10955_ (.A(net1093),
    .B(_05153_),
    .X(_00816_));
 sky130_fd_sc_hd__a22o_1 _10956_ (.A1(_04405_),
    .A2(net445),
    .B1(net304),
    .B2(\reg_module.gprf[715] ),
    .X(_05154_));
 sky130_fd_sc_hd__and2_1 _10957_ (.A(net1100),
    .B(_05154_),
    .X(_00817_));
 sky130_fd_sc_hd__a22o_1 _10958_ (.A1(_04407_),
    .A2(net445),
    .B1(net305),
    .B2(\reg_module.gprf[716] ),
    .X(_05155_));
 sky130_fd_sc_hd__and2_1 _10959_ (.A(net1104),
    .B(_05155_),
    .X(_00818_));
 sky130_fd_sc_hd__a22o_1 _10960_ (.A1(_04409_),
    .A2(net444),
    .B1(net304),
    .B2(\reg_module.gprf[717] ),
    .X(_05156_));
 sky130_fd_sc_hd__and2_1 _10961_ (.A(net1105),
    .B(_05156_),
    .X(_00819_));
 sky130_fd_sc_hd__a22o_1 _10962_ (.A1(_04411_),
    .A2(net450),
    .B1(net304),
    .B2(\reg_module.gprf[718] ),
    .X(_05157_));
 sky130_fd_sc_hd__and2_1 _10963_ (.A(net1116),
    .B(_05157_),
    .X(_00820_));
 sky130_fd_sc_hd__a22o_1 _10964_ (.A1(_04413_),
    .A2(net465),
    .B1(net306),
    .B2(\reg_module.gprf[719] ),
    .X(_05158_));
 sky130_fd_sc_hd__and2_1 _10965_ (.A(net1155),
    .B(_05158_),
    .X(_00821_));
 sky130_fd_sc_hd__a22o_1 _10966_ (.A1(_04415_),
    .A2(net483),
    .B1(net307),
    .B2(\reg_module.gprf[720] ),
    .X(_05159_));
 sky130_fd_sc_hd__and2_1 _10967_ (.A(net1200),
    .B(_05159_),
    .X(_00822_));
 sky130_fd_sc_hd__a22o_1 _10968_ (.A1(_04417_),
    .A2(net460),
    .B1(net306),
    .B2(\reg_module.gprf[721] ),
    .X(_05160_));
 sky130_fd_sc_hd__and2_1 _10969_ (.A(net1142),
    .B(_05160_),
    .X(_00823_));
 sky130_fd_sc_hd__a22o_1 _10970_ (.A1(_04419_),
    .A2(net445),
    .B1(net306),
    .B2(\reg_module.gprf[722] ),
    .X(_05161_));
 sky130_fd_sc_hd__and2_1 _10971_ (.A(net1103),
    .B(_05161_),
    .X(_00824_));
 sky130_fd_sc_hd__a22o_1 _10972_ (.A1(_04421_),
    .A2(net463),
    .B1(net306),
    .B2(\reg_module.gprf[723] ),
    .X(_05162_));
 sky130_fd_sc_hd__and2_1 _10973_ (.A(net1150),
    .B(_05162_),
    .X(_00825_));
 sky130_fd_sc_hd__a22o_1 _10974_ (.A1(_04423_),
    .A2(net449),
    .B1(net305),
    .B2(\reg_module.gprf[724] ),
    .X(_05163_));
 sky130_fd_sc_hd__and2_1 _10975_ (.A(net1113),
    .B(_05163_),
    .X(_00826_));
 sky130_fd_sc_hd__a22o_1 _10976_ (.A1(_04425_),
    .A2(net485),
    .B1(net307),
    .B2(\reg_module.gprf[725] ),
    .X(_05164_));
 sky130_fd_sc_hd__and2_1 _10977_ (.A(net1200),
    .B(_05164_),
    .X(_00827_));
 sky130_fd_sc_hd__a22o_1 _10978_ (.A1(_04427_),
    .A2(net480),
    .B1(net307),
    .B2(\reg_module.gprf[726] ),
    .X(_05165_));
 sky130_fd_sc_hd__and2_1 _10979_ (.A(net1194),
    .B(_05165_),
    .X(_00828_));
 sky130_fd_sc_hd__a22o_1 _10980_ (.A1(_04429_),
    .A2(net471),
    .B1(net306),
    .B2(\reg_module.gprf[727] ),
    .X(_05166_));
 sky130_fd_sc_hd__and2_1 _10981_ (.A(net1168),
    .B(_05166_),
    .X(_00829_));
 sky130_fd_sc_hd__a22o_1 _10982_ (.A1(_04431_),
    .A2(net477),
    .B1(net306),
    .B2(\reg_module.gprf[728] ),
    .X(_05167_));
 sky130_fd_sc_hd__and2_1 _10983_ (.A(net1181),
    .B(_05167_),
    .X(_00830_));
 sky130_fd_sc_hd__a22o_1 _10984_ (.A1(_04433_),
    .A2(net473),
    .B1(net306),
    .B2(\reg_module.gprf[729] ),
    .X(_05168_));
 sky130_fd_sc_hd__and2_1 _10985_ (.A(net1173),
    .B(_05168_),
    .X(_00831_));
 sky130_fd_sc_hd__a22o_1 _10986_ (.A1(_04435_),
    .A2(net467),
    .B1(net306),
    .B2(\reg_module.gprf[730] ),
    .X(_05169_));
 sky130_fd_sc_hd__and2_1 _10987_ (.A(net1162),
    .B(_05169_),
    .X(_00832_));
 sky130_fd_sc_hd__a22o_1 _10988_ (.A1(_04437_),
    .A2(net463),
    .B1(net306),
    .B2(\reg_module.gprf[731] ),
    .X(_05170_));
 sky130_fd_sc_hd__and2_1 _10989_ (.A(net1149),
    .B(_05170_),
    .X(_00833_));
 sky130_fd_sc_hd__a22o_1 _10990_ (.A1(_04439_),
    .A2(net474),
    .B1(net307),
    .B2(\reg_module.gprf[732] ),
    .X(_05171_));
 sky130_fd_sc_hd__and2_1 _10991_ (.A(net1171),
    .B(_05171_),
    .X(_00834_));
 sky130_fd_sc_hd__a22o_1 _10992_ (.A1(_04441_),
    .A2(net475),
    .B1(net307),
    .B2(\reg_module.gprf[733] ),
    .X(_05172_));
 sky130_fd_sc_hd__and2_1 _10993_ (.A(net1175),
    .B(_05172_),
    .X(_00835_));
 sky130_fd_sc_hd__a22o_1 _10994_ (.A1(_04443_),
    .A2(net477),
    .B1(net306),
    .B2(\reg_module.gprf[734] ),
    .X(_05173_));
 sky130_fd_sc_hd__and2_1 _10995_ (.A(net1184),
    .B(_05173_),
    .X(_00836_));
 sky130_fd_sc_hd__a22o_1 _10996_ (.A1(_04445_),
    .A2(net481),
    .B1(net307),
    .B2(\reg_module.gprf[735] ),
    .X(_05174_));
 sky130_fd_sc_hd__and2_1 _10997_ (.A(net1195),
    .B(_05174_),
    .X(_00837_));
 sky130_fd_sc_hd__nand3_4 _10998_ (.A(net967),
    .B(net777),
    .C(net457),
    .Y(_05175_));
 sky130_fd_sc_hd__a32o_1 _10999_ (.A1(net776),
    .A2(net418),
    .A3(net447),
    .B1(net300),
    .B2(\reg_module.gprf[736] ),
    .X(_05176_));
 sky130_fd_sc_hd__and2_1 _11000_ (.A(net1111),
    .B(_05176_),
    .X(_00838_));
 sky130_fd_sc_hd__a32o_1 _11001_ (.A1(net777),
    .A2(net417),
    .A3(net457),
    .B1(net301),
    .B2(\reg_module.gprf[737] ),
    .X(_05177_));
 sky130_fd_sc_hd__and2_1 _11002_ (.A(net1133),
    .B(_05177_),
    .X(_00839_));
 sky130_fd_sc_hd__a32o_1 _11003_ (.A1(net776),
    .A2(net416),
    .A3(net448),
    .B1(net300),
    .B2(\reg_module.gprf[738] ),
    .X(_05178_));
 sky130_fd_sc_hd__and2_1 _11004_ (.A(net1106),
    .B(_05178_),
    .X(_00840_));
 sky130_fd_sc_hd__a32o_1 _11005_ (.A1(net774),
    .A2(_04187_),
    .A3(net440),
    .B1(net300),
    .B2(\reg_module.gprf[739] ),
    .X(_05179_));
 sky130_fd_sc_hd__and2_1 _11006_ (.A(net1087),
    .B(_05179_),
    .X(_00841_));
 sky130_fd_sc_hd__a32o_1 _11007_ (.A1(net777),
    .A2(net414),
    .A3(net456),
    .B1(net301),
    .B2(\reg_module.gprf[740] ),
    .X(_05180_));
 sky130_fd_sc_hd__and2_1 _11008_ (.A(net1131),
    .B(_05180_),
    .X(_00842_));
 sky130_fd_sc_hd__a32o_1 _11009_ (.A1(net774),
    .A2(net413),
    .A3(net438),
    .B1(net300),
    .B2(\reg_module.gprf[741] ),
    .X(_05181_));
 sky130_fd_sc_hd__and2_1 _11010_ (.A(net1086),
    .B(_05181_),
    .X(_00843_));
 sky130_fd_sc_hd__a32o_1 _11011_ (.A1(net774),
    .A2(net412),
    .A3(net436),
    .B1(net300),
    .B2(\reg_module.gprf[742] ),
    .X(_05182_));
 sky130_fd_sc_hd__and2_1 _11012_ (.A(net1073),
    .B(_05182_),
    .X(_00844_));
 sky130_fd_sc_hd__a32o_1 _11013_ (.A1(net774),
    .A2(_04195_),
    .A3(net438),
    .B1(net300),
    .B2(\reg_module.gprf[743] ),
    .X(_05183_));
 sky130_fd_sc_hd__and2_1 _11014_ (.A(net1086),
    .B(_05183_),
    .X(_00845_));
 sky130_fd_sc_hd__a32o_1 _11015_ (.A1(net777),
    .A2(net410),
    .A3(net454),
    .B1(net301),
    .B2(\reg_module.gprf[744] ),
    .X(_05184_));
 sky130_fd_sc_hd__and2_1 _11016_ (.A(net1124),
    .B(_05184_),
    .X(_00846_));
 sky130_fd_sc_hd__a32o_1 _11017_ (.A1(net774),
    .A2(net409),
    .A3(net435),
    .B1(net300),
    .B2(\reg_module.gprf[745] ),
    .X(_05185_));
 sky130_fd_sc_hd__and2_1 _11018_ (.A(net1076),
    .B(_05185_),
    .X(_00847_));
 sky130_fd_sc_hd__a32o_1 _11019_ (.A1(net774),
    .A2(net408),
    .A3(net434),
    .B1(net300),
    .B2(\reg_module.gprf[746] ),
    .X(_05186_));
 sky130_fd_sc_hd__and2_1 _11020_ (.A(net1077),
    .B(_05186_),
    .X(_00848_));
 sky130_fd_sc_hd__a32o_1 _11021_ (.A1(net775),
    .A2(net407),
    .A3(net443),
    .B1(net300),
    .B2(\reg_module.gprf[747] ),
    .X(_05187_));
 sky130_fd_sc_hd__and2_1 _11022_ (.A(net1096),
    .B(_05187_),
    .X(_00849_));
 sky130_fd_sc_hd__a32o_1 _11023_ (.A1(net775),
    .A2(_04205_),
    .A3(net445),
    .B1(net301),
    .B2(\reg_module.gprf[748] ),
    .X(_05188_));
 sky130_fd_sc_hd__and2_1 _11024_ (.A(net1104),
    .B(_05188_),
    .X(_00850_));
 sky130_fd_sc_hd__a32o_1 _11025_ (.A1(net775),
    .A2(net405),
    .A3(net446),
    .B1(net300),
    .B2(\reg_module.gprf[749] ),
    .X(_05189_));
 sky130_fd_sc_hd__and2_1 _11026_ (.A(net1104),
    .B(_05189_),
    .X(_00851_));
 sky130_fd_sc_hd__a32o_1 _11027_ (.A1(net777),
    .A2(net404),
    .A3(net459),
    .B1(net301),
    .B2(\reg_module.gprf[750] ),
    .X(_05190_));
 sky130_fd_sc_hd__and2_1 _11028_ (.A(net1136),
    .B(_05190_),
    .X(_00852_));
 sky130_fd_sc_hd__a32o_1 _11029_ (.A1(net780),
    .A2(_04211_),
    .A3(net466),
    .B1(net302),
    .B2(\reg_module.gprf[751] ),
    .X(_05191_));
 sky130_fd_sc_hd__and2_1 _11030_ (.A(net1156),
    .B(_05191_),
    .X(_00853_));
 sky130_fd_sc_hd__a32o_1 _11031_ (.A1(net781),
    .A2(_04213_),
    .A3(net483),
    .B1(net303),
    .B2(\reg_module.gprf[752] ),
    .X(_05192_));
 sky130_fd_sc_hd__and2_1 _11032_ (.A(net1200),
    .B(_05192_),
    .X(_00854_));
 sky130_fd_sc_hd__a32o_1 _11033_ (.A1(net778),
    .A2(net401),
    .A3(net462),
    .B1(net302),
    .B2(\reg_module.gprf[753] ),
    .X(_05193_));
 sky130_fd_sc_hd__and2_1 _11034_ (.A(net1147),
    .B(_05193_),
    .X(_00855_));
 sky130_fd_sc_hd__a32o_1 _11035_ (.A1(net775),
    .A2(net400),
    .A3(net460),
    .B1(net302),
    .B2(\reg_module.gprf[754] ),
    .X(_05194_));
 sky130_fd_sc_hd__and2_1 _11036_ (.A(net1103),
    .B(_05194_),
    .X(_00856_));
 sky130_fd_sc_hd__a32o_1 _11037_ (.A1(net778),
    .A2(net399),
    .A3(net463),
    .B1(net302),
    .B2(\reg_module.gprf[755] ),
    .X(_05195_));
 sky130_fd_sc_hd__and2_1 _11038_ (.A(net1150),
    .B(_05195_),
    .X(_00857_));
 sky130_fd_sc_hd__a32o_1 _11039_ (.A1(net776),
    .A2(_04221_),
    .A3(net450),
    .B1(net301),
    .B2(\reg_module.gprf[756] ),
    .X(_05196_));
 sky130_fd_sc_hd__and2_1 _11040_ (.A(net1115),
    .B(_05196_),
    .X(_00858_));
 sky130_fd_sc_hd__a32o_1 _11041_ (.A1(net781),
    .A2(net397),
    .A3(net486),
    .B1(net303),
    .B2(\reg_module.gprf[757] ),
    .X(_05197_));
 sky130_fd_sc_hd__and2_1 _11042_ (.A(net1200),
    .B(_05197_),
    .X(_00859_));
 sky130_fd_sc_hd__a32o_1 _11043_ (.A1(net781),
    .A2(net396),
    .A3(net480),
    .B1(net303),
    .B2(\reg_module.gprf[758] ),
    .X(_05198_));
 sky130_fd_sc_hd__and2_1 _11044_ (.A(net1191),
    .B(_05198_),
    .X(_00860_));
 sky130_fd_sc_hd__a32o_1 _11045_ (.A1(net779),
    .A2(_04227_),
    .A3(net470),
    .B1(net302),
    .B2(\reg_module.gprf[759] ),
    .X(_05199_));
 sky130_fd_sc_hd__and2_1 _11046_ (.A(net1168),
    .B(_05199_),
    .X(_00861_));
 sky130_fd_sc_hd__a32o_1 _11047_ (.A1(net779),
    .A2(net394),
    .A3(net477),
    .B1(net302),
    .B2(\reg_module.gprf[760] ),
    .X(_05200_));
 sky130_fd_sc_hd__and2_1 _11048_ (.A(net1177),
    .B(_05200_),
    .X(_00862_));
 sky130_fd_sc_hd__a32o_1 _11049_ (.A1(net779),
    .A2(net393),
    .A3(net474),
    .B1(net302),
    .B2(\reg_module.gprf[761] ),
    .X(_05201_));
 sky130_fd_sc_hd__and2_1 _11050_ (.A(net1169),
    .B(_05201_),
    .X(_00863_));
 sky130_fd_sc_hd__a32o_1 _11051_ (.A1(net778),
    .A2(_04233_),
    .A3(net468),
    .B1(net302),
    .B2(\reg_module.gprf[762] ),
    .X(_05202_));
 sky130_fd_sc_hd__and2_1 _11052_ (.A(net1162),
    .B(_05202_),
    .X(_00864_));
 sky130_fd_sc_hd__a32o_1 _11053_ (.A1(net778),
    .A2(net391),
    .A3(net463),
    .B1(net302),
    .B2(\reg_module.gprf[763] ),
    .X(_05203_));
 sky130_fd_sc_hd__and2_1 _11054_ (.A(net1149),
    .B(_05203_),
    .X(_00865_));
 sky130_fd_sc_hd__a32o_1 _11055_ (.A1(net779),
    .A2(net390),
    .A3(net473),
    .B1(net303),
    .B2(\reg_module.gprf[764] ),
    .X(_05204_));
 sky130_fd_sc_hd__and2_1 _11056_ (.A(net1166),
    .B(_05204_),
    .X(_00866_));
 sky130_fd_sc_hd__a32o_1 _11057_ (.A1(net779),
    .A2(_04239_),
    .A3(net476),
    .B1(net303),
    .B2(\reg_module.gprf[765] ),
    .X(_05205_));
 sky130_fd_sc_hd__and2_1 _11058_ (.A(net1176),
    .B(_05205_),
    .X(_00867_));
 sky130_fd_sc_hd__a32o_1 _11059_ (.A1(net779),
    .A2(net388),
    .A3(net477),
    .B1(net302),
    .B2(\reg_module.gprf[766] ),
    .X(_05206_));
 sky130_fd_sc_hd__and2_1 _11060_ (.A(net1184),
    .B(_05206_),
    .X(_00868_));
 sky130_fd_sc_hd__a32o_1 _11061_ (.A1(net781),
    .A2(net387),
    .A3(net480),
    .B1(net303),
    .B2(\reg_module.gprf[767] ),
    .X(_05207_));
 sky130_fd_sc_hd__and2_1 _11062_ (.A(net1198),
    .B(_05207_),
    .X(_00869_));
 sky130_fd_sc_hd__nor2_4 _11063_ (.A(_04178_),
    .B(_04976_),
    .Y(_05208_));
 sky130_fd_sc_hd__or2_1 _11064_ (.A(\reg_module.gprf[768] ),
    .B(net295),
    .X(_05209_));
 sky130_fd_sc_hd__o311a_1 _11065_ (.A1(_02686_),
    .A2(_04178_),
    .A3(_04976_),
    .B1(_05209_),
    .C1(net1125),
    .X(_00870_));
 sky130_fd_sc_hd__nand2_1 _11066_ (.A(net721),
    .B(net295),
    .Y(_05210_));
 sky130_fd_sc_hd__o211a_1 _11067_ (.A1(net1421),
    .A2(net295),
    .B1(_05210_),
    .C1(net1129),
    .X(_00871_));
 sky130_fd_sc_hd__nand2_1 _11068_ (.A(net713),
    .B(net294),
    .Y(_05211_));
 sky130_fd_sc_hd__o211a_1 _11069_ (.A1(net1350),
    .A2(net294),
    .B1(_05211_),
    .C1(net1107),
    .X(_00872_));
 sky130_fd_sc_hd__nand2_1 _11070_ (.A(_02717_),
    .B(net294),
    .Y(_05212_));
 sky130_fd_sc_hd__o211a_1 _11071_ (.A1(net1391),
    .A2(net294),
    .B1(_05212_),
    .C1(net1088),
    .X(_00873_));
 sky130_fd_sc_hd__nand2_1 _11072_ (.A(net723),
    .B(net295),
    .Y(_05213_));
 sky130_fd_sc_hd__o211a_1 _11073_ (.A1(net1359),
    .A2(net295),
    .B1(_05213_),
    .C1(net1129),
    .X(_00874_));
 sky130_fd_sc_hd__nand2_1 _11074_ (.A(net722),
    .B(net295),
    .Y(_05214_));
 sky130_fd_sc_hd__o211a_1 _11075_ (.A1(net1429),
    .A2(net295),
    .B1(_05214_),
    .C1(net1119),
    .X(_00875_));
 sky130_fd_sc_hd__nand2_1 _11076_ (.A(net725),
    .B(net293),
    .Y(_05215_));
 sky130_fd_sc_hd__o211a_1 _11077_ (.A1(net1364),
    .A2(net293),
    .B1(_05215_),
    .C1(net1081),
    .X(_00876_));
 sky130_fd_sc_hd__nand2_1 _11078_ (.A(net724),
    .B(net293),
    .Y(_05216_));
 sky130_fd_sc_hd__o211a_1 _11079_ (.A1(net1373),
    .A2(net293),
    .B1(_05216_),
    .C1(net1085),
    .X(_00877_));
 sky130_fd_sc_hd__nand2_1 _11080_ (.A(net689),
    .B(_05208_),
    .Y(_05217_));
 sky130_fd_sc_hd__o211a_1 _11081_ (.A1(net1438),
    .A2(net295),
    .B1(_05217_),
    .C1(net1121),
    .X(_00878_));
 sky130_fd_sc_hd__nand2_1 _11082_ (.A(net690),
    .B(net293),
    .Y(_05218_));
 sky130_fd_sc_hd__o211a_1 _11083_ (.A1(net1436),
    .A2(net293),
    .B1(_05218_),
    .C1(net1075),
    .X(_00879_));
 sky130_fd_sc_hd__nand2_1 _11084_ (.A(net692),
    .B(net293),
    .Y(_05219_));
 sky130_fd_sc_hd__o211a_1 _11085_ (.A1(net1444),
    .A2(net293),
    .B1(_05219_),
    .C1(net1073),
    .X(_00880_));
 sky130_fd_sc_hd__nand2_1 _11086_ (.A(net691),
    .B(net294),
    .Y(_05220_));
 sky130_fd_sc_hd__o211a_1 _11087_ (.A1(net1443),
    .A2(net294),
    .B1(_05220_),
    .C1(net1095),
    .X(_00881_));
 sky130_fd_sc_hd__nand2_1 _11088_ (.A(net693),
    .B(net296),
    .Y(_05221_));
 sky130_fd_sc_hd__o211a_1 _11089_ (.A1(net1356),
    .A2(net296),
    .B1(_05221_),
    .C1(net1143),
    .X(_00882_));
 sky130_fd_sc_hd__nand2_1 _11090_ (.A(net694),
    .B(net293),
    .Y(_05222_));
 sky130_fd_sc_hd__o211a_1 _11091_ (.A1(net1390),
    .A2(net293),
    .B1(_05222_),
    .C1(net1078),
    .X(_00883_));
 sky130_fd_sc_hd__nand2_1 _11092_ (.A(net696),
    .B(net295),
    .Y(_05223_));
 sky130_fd_sc_hd__o211a_1 _11093_ (.A1(net1357),
    .A2(net294),
    .B1(_05223_),
    .C1(net1116),
    .X(_00884_));
 sky130_fd_sc_hd__nand2_1 _11094_ (.A(net695),
    .B(net298),
    .Y(_05224_));
 sky130_fd_sc_hd__o211a_1 _11095_ (.A1(net1427),
    .A2(net298),
    .B1(_05224_),
    .C1(net1153),
    .X(_00885_));
 sky130_fd_sc_hd__nand2_1 _11096_ (.A(_02938_),
    .B(net299),
    .Y(_05225_));
 sky130_fd_sc_hd__o211a_1 _11097_ (.A1(net1397),
    .A2(net299),
    .B1(_05225_),
    .C1(net1202),
    .X(_00886_));
 sky130_fd_sc_hd__nand2_1 _11098_ (.A(net697),
    .B(net296),
    .Y(_05226_));
 sky130_fd_sc_hd__o211a_1 _11099_ (.A1(net1370),
    .A2(net296),
    .B1(_05226_),
    .C1(net1145),
    .X(_00887_));
 sky130_fd_sc_hd__nand2_1 _11100_ (.A(net700),
    .B(net296),
    .Y(_05227_));
 sky130_fd_sc_hd__o211a_1 _11101_ (.A1(net1425),
    .A2(net296),
    .B1(_05227_),
    .C1(net1139),
    .X(_00888_));
 sky130_fd_sc_hd__nand2_1 _11102_ (.A(_02923_),
    .B(net296),
    .Y(_05228_));
 sky130_fd_sc_hd__o211a_1 _11103_ (.A1(net1416),
    .A2(net296),
    .B1(_05228_),
    .C1(net1160),
    .X(_00889_));
 sky130_fd_sc_hd__nand2_1 _11104_ (.A(net702),
    .B(net294),
    .Y(_05229_));
 sky130_fd_sc_hd__o211a_1 _11105_ (.A1(net1377),
    .A2(net294),
    .B1(_05229_),
    .C1(net1113),
    .X(_00890_));
 sky130_fd_sc_hd__nand2_1 _11106_ (.A(_02894_),
    .B(net299),
    .Y(_05230_));
 sky130_fd_sc_hd__o211a_1 _11107_ (.A1(net1354),
    .A2(net299),
    .B1(_05230_),
    .C1(net1207),
    .X(_00891_));
 sky130_fd_sc_hd__nand2_1 _11108_ (.A(_02850_),
    .B(net299),
    .Y(_05231_));
 sky130_fd_sc_hd__o211a_1 _11109_ (.A1(net1366),
    .A2(net299),
    .B1(_05231_),
    .C1(net1196),
    .X(_00892_));
 sky130_fd_sc_hd__nand2_1 _11110_ (.A(net703),
    .B(net297),
    .Y(_05232_));
 sky130_fd_sc_hd__o211a_1 _11111_ (.A1(net1410),
    .A2(net297),
    .B1(_05232_),
    .C1(net1164),
    .X(_00893_));
 sky130_fd_sc_hd__nand2_1 _11112_ (.A(_02832_),
    .B(net297),
    .Y(_05233_));
 sky130_fd_sc_hd__o211a_1 _11113_ (.A1(net1395),
    .A2(net297),
    .B1(_05233_),
    .C1(net1183),
    .X(_00894_));
 sky130_fd_sc_hd__nand2_1 _11114_ (.A(_02816_),
    .B(net297),
    .Y(_05234_));
 sky130_fd_sc_hd__o211a_1 _11115_ (.A1(net1400),
    .A2(net297),
    .B1(_05234_),
    .C1(net1172),
    .X(_00895_));
 sky130_fd_sc_hd__nand2_1 _11116_ (.A(net708),
    .B(net298),
    .Y(_05235_));
 sky130_fd_sc_hd__o211a_1 _11117_ (.A1(net1389),
    .A2(net298),
    .B1(_05235_),
    .C1(net1163),
    .X(_00896_));
 sky130_fd_sc_hd__nand2_1 _11118_ (.A(net707),
    .B(net296),
    .Y(_05236_));
 sky130_fd_sc_hd__o211a_1 _11119_ (.A1(net1437),
    .A2(net296),
    .B1(_05236_),
    .C1(net1146),
    .X(_00897_));
 sky130_fd_sc_hd__nand2_1 _11120_ (.A(net710),
    .B(net297),
    .Y(_05237_));
 sky130_fd_sc_hd__o211a_1 _11121_ (.A1(net1361),
    .A2(net297),
    .B1(_05237_),
    .C1(net1174),
    .X(_00898_));
 sky130_fd_sc_hd__nand2_1 _11122_ (.A(net709),
    .B(net298),
    .Y(_05238_));
 sky130_fd_sc_hd__o211a_1 _11123_ (.A1(net1363),
    .A2(net298),
    .B1(_05238_),
    .C1(net1177),
    .X(_00899_));
 sky130_fd_sc_hd__nand2_1 _11124_ (.A(net711),
    .B(net297),
    .Y(_05239_));
 sky130_fd_sc_hd__o211a_1 _11125_ (.A1(net1432),
    .A2(net297),
    .B1(_05239_),
    .C1(net1183),
    .X(_00900_));
 sky130_fd_sc_hd__nand2_1 _11126_ (.A(_02585_),
    .B(net299),
    .Y(_05240_));
 sky130_fd_sc_hd__o211a_1 _11127_ (.A1(net1358),
    .A2(net299),
    .B1(_05240_),
    .C1(net1196),
    .X(_00901_));
 sky130_fd_sc_hd__or2_4 _11128_ (.A(net502),
    .B(_04976_),
    .X(_05241_));
 sky130_fd_sc_hd__a22o_1 _11129_ (.A1(_04515_),
    .A2(net453),
    .B1(net290),
    .B2(\reg_module.gprf[800] ),
    .X(_05242_));
 sky130_fd_sc_hd__and2_1 _11130_ (.A(net1124),
    .B(_05242_),
    .X(_00902_));
 sky130_fd_sc_hd__a22o_1 _11131_ (.A1(_04517_),
    .A2(net455),
    .B1(net290),
    .B2(\reg_module.gprf[801] ),
    .X(_05243_));
 sky130_fd_sc_hd__and2_1 _11132_ (.A(net1129),
    .B(_05243_),
    .X(_00903_));
 sky130_fd_sc_hd__a22o_1 _11133_ (.A1(_04519_),
    .A2(net448),
    .B1(net289),
    .B2(\reg_module.gprf[802] ),
    .X(_05244_));
 sky130_fd_sc_hd__and2_1 _11134_ (.A(net1107),
    .B(_05244_),
    .X(_00904_));
 sky130_fd_sc_hd__a22o_1 _11135_ (.A1(_04521_),
    .A2(net440),
    .B1(net289),
    .B2(\reg_module.gprf[803] ),
    .X(_05245_));
 sky130_fd_sc_hd__and2_1 _11136_ (.A(net1087),
    .B(_05245_),
    .X(_00905_));
 sky130_fd_sc_hd__a22o_1 _11137_ (.A1(_04523_),
    .A2(net455),
    .B1(net290),
    .B2(\reg_module.gprf[804] ),
    .X(_05246_));
 sky130_fd_sc_hd__and2_1 _11138_ (.A(net1127),
    .B(_05246_),
    .X(_00906_));
 sky130_fd_sc_hd__a22o_1 _11139_ (.A1(_04525_),
    .A2(net452),
    .B1(net290),
    .B2(\reg_module.gprf[805] ),
    .X(_05247_));
 sky130_fd_sc_hd__and2_1 _11140_ (.A(net1119),
    .B(_05247_),
    .X(_00907_));
 sky130_fd_sc_hd__a22o_1 _11141_ (.A1(_04527_),
    .A2(net439),
    .B1(net289),
    .B2(\reg_module.gprf[806] ),
    .X(_05248_));
 sky130_fd_sc_hd__and2_1 _11142_ (.A(net1081),
    .B(_05248_),
    .X(_00908_));
 sky130_fd_sc_hd__a22o_1 _11143_ (.A1(_04529_),
    .A2(net437),
    .B1(net289),
    .B2(\reg_module.gprf[807] ),
    .X(_05249_));
 sky130_fd_sc_hd__and2_1 _11144_ (.A(net1085),
    .B(_05249_),
    .X(_00909_));
 sky130_fd_sc_hd__a22o_1 _11145_ (.A1(_04531_),
    .A2(net456),
    .B1(net290),
    .B2(\reg_module.gprf[808] ),
    .X(_05250_));
 sky130_fd_sc_hd__and2_1 _11146_ (.A(net1122),
    .B(_05250_),
    .X(_00910_));
 sky130_fd_sc_hd__a22o_1 _11147_ (.A1(_04533_),
    .A2(net435),
    .B1(net289),
    .B2(\reg_module.gprf[809] ),
    .X(_05251_));
 sky130_fd_sc_hd__and2_1 _11148_ (.A(net1075),
    .B(_05251_),
    .X(_00911_));
 sky130_fd_sc_hd__a22o_1 _11149_ (.A1(_04535_),
    .A2(net435),
    .B1(net289),
    .B2(\reg_module.gprf[810] ),
    .X(_05252_));
 sky130_fd_sc_hd__and2_1 _11150_ (.A(net1074),
    .B(_05252_),
    .X(_00912_));
 sky130_fd_sc_hd__a22o_1 _11151_ (.A1(_04537_),
    .A2(net443),
    .B1(net289),
    .B2(\reg_module.gprf[811] ),
    .X(_05253_));
 sky130_fd_sc_hd__and2_1 _11152_ (.A(net1095),
    .B(_05253_),
    .X(_00913_));
 sky130_fd_sc_hd__a22o_1 _11153_ (.A1(_04539_),
    .A2(net460),
    .B1(net291),
    .B2(\reg_module.gprf[812] ),
    .X(_05254_));
 sky130_fd_sc_hd__and2_1 _11154_ (.A(net1143),
    .B(_05254_),
    .X(_00914_));
 sky130_fd_sc_hd__a22o_1 _11155_ (.A1(_04541_),
    .A2(net434),
    .B1(net289),
    .B2(\reg_module.gprf[813] ),
    .X(_05255_));
 sky130_fd_sc_hd__and2_1 _11156_ (.A(net1078),
    .B(_05255_),
    .X(_00915_));
 sky130_fd_sc_hd__a22o_1 _11157_ (.A1(_04543_),
    .A2(net450),
    .B1(net289),
    .B2(\reg_module.gprf[814] ),
    .X(_05256_));
 sky130_fd_sc_hd__and2_1 _11158_ (.A(net1116),
    .B(_05256_),
    .X(_00916_));
 sky130_fd_sc_hd__a22o_1 _11159_ (.A1(_04545_),
    .A2(net466),
    .B1(net291),
    .B2(\reg_module.gprf[815] ),
    .X(_05257_));
 sky130_fd_sc_hd__and2_1 _11160_ (.A(net1153),
    .B(_05257_),
    .X(_00917_));
 sky130_fd_sc_hd__a22o_1 _11161_ (.A1(_04547_),
    .A2(net484),
    .B1(net292),
    .B2(\reg_module.gprf[816] ),
    .X(_05258_));
 sky130_fd_sc_hd__and2_1 _11162_ (.A(net1202),
    .B(_05258_),
    .X(_00918_));
 sky130_fd_sc_hd__a22o_1 _11163_ (.A1(_04549_),
    .A2(net461),
    .B1(net291),
    .B2(\reg_module.gprf[817] ),
    .X(_05259_));
 sky130_fd_sc_hd__and2_1 _11164_ (.A(net1140),
    .B(_05259_),
    .X(_00919_));
 sky130_fd_sc_hd__a22o_1 _11165_ (.A1(_04551_),
    .A2(net461),
    .B1(net291),
    .B2(\reg_module.gprf[818] ),
    .X(_05260_));
 sky130_fd_sc_hd__and2_1 _11166_ (.A(net1139),
    .B(_05260_),
    .X(_00920_));
 sky130_fd_sc_hd__a22o_1 _11167_ (.A1(_04553_),
    .A2(net467),
    .B1(net291),
    .B2(\reg_module.gprf[819] ),
    .X(_05261_));
 sky130_fd_sc_hd__and2_1 _11168_ (.A(net1158),
    .B(_05261_),
    .X(_00921_));
 sky130_fd_sc_hd__a22o_1 _11169_ (.A1(_04555_),
    .A2(net449),
    .B1(net289),
    .B2(\reg_module.gprf[820] ),
    .X(_05262_));
 sky130_fd_sc_hd__and2_1 _11170_ (.A(net1117),
    .B(_05262_),
    .X(_00922_));
 sky130_fd_sc_hd__a22o_1 _11171_ (.A1(_04557_),
    .A2(net485),
    .B1(net292),
    .B2(\reg_module.gprf[821] ),
    .X(_05263_));
 sky130_fd_sc_hd__and2_1 _11172_ (.A(net1207),
    .B(_05263_),
    .X(_00923_));
 sky130_fd_sc_hd__a22o_1 _11173_ (.A1(_04559_),
    .A2(net481),
    .B1(net292),
    .B2(\reg_module.gprf[822] ),
    .X(_05264_));
 sky130_fd_sc_hd__and2_1 _11174_ (.A(net1196),
    .B(_05264_),
    .X(_00924_));
 sky130_fd_sc_hd__a22o_1 _11175_ (.A1(_04561_),
    .A2(net472),
    .B1(net291),
    .B2(\reg_module.gprf[823] ),
    .X(_05265_));
 sky130_fd_sc_hd__and2_1 _11176_ (.A(net1165),
    .B(_05265_),
    .X(_00925_));
 sky130_fd_sc_hd__a22o_1 _11177_ (.A1(_04563_),
    .A2(net478),
    .B1(net291),
    .B2(\reg_module.gprf[824] ),
    .X(_05266_));
 sky130_fd_sc_hd__and2_1 _11178_ (.A(net1183),
    .B(_05266_),
    .X(_00926_));
 sky130_fd_sc_hd__a22o_1 _11179_ (.A1(_04565_),
    .A2(net473),
    .B1(net292),
    .B2(\reg_module.gprf[825] ),
    .X(_05267_));
 sky130_fd_sc_hd__and2_1 _11180_ (.A(net1173),
    .B(_05267_),
    .X(_00927_));
 sky130_fd_sc_hd__a22o_1 _11181_ (.A1(_04567_),
    .A2(net467),
    .B1(net291),
    .B2(\reg_module.gprf[826] ),
    .X(_05268_));
 sky130_fd_sc_hd__and2_1 _11182_ (.A(net1163),
    .B(_05268_),
    .X(_00928_));
 sky130_fd_sc_hd__a22o_1 _11183_ (.A1(_04569_),
    .A2(net462),
    .B1(net292),
    .B2(\reg_module.gprf[827] ),
    .X(_05269_));
 sky130_fd_sc_hd__and2_1 _11184_ (.A(net1146),
    .B(_05269_),
    .X(_00929_));
 sky130_fd_sc_hd__a22o_1 _11185_ (.A1(_04571_),
    .A2(net473),
    .B1(net291),
    .B2(\reg_module.gprf[828] ),
    .X(_05270_));
 sky130_fd_sc_hd__and2_1 _11186_ (.A(net1174),
    .B(_05270_),
    .X(_00930_));
 sky130_fd_sc_hd__a22o_1 _11187_ (.A1(_04573_),
    .A2(net479),
    .B1(net291),
    .B2(\reg_module.gprf[829] ),
    .X(_05271_));
 sky130_fd_sc_hd__and2_1 _11188_ (.A(net1178),
    .B(_05271_),
    .X(_00931_));
 sky130_fd_sc_hd__a22o_1 _11189_ (.A1(_04575_),
    .A2(net480),
    .B1(net292),
    .B2(\reg_module.gprf[830] ),
    .X(_05272_));
 sky130_fd_sc_hd__and2_1 _11190_ (.A(net1192),
    .B(_05272_),
    .X(_00932_));
 sky130_fd_sc_hd__a22o_1 _11191_ (.A1(_04577_),
    .A2(net485),
    .B1(net292),
    .B2(\reg_module.gprf[831] ),
    .X(_05273_));
 sky130_fd_sc_hd__and2_1 _11192_ (.A(net1196),
    .B(_05273_),
    .X(_00933_));
 sky130_fd_sc_hd__or2_4 _11193_ (.A(net640),
    .B(_04976_),
    .X(_05274_));
 sky130_fd_sc_hd__a22o_1 _11194_ (.A1(_04581_),
    .A2(net453),
    .B1(net286),
    .B2(\reg_module.gprf[832] ),
    .X(_05275_));
 sky130_fd_sc_hd__and2_1 _11195_ (.A(net1124),
    .B(_05275_),
    .X(_00934_));
 sky130_fd_sc_hd__a22o_1 _11196_ (.A1(_04583_),
    .A2(net455),
    .B1(net286),
    .B2(\reg_module.gprf[833] ),
    .X(_05276_));
 sky130_fd_sc_hd__and2_1 _11197_ (.A(net1129),
    .B(_05276_),
    .X(_00935_));
 sky130_fd_sc_hd__a22o_1 _11198_ (.A1(_04585_),
    .A2(net448),
    .B1(net285),
    .B2(\reg_module.gprf[834] ),
    .X(_05277_));
 sky130_fd_sc_hd__and2_1 _11199_ (.A(net1110),
    .B(_05277_),
    .X(_00936_));
 sky130_fd_sc_hd__a22o_1 _11200_ (.A1(_04587_),
    .A2(net440),
    .B1(net285),
    .B2(\reg_module.gprf[835] ),
    .X(_05278_));
 sky130_fd_sc_hd__and2_1 _11201_ (.A(net1088),
    .B(_05278_),
    .X(_00937_));
 sky130_fd_sc_hd__a22o_1 _11202_ (.A1(_04589_),
    .A2(net455),
    .B1(net286),
    .B2(\reg_module.gprf[836] ),
    .X(_05279_));
 sky130_fd_sc_hd__and2_1 _11203_ (.A(net1127),
    .B(_05279_),
    .X(_00938_));
 sky130_fd_sc_hd__a22o_1 _11204_ (.A1(_04591_),
    .A2(net452),
    .B1(net286),
    .B2(\reg_module.gprf[837] ),
    .X(_05280_));
 sky130_fd_sc_hd__and2_1 _11205_ (.A(net1119),
    .B(_05280_),
    .X(_00939_));
 sky130_fd_sc_hd__a22o_1 _11206_ (.A1(_04593_),
    .A2(net439),
    .B1(net285),
    .B2(\reg_module.gprf[838] ),
    .X(_05281_));
 sky130_fd_sc_hd__and2_1 _11207_ (.A(net1081),
    .B(_05281_),
    .X(_00940_));
 sky130_fd_sc_hd__a22o_1 _11208_ (.A1(_04595_),
    .A2(net437),
    .B1(net285),
    .B2(\reg_module.gprf[839] ),
    .X(_05282_));
 sky130_fd_sc_hd__and2_1 _11209_ (.A(net1085),
    .B(_05282_),
    .X(_00941_));
 sky130_fd_sc_hd__a22o_1 _11210_ (.A1(_04597_),
    .A2(net456),
    .B1(net286),
    .B2(\reg_module.gprf[840] ),
    .X(_05283_));
 sky130_fd_sc_hd__and2_1 _11211_ (.A(net1122),
    .B(_05283_),
    .X(_00942_));
 sky130_fd_sc_hd__a22o_1 _11212_ (.A1(_04599_),
    .A2(net443),
    .B1(net285),
    .B2(\reg_module.gprf[841] ),
    .X(_05284_));
 sky130_fd_sc_hd__and2_1 _11213_ (.A(net1094),
    .B(_05284_),
    .X(_00943_));
 sky130_fd_sc_hd__a22o_1 _11214_ (.A1(_04601_),
    .A2(net435),
    .B1(net285),
    .B2(\reg_module.gprf[842] ),
    .X(_05285_));
 sky130_fd_sc_hd__and2_1 _11215_ (.A(net1074),
    .B(_05285_),
    .X(_00944_));
 sky130_fd_sc_hd__a22o_1 _11216_ (.A1(_04603_),
    .A2(net445),
    .B1(net285),
    .B2(\reg_module.gprf[843] ),
    .X(_05286_));
 sky130_fd_sc_hd__and2_1 _11217_ (.A(net1099),
    .B(_05286_),
    .X(_00945_));
 sky130_fd_sc_hd__a22o_1 _11218_ (.A1(_04605_),
    .A2(net460),
    .B1(net287),
    .B2(\reg_module.gprf[844] ),
    .X(_05287_));
 sky130_fd_sc_hd__and2_1 _11219_ (.A(net1143),
    .B(_05287_),
    .X(_00946_));
 sky130_fd_sc_hd__a22o_1 _11220_ (.A1(_04607_),
    .A2(net448),
    .B1(net285),
    .B2(\reg_module.gprf[845] ),
    .X(_05288_));
 sky130_fd_sc_hd__and2_1 _11221_ (.A(net1106),
    .B(_05288_),
    .X(_00947_));
 sky130_fd_sc_hd__a22o_1 _11222_ (.A1(_04609_),
    .A2(net450),
    .B1(net285),
    .B2(\reg_module.gprf[846] ),
    .X(_05289_));
 sky130_fd_sc_hd__and2_1 _11223_ (.A(net1116),
    .B(_05289_),
    .X(_00948_));
 sky130_fd_sc_hd__a22o_1 _11224_ (.A1(_04611_),
    .A2(net466),
    .B1(net287),
    .B2(\reg_module.gprf[847] ),
    .X(_05290_));
 sky130_fd_sc_hd__and2_1 _11225_ (.A(net1153),
    .B(_05290_),
    .X(_00949_));
 sky130_fd_sc_hd__a22o_1 _11226_ (.A1(_04613_),
    .A2(net483),
    .B1(net288),
    .B2(\reg_module.gprf[848] ),
    .X(_05291_));
 sky130_fd_sc_hd__and2_1 _11227_ (.A(net1201),
    .B(_05291_),
    .X(_00950_));
 sky130_fd_sc_hd__a22o_1 _11228_ (.A1(_04615_),
    .A2(net462),
    .B1(net287),
    .B2(\reg_module.gprf[849] ),
    .X(_05292_));
 sky130_fd_sc_hd__and2_1 _11229_ (.A(net1145),
    .B(_05292_),
    .X(_00951_));
 sky130_fd_sc_hd__a22o_1 _11230_ (.A1(_04617_),
    .A2(net461),
    .B1(net287),
    .B2(\reg_module.gprf[850] ),
    .X(_05293_));
 sky130_fd_sc_hd__and2_1 _11231_ (.A(net1139),
    .B(_05293_),
    .X(_00952_));
 sky130_fd_sc_hd__a22o_1 _11232_ (.A1(_04619_),
    .A2(net467),
    .B1(net287),
    .B2(\reg_module.gprf[851] ),
    .X(_05294_));
 sky130_fd_sc_hd__and2_1 _11233_ (.A(net1160),
    .B(_05294_),
    .X(_00953_));
 sky130_fd_sc_hd__a22o_1 _11234_ (.A1(_04621_),
    .A2(net449),
    .B1(net285),
    .B2(\reg_module.gprf[852] ),
    .X(_05295_));
 sky130_fd_sc_hd__and2_1 _11235_ (.A(net1114),
    .B(_05295_),
    .X(_00954_));
 sky130_fd_sc_hd__a22o_1 _11236_ (.A1(_04623_),
    .A2(net485),
    .B1(net288),
    .B2(\reg_module.gprf[853] ),
    .X(_05296_));
 sky130_fd_sc_hd__and2_1 _11237_ (.A(net1208),
    .B(_05296_),
    .X(_00955_));
 sky130_fd_sc_hd__a22o_1 _11238_ (.A1(_04625_),
    .A2(net480),
    .B1(net288),
    .B2(\reg_module.gprf[854] ),
    .X(_05297_));
 sky130_fd_sc_hd__and2_1 _11239_ (.A(net1196),
    .B(_05297_),
    .X(_00956_));
 sky130_fd_sc_hd__a22o_1 _11240_ (.A1(_04627_),
    .A2(net472),
    .B1(net287),
    .B2(\reg_module.gprf[855] ),
    .X(_05298_));
 sky130_fd_sc_hd__and2_1 _11241_ (.A(net1165),
    .B(_05298_),
    .X(_00957_));
 sky130_fd_sc_hd__a22o_1 _11242_ (.A1(_04629_),
    .A2(net478),
    .B1(net287),
    .B2(\reg_module.gprf[856] ),
    .X(_05299_));
 sky130_fd_sc_hd__and2_1 _11243_ (.A(net1183),
    .B(_05299_),
    .X(_00958_));
 sky130_fd_sc_hd__a22o_1 _11244_ (.A1(_04631_),
    .A2(net474),
    .B1(net287),
    .B2(\reg_module.gprf[857] ),
    .X(_05300_));
 sky130_fd_sc_hd__and2_1 _11245_ (.A(net1173),
    .B(_05300_),
    .X(_00959_));
 sky130_fd_sc_hd__a22o_1 _11246_ (.A1(_04633_),
    .A2(net467),
    .B1(net287),
    .B2(\reg_module.gprf[858] ),
    .X(_05301_));
 sky130_fd_sc_hd__and2_1 _11247_ (.A(net1160),
    .B(_05301_),
    .X(_00960_));
 sky130_fd_sc_hd__a22o_1 _11248_ (.A1(_04635_),
    .A2(net464),
    .B1(net287),
    .B2(\reg_module.gprf[859] ),
    .X(_05302_));
 sky130_fd_sc_hd__and2_1 _11249_ (.A(net1146),
    .B(_05302_),
    .X(_00961_));
 sky130_fd_sc_hd__a22o_1 _11250_ (.A1(_04637_),
    .A2(net473),
    .B1(net288),
    .B2(\reg_module.gprf[860] ),
    .X(_05303_));
 sky130_fd_sc_hd__and2_1 _11251_ (.A(net1174),
    .B(_05303_),
    .X(_00962_));
 sky130_fd_sc_hd__a22o_1 _11252_ (.A1(_04639_),
    .A2(net476),
    .B1(net288),
    .B2(\reg_module.gprf[861] ),
    .X(_05304_));
 sky130_fd_sc_hd__and2_1 _11253_ (.A(net1179),
    .B(_05304_),
    .X(_00963_));
 sky130_fd_sc_hd__a22o_1 _11254_ (.A1(_04641_),
    .A2(net480),
    .B1(net288),
    .B2(\reg_module.gprf[862] ),
    .X(_05305_));
 sky130_fd_sc_hd__and2_1 _11255_ (.A(net1193),
    .B(_05305_),
    .X(_00964_));
 sky130_fd_sc_hd__a22o_1 _11256_ (.A1(_04643_),
    .A2(net485),
    .B1(net288),
    .B2(\reg_module.gprf[863] ),
    .X(_05306_));
 sky130_fd_sc_hd__and2_1 _11257_ (.A(net1196),
    .B(_05306_),
    .X(_00965_));
 sky130_fd_sc_hd__or2_4 _11258_ (.A(net636),
    .B(_04976_),
    .X(_05307_));
 sky130_fd_sc_hd__a22o_1 _11259_ (.A1(_04647_),
    .A2(net453),
    .B1(net282),
    .B2(\reg_module.gprf[864] ),
    .X(_05308_));
 sky130_fd_sc_hd__and2_1 _11260_ (.A(net1125),
    .B(_05308_),
    .X(_00966_));
 sky130_fd_sc_hd__a22o_1 _11261_ (.A1(_04649_),
    .A2(net455),
    .B1(net282),
    .B2(\reg_module.gprf[865] ),
    .X(_05309_));
 sky130_fd_sc_hd__and2_1 _11262_ (.A(net1131),
    .B(_05309_),
    .X(_00967_));
 sky130_fd_sc_hd__a22o_1 _11263_ (.A1(_04651_),
    .A2(net448),
    .B1(net281),
    .B2(\reg_module.gprf[866] ),
    .X(_05310_));
 sky130_fd_sc_hd__and2_1 _11264_ (.A(net1107),
    .B(_05310_),
    .X(_00968_));
 sky130_fd_sc_hd__a22o_1 _11265_ (.A1(_04653_),
    .A2(net440),
    .B1(net281),
    .B2(\reg_module.gprf[867] ),
    .X(_05311_));
 sky130_fd_sc_hd__and2_1 _11266_ (.A(net1092),
    .B(_05311_),
    .X(_00969_));
 sky130_fd_sc_hd__a22o_1 _11267_ (.A1(_04655_),
    .A2(net455),
    .B1(net282),
    .B2(\reg_module.gprf[868] ),
    .X(_05312_));
 sky130_fd_sc_hd__and2_1 _11268_ (.A(net1127),
    .B(_05312_),
    .X(_00970_));
 sky130_fd_sc_hd__a22o_1 _11269_ (.A1(_04657_),
    .A2(net452),
    .B1(net282),
    .B2(\reg_module.gprf[869] ),
    .X(_05313_));
 sky130_fd_sc_hd__and2_1 _11270_ (.A(net1119),
    .B(_05313_),
    .X(_00971_));
 sky130_fd_sc_hd__a22o_1 _11271_ (.A1(_04659_),
    .A2(net439),
    .B1(net281),
    .B2(\reg_module.gprf[870] ),
    .X(_05314_));
 sky130_fd_sc_hd__and2_1 _11272_ (.A(net1081),
    .B(_05314_),
    .X(_00972_));
 sky130_fd_sc_hd__a22o_1 _11273_ (.A1(_04661_),
    .A2(net437),
    .B1(net281),
    .B2(\reg_module.gprf[871] ),
    .X(_05315_));
 sky130_fd_sc_hd__and2_1 _11274_ (.A(net1085),
    .B(_05315_),
    .X(_00973_));
 sky130_fd_sc_hd__a22o_1 _11275_ (.A1(_04663_),
    .A2(net456),
    .B1(net282),
    .B2(\reg_module.gprf[872] ),
    .X(_05316_));
 sky130_fd_sc_hd__and2_1 _11276_ (.A(net1122),
    .B(_05316_),
    .X(_00974_));
 sky130_fd_sc_hd__a22o_1 _11277_ (.A1(_04665_),
    .A2(net443),
    .B1(net281),
    .B2(\reg_module.gprf[873] ),
    .X(_05317_));
 sky130_fd_sc_hd__and2_1 _11278_ (.A(net1094),
    .B(_05317_),
    .X(_00975_));
 sky130_fd_sc_hd__a22o_1 _11279_ (.A1(_04667_),
    .A2(net435),
    .B1(net281),
    .B2(\reg_module.gprf[874] ),
    .X(_05318_));
 sky130_fd_sc_hd__and2_1 _11280_ (.A(net1075),
    .B(_05318_),
    .X(_00976_));
 sky130_fd_sc_hd__a22o_1 _11281_ (.A1(_04669_),
    .A2(net445),
    .B1(net281),
    .B2(\reg_module.gprf[875] ),
    .X(_05319_));
 sky130_fd_sc_hd__and2_1 _11282_ (.A(net1099),
    .B(_05319_),
    .X(_00977_));
 sky130_fd_sc_hd__a22o_1 _11283_ (.A1(_04671_),
    .A2(net461),
    .B1(net283),
    .B2(\reg_module.gprf[876] ),
    .X(_05320_));
 sky130_fd_sc_hd__and2_1 _11284_ (.A(net1144),
    .B(_05320_),
    .X(_00978_));
 sky130_fd_sc_hd__a22o_1 _11285_ (.A1(_04673_),
    .A2(net443),
    .B1(net281),
    .B2(\reg_module.gprf[877] ),
    .X(_05321_));
 sky130_fd_sc_hd__and2_1 _11286_ (.A(net1097),
    .B(_05321_),
    .X(_00979_));
 sky130_fd_sc_hd__a22o_1 _11287_ (.A1(_04675_),
    .A2(net465),
    .B1(net281),
    .B2(\reg_module.gprf[878] ),
    .X(_05322_));
 sky130_fd_sc_hd__and2_1 _11288_ (.A(net1116),
    .B(_05322_),
    .X(_00980_));
 sky130_fd_sc_hd__a22o_1 _11289_ (.A1(_04677_),
    .A2(net467),
    .B1(net283),
    .B2(\reg_module.gprf[879] ),
    .X(_05323_));
 sky130_fd_sc_hd__and2_1 _11290_ (.A(net1160),
    .B(_05323_),
    .X(_00981_));
 sky130_fd_sc_hd__a22o_1 _11291_ (.A1(_04679_),
    .A2(net483),
    .B1(net284),
    .B2(\reg_module.gprf[880] ),
    .X(_05324_));
 sky130_fd_sc_hd__and2_1 _11292_ (.A(net1201),
    .B(_05324_),
    .X(_00982_));
 sky130_fd_sc_hd__a22o_1 _11293_ (.A1(_04681_),
    .A2(net462),
    .B1(net283),
    .B2(\reg_module.gprf[881] ),
    .X(_05325_));
 sky130_fd_sc_hd__and2_1 _11294_ (.A(net1145),
    .B(_05325_),
    .X(_00983_));
 sky130_fd_sc_hd__a22o_1 _11295_ (.A1(_04683_),
    .A2(net461),
    .B1(net283),
    .B2(\reg_module.gprf[882] ),
    .X(_05326_));
 sky130_fd_sc_hd__and2_1 _11296_ (.A(net1139),
    .B(_05326_),
    .X(_00984_));
 sky130_fd_sc_hd__a22o_1 _11297_ (.A1(_04685_),
    .A2(net467),
    .B1(net283),
    .B2(\reg_module.gprf[883] ),
    .X(_05327_));
 sky130_fd_sc_hd__and2_1 _11298_ (.A(net1159),
    .B(_05327_),
    .X(_00985_));
 sky130_fd_sc_hd__a22o_1 _11299_ (.A1(_04687_),
    .A2(net449),
    .B1(net281),
    .B2(\reg_module.gprf[884] ),
    .X(_05328_));
 sky130_fd_sc_hd__and2_1 _11300_ (.A(net1114),
    .B(_05328_),
    .X(_00986_));
 sky130_fd_sc_hd__a22o_1 _11301_ (.A1(_04689_),
    .A2(net486),
    .B1(net284),
    .B2(\reg_module.gprf[885] ),
    .X(_05329_));
 sky130_fd_sc_hd__and2_1 _11302_ (.A(net1208),
    .B(_05329_),
    .X(_00987_));
 sky130_fd_sc_hd__a22o_1 _11303_ (.A1(_04691_),
    .A2(net480),
    .B1(net284),
    .B2(\reg_module.gprf[886] ),
    .X(_05330_));
 sky130_fd_sc_hd__and2_1 _11304_ (.A(net1196),
    .B(_05330_),
    .X(_00988_));
 sky130_fd_sc_hd__a22o_1 _11305_ (.A1(_04693_),
    .A2(net472),
    .B1(net283),
    .B2(\reg_module.gprf[887] ),
    .X(_05331_));
 sky130_fd_sc_hd__and2_1 _11306_ (.A(net1165),
    .B(_05331_),
    .X(_00989_));
 sky130_fd_sc_hd__a22o_1 _11307_ (.A1(_04695_),
    .A2(net478),
    .B1(net283),
    .B2(\reg_module.gprf[888] ),
    .X(_05332_));
 sky130_fd_sc_hd__and2_1 _11308_ (.A(net1185),
    .B(_05332_),
    .X(_00990_));
 sky130_fd_sc_hd__a22o_1 _11309_ (.A1(_04697_),
    .A2(net474),
    .B1(net283),
    .B2(\reg_module.gprf[889] ),
    .X(_05333_));
 sky130_fd_sc_hd__and2_1 _11310_ (.A(net1173),
    .B(_05333_),
    .X(_00991_));
 sky130_fd_sc_hd__a22o_1 _11311_ (.A1(_04699_),
    .A2(net479),
    .B1(net283),
    .B2(\reg_module.gprf[890] ),
    .X(_05334_));
 sky130_fd_sc_hd__and2_1 _11312_ (.A(net1178),
    .B(_05334_),
    .X(_00992_));
 sky130_fd_sc_hd__a22o_1 _11313_ (.A1(_04701_),
    .A2(net472),
    .B1(net283),
    .B2(\reg_module.gprf[891] ),
    .X(_05335_));
 sky130_fd_sc_hd__and2_1 _11314_ (.A(net1164),
    .B(_05335_),
    .X(_00993_));
 sky130_fd_sc_hd__a22o_1 _11315_ (.A1(_04703_),
    .A2(net473),
    .B1(net284),
    .B2(\reg_module.gprf[892] ),
    .X(_05336_));
 sky130_fd_sc_hd__and2_1 _11316_ (.A(net1174),
    .B(_05336_),
    .X(_00994_));
 sky130_fd_sc_hd__a22o_1 _11317_ (.A1(_04705_),
    .A2(net476),
    .B1(net284),
    .B2(\reg_module.gprf[893] ),
    .X(_05337_));
 sky130_fd_sc_hd__and2_1 _11318_ (.A(net1179),
    .B(_05337_),
    .X(_00995_));
 sky130_fd_sc_hd__a22o_1 _11319_ (.A1(_04707_),
    .A2(net478),
    .B1(net284),
    .B2(\reg_module.gprf[894] ),
    .X(_05338_));
 sky130_fd_sc_hd__and2_1 _11320_ (.A(net1184),
    .B(_05338_),
    .X(_00996_));
 sky130_fd_sc_hd__a22o_1 _11321_ (.A1(_04709_),
    .A2(net485),
    .B1(net284),
    .B2(\reg_module.gprf[895] ),
    .X(_05339_));
 sky130_fd_sc_hd__and2_1 _11322_ (.A(net1197),
    .B(_05339_),
    .X(_00997_));
 sky130_fd_sc_hd__or2_2 _11323_ (.A(net498),
    .B(_04976_),
    .X(_05340_));
 sky130_fd_sc_hd__a22o_1 _11324_ (.A1(_04713_),
    .A2(net453),
    .B1(net278),
    .B2(\reg_module.gprf[896] ),
    .X(_05341_));
 sky130_fd_sc_hd__and2_1 _11325_ (.A(net1124),
    .B(_05341_),
    .X(_00998_));
 sky130_fd_sc_hd__a22o_1 _11326_ (.A1(_04715_),
    .A2(net458),
    .B1(net278),
    .B2(\reg_module.gprf[897] ),
    .X(_05342_));
 sky130_fd_sc_hd__and2_1 _11327_ (.A(net1132),
    .B(_05342_),
    .X(_00999_));
 sky130_fd_sc_hd__a22o_1 _11328_ (.A1(_04717_),
    .A2(net447),
    .B1(net277),
    .B2(\reg_module.gprf[898] ),
    .X(_05343_));
 sky130_fd_sc_hd__and2_1 _11329_ (.A(net1111),
    .B(_05343_),
    .X(_01000_));
 sky130_fd_sc_hd__a22o_1 _11330_ (.A1(_04719_),
    .A2(net441),
    .B1(net277),
    .B2(\reg_module.gprf[899] ),
    .X(_05344_));
 sky130_fd_sc_hd__and2_1 _11331_ (.A(net1090),
    .B(_05344_),
    .X(_01001_));
 sky130_fd_sc_hd__a22o_1 _11332_ (.A1(_04721_),
    .A2(net458),
    .B1(net278),
    .B2(\reg_module.gprf[900] ),
    .X(_05345_));
 sky130_fd_sc_hd__and2_1 _11333_ (.A(net1130),
    .B(_05345_),
    .X(_01002_));
 sky130_fd_sc_hd__a22o_1 _11334_ (.A1(_04723_),
    .A2(net452),
    .B1(net278),
    .B2(\reg_module.gprf[901] ),
    .X(_05346_));
 sky130_fd_sc_hd__and2_1 _11335_ (.A(net1119),
    .B(_05346_),
    .X(_01003_));
 sky130_fd_sc_hd__a22o_1 _11336_ (.A1(_04725_),
    .A2(net439),
    .B1(net277),
    .B2(\reg_module.gprf[902] ),
    .X(_05347_));
 sky130_fd_sc_hd__and2_1 _11337_ (.A(net1081),
    .B(_05347_),
    .X(_01004_));
 sky130_fd_sc_hd__a22o_1 _11338_ (.A1(_04727_),
    .A2(net438),
    .B1(net277),
    .B2(\reg_module.gprf[903] ),
    .X(_05348_));
 sky130_fd_sc_hd__and2_1 _11339_ (.A(net1084),
    .B(_05348_),
    .X(_01005_));
 sky130_fd_sc_hd__a22o_1 _11340_ (.A1(_04729_),
    .A2(net452),
    .B1(net278),
    .B2(\reg_module.gprf[904] ),
    .X(_05349_));
 sky130_fd_sc_hd__and2_1 _11341_ (.A(net1123),
    .B(_05349_),
    .X(_01006_));
 sky130_fd_sc_hd__a22o_1 _11342_ (.A1(_04731_),
    .A2(net435),
    .B1(net277),
    .B2(\reg_module.gprf[905] ),
    .X(_05350_));
 sky130_fd_sc_hd__and2_1 _11343_ (.A(net1076),
    .B(_05350_),
    .X(_01007_));
 sky130_fd_sc_hd__a22o_1 _11344_ (.A1(_04733_),
    .A2(net433),
    .B1(net277),
    .B2(\reg_module.gprf[906] ),
    .X(_05351_));
 sky130_fd_sc_hd__and2_1 _11345_ (.A(net1073),
    .B(_05351_),
    .X(_01008_));
 sky130_fd_sc_hd__a22o_1 _11346_ (.A1(_04735_),
    .A2(net443),
    .B1(net277),
    .B2(\reg_module.gprf[907] ),
    .X(_05352_));
 sky130_fd_sc_hd__and2_1 _11347_ (.A(net1096),
    .B(_05352_),
    .X(_01009_));
 sky130_fd_sc_hd__a22o_1 _11348_ (.A1(_04737_),
    .A2(net466),
    .B1(net279),
    .B2(\reg_module.gprf[908] ),
    .X(_05353_));
 sky130_fd_sc_hd__and2_1 _11349_ (.A(net1152),
    .B(_05353_),
    .X(_01010_));
 sky130_fd_sc_hd__a22o_1 _11350_ (.A1(_04739_),
    .A2(net434),
    .B1(net277),
    .B2(\reg_module.gprf[909] ),
    .X(_05354_));
 sky130_fd_sc_hd__and2_1 _11351_ (.A(net1078),
    .B(_05354_),
    .X(_01011_));
 sky130_fd_sc_hd__a22o_1 _11352_ (.A1(_04741_),
    .A2(net459),
    .B1(net278),
    .B2(\reg_module.gprf[910] ),
    .X(_05355_));
 sky130_fd_sc_hd__and2_1 _11353_ (.A(net1136),
    .B(_05355_),
    .X(_01012_));
 sky130_fd_sc_hd__a22o_1 _11354_ (.A1(_04743_),
    .A2(net465),
    .B1(net279),
    .B2(\reg_module.gprf[911] ),
    .X(_05356_));
 sky130_fd_sc_hd__and2_1 _11355_ (.A(net1157),
    .B(_05356_),
    .X(_01013_));
 sky130_fd_sc_hd__a22o_1 _11356_ (.A1(_04745_),
    .A2(net487),
    .B1(net280),
    .B2(\reg_module.gprf[912] ),
    .X(_05357_));
 sky130_fd_sc_hd__and2_1 _11357_ (.A(net1189),
    .B(_05357_),
    .X(_01014_));
 sky130_fd_sc_hd__a22o_1 _11358_ (.A1(_04747_),
    .A2(net462),
    .B1(net279),
    .B2(\reg_module.gprf[913] ),
    .X(_05358_));
 sky130_fd_sc_hd__and2_1 _11359_ (.A(net1140),
    .B(_05358_),
    .X(_01015_));
 sky130_fd_sc_hd__a22o_1 _11360_ (.A1(_04749_),
    .A2(net445),
    .B1(net277),
    .B2(\reg_module.gprf[914] ),
    .X(_05359_));
 sky130_fd_sc_hd__and2_1 _11361_ (.A(net1101),
    .B(_05359_),
    .X(_01016_));
 sky130_fd_sc_hd__a22o_1 _11362_ (.A1(_04751_),
    .A2(net467),
    .B1(net279),
    .B2(\reg_module.gprf[915] ),
    .X(_05360_));
 sky130_fd_sc_hd__and2_1 _11363_ (.A(net1158),
    .B(_05360_),
    .X(_01017_));
 sky130_fd_sc_hd__a22o_1 _11364_ (.A1(_04753_),
    .A2(net449),
    .B1(net277),
    .B2(\reg_module.gprf[916] ),
    .X(_05361_));
 sky130_fd_sc_hd__and2_1 _11365_ (.A(net1114),
    .B(_05361_),
    .X(_01018_));
 sky130_fd_sc_hd__a22o_1 _11366_ (.A1(_04755_),
    .A2(net484),
    .B1(net280),
    .B2(\reg_module.gprf[917] ),
    .X(_05362_));
 sky130_fd_sc_hd__and2_1 _11367_ (.A(net1203),
    .B(_05362_),
    .X(_01019_));
 sky130_fd_sc_hd__a22o_1 _11368_ (.A1(_04757_),
    .A2(net481),
    .B1(net280),
    .B2(\reg_module.gprf[918] ),
    .X(_05363_));
 sky130_fd_sc_hd__and2_1 _11369_ (.A(net1197),
    .B(_05363_),
    .X(_01020_));
 sky130_fd_sc_hd__a22o_1 _11370_ (.A1(_04759_),
    .A2(net472),
    .B1(net279),
    .B2(\reg_module.gprf[919] ),
    .X(_05364_));
 sky130_fd_sc_hd__and2_1 _11371_ (.A(net1164),
    .B(_05364_),
    .X(_01021_));
 sky130_fd_sc_hd__a22o_1 _11372_ (.A1(_04761_),
    .A2(net477),
    .B1(net279),
    .B2(\reg_module.gprf[920] ),
    .X(_05365_));
 sky130_fd_sc_hd__and2_1 _11373_ (.A(net1183),
    .B(_05365_),
    .X(_01022_));
 sky130_fd_sc_hd__a22o_1 _11374_ (.A1(_04763_),
    .A2(net477),
    .B1(net279),
    .B2(\reg_module.gprf[921] ),
    .X(_05366_));
 sky130_fd_sc_hd__and2_1 _11375_ (.A(net1180),
    .B(_05366_),
    .X(_01023_));
 sky130_fd_sc_hd__a22o_1 _11376_ (.A1(_04765_),
    .A2(net467),
    .B1(net280),
    .B2(\reg_module.gprf[922] ),
    .X(_05367_));
 sky130_fd_sc_hd__and2_1 _11377_ (.A(net1163),
    .B(_05367_),
    .X(_01024_));
 sky130_fd_sc_hd__a22o_1 _11378_ (.A1(_04767_),
    .A2(net462),
    .B1(net279),
    .B2(\reg_module.gprf[923] ),
    .X(_05368_));
 sky130_fd_sc_hd__and2_1 _11379_ (.A(net1145),
    .B(_05368_),
    .X(_01025_));
 sky130_fd_sc_hd__a22o_1 _11380_ (.A1(_04769_),
    .A2(net473),
    .B1(net279),
    .B2(\reg_module.gprf[924] ),
    .X(_05369_));
 sky130_fd_sc_hd__and2_1 _11381_ (.A(net1172),
    .B(_05369_),
    .X(_01026_));
 sky130_fd_sc_hd__a22o_1 _11382_ (.A1(_04771_),
    .A2(net475),
    .B1(net279),
    .B2(\reg_module.gprf[925] ),
    .X(_05370_));
 sky130_fd_sc_hd__and2_1 _11383_ (.A(net1175),
    .B(_05370_),
    .X(_01027_));
 sky130_fd_sc_hd__a22o_1 _11384_ (.A1(_04773_),
    .A2(net480),
    .B1(net280),
    .B2(\reg_module.gprf[926] ),
    .X(_05371_));
 sky130_fd_sc_hd__and2_1 _11385_ (.A(net1193),
    .B(_05371_),
    .X(_01028_));
 sky130_fd_sc_hd__a22o_1 _11386_ (.A1(_04775_),
    .A2(net485),
    .B1(net280),
    .B2(\reg_module.gprf[927] ),
    .X(_05372_));
 sky130_fd_sc_hd__and2_1 _11387_ (.A(net1205),
    .B(_05372_),
    .X(_01029_));
 sky130_fd_sc_hd__or2_2 _11388_ (.A(net494),
    .B(_04976_),
    .X(_05373_));
 sky130_fd_sc_hd__a22o_1 _11389_ (.A1(_04779_),
    .A2(net453),
    .B1(net274),
    .B2(\reg_module.gprf[928] ),
    .X(_05374_));
 sky130_fd_sc_hd__and2_1 _11390_ (.A(net1124),
    .B(_05374_),
    .X(_01030_));
 sky130_fd_sc_hd__a22o_1 _11391_ (.A1(_04781_),
    .A2(net457),
    .B1(net274),
    .B2(\reg_module.gprf[929] ),
    .X(_05375_));
 sky130_fd_sc_hd__and2_1 _11392_ (.A(net1132),
    .B(_05375_),
    .X(_01031_));
 sky130_fd_sc_hd__a22o_1 _11393_ (.A1(_04783_),
    .A2(net447),
    .B1(net273),
    .B2(\reg_module.gprf[930] ),
    .X(_05376_));
 sky130_fd_sc_hd__and2_1 _11394_ (.A(net1111),
    .B(_05376_),
    .X(_01032_));
 sky130_fd_sc_hd__a22o_1 _11395_ (.A1(_04785_),
    .A2(net441),
    .B1(net273),
    .B2(\reg_module.gprf[931] ),
    .X(_05377_));
 sky130_fd_sc_hd__and2_1 _11396_ (.A(net1089),
    .B(_05377_),
    .X(_01033_));
 sky130_fd_sc_hd__a22o_1 _11397_ (.A1(_04787_),
    .A2(net455),
    .B1(net274),
    .B2(\reg_module.gprf[932] ),
    .X(_05378_));
 sky130_fd_sc_hd__and2_1 _11398_ (.A(net1130),
    .B(_05378_),
    .X(_01034_));
 sky130_fd_sc_hd__a22o_1 _11399_ (.A1(_04789_),
    .A2(net452),
    .B1(net274),
    .B2(\reg_module.gprf[933] ),
    .X(_05379_));
 sky130_fd_sc_hd__and2_1 _11400_ (.A(net1119),
    .B(_05379_),
    .X(_01035_));
 sky130_fd_sc_hd__a22o_1 _11401_ (.A1(_04791_),
    .A2(net439),
    .B1(net273),
    .B2(\reg_module.gprf[934] ),
    .X(_05380_));
 sky130_fd_sc_hd__and2_1 _11402_ (.A(net1081),
    .B(_05380_),
    .X(_01036_));
 sky130_fd_sc_hd__a22o_1 _11403_ (.A1(_04793_),
    .A2(net437),
    .B1(net273),
    .B2(\reg_module.gprf[935] ),
    .X(_05381_));
 sky130_fd_sc_hd__and2_1 _11404_ (.A(net1084),
    .B(_05381_),
    .X(_01037_));
 sky130_fd_sc_hd__a22o_1 _11405_ (.A1(_04795_),
    .A2(net454),
    .B1(net274),
    .B2(\reg_module.gprf[936] ),
    .X(_05382_));
 sky130_fd_sc_hd__and2_1 _11406_ (.A(net1123),
    .B(_05382_),
    .X(_01038_));
 sky130_fd_sc_hd__a22o_1 _11407_ (.A1(_04797_),
    .A2(net435),
    .B1(net273),
    .B2(\reg_module.gprf[937] ),
    .X(_05383_));
 sky130_fd_sc_hd__and2_1 _11408_ (.A(net1075),
    .B(_05383_),
    .X(_01039_));
 sky130_fd_sc_hd__a22o_1 _11409_ (.A1(_04799_),
    .A2(net433),
    .B1(net273),
    .B2(\reg_module.gprf[938] ),
    .X(_05384_));
 sky130_fd_sc_hd__and2_1 _11410_ (.A(net1073),
    .B(_05384_),
    .X(_01040_));
 sky130_fd_sc_hd__a22o_1 _11411_ (.A1(_04801_),
    .A2(net443),
    .B1(net273),
    .B2(\reg_module.gprf[939] ),
    .X(_05385_));
 sky130_fd_sc_hd__and2_1 _11412_ (.A(net1095),
    .B(_05385_),
    .X(_01041_));
 sky130_fd_sc_hd__a22o_1 _11413_ (.A1(_04803_),
    .A2(net466),
    .B1(net275),
    .B2(\reg_module.gprf[940] ),
    .X(_05386_));
 sky130_fd_sc_hd__and2_1 _11414_ (.A(net1152),
    .B(_05386_),
    .X(_01042_));
 sky130_fd_sc_hd__a22o_1 _11415_ (.A1(_04805_),
    .A2(net434),
    .B1(net273),
    .B2(\reg_module.gprf[941] ),
    .X(_05387_));
 sky130_fd_sc_hd__and2_1 _11416_ (.A(net1079),
    .B(_05387_),
    .X(_01043_));
 sky130_fd_sc_hd__a22o_1 _11417_ (.A1(_04807_),
    .A2(net450),
    .B1(net273),
    .B2(\reg_module.gprf[942] ),
    .X(_05388_));
 sky130_fd_sc_hd__and2_1 _11418_ (.A(net1116),
    .B(_05388_),
    .X(_01044_));
 sky130_fd_sc_hd__a22o_1 _11419_ (.A1(_04809_),
    .A2(net465),
    .B1(net275),
    .B2(\reg_module.gprf[943] ),
    .X(_05389_));
 sky130_fd_sc_hd__and2_1 _11420_ (.A(net1156),
    .B(_05389_),
    .X(_01045_));
 sky130_fd_sc_hd__a22o_1 _11421_ (.A1(_04811_),
    .A2(net487),
    .B1(net276),
    .B2(\reg_module.gprf[944] ),
    .X(_05390_));
 sky130_fd_sc_hd__and2_1 _11422_ (.A(net1189),
    .B(_05390_),
    .X(_01046_));
 sky130_fd_sc_hd__a22o_1 _11423_ (.A1(_04813_),
    .A2(net461),
    .B1(net275),
    .B2(\reg_module.gprf[945] ),
    .X(_05391_));
 sky130_fd_sc_hd__and2_1 _11424_ (.A(net1140),
    .B(_05391_),
    .X(_01047_));
 sky130_fd_sc_hd__a22o_1 _11425_ (.A1(_04815_),
    .A2(net445),
    .B1(net274),
    .B2(\reg_module.gprf[946] ),
    .X(_05392_));
 sky130_fd_sc_hd__and2_1 _11426_ (.A(net1101),
    .B(_05392_),
    .X(_01048_));
 sky130_fd_sc_hd__a22o_1 _11427_ (.A1(_04817_),
    .A2(net466),
    .B1(net275),
    .B2(\reg_module.gprf[947] ),
    .X(_05393_));
 sky130_fd_sc_hd__and2_1 _11428_ (.A(net1153),
    .B(_05393_),
    .X(_01049_));
 sky130_fd_sc_hd__a22o_1 _11429_ (.A1(_04819_),
    .A2(net449),
    .B1(net273),
    .B2(\reg_module.gprf[948] ),
    .X(_05394_));
 sky130_fd_sc_hd__and2_1 _11430_ (.A(net1117),
    .B(_05394_),
    .X(_01050_));
 sky130_fd_sc_hd__a22o_1 _11431_ (.A1(_04821_),
    .A2(net484),
    .B1(net276),
    .B2(\reg_module.gprf[949] ),
    .X(_05395_));
 sky130_fd_sc_hd__and2_1 _11432_ (.A(net1203),
    .B(_05395_),
    .X(_01051_));
 sky130_fd_sc_hd__a22o_1 _11433_ (.A1(_04823_),
    .A2(net481),
    .B1(net276),
    .B2(\reg_module.gprf[950] ),
    .X(_05396_));
 sky130_fd_sc_hd__and2_1 _11434_ (.A(net1197),
    .B(_05396_),
    .X(_01052_));
 sky130_fd_sc_hd__a22o_1 _11435_ (.A1(_04825_),
    .A2(net472),
    .B1(net275),
    .B2(\reg_module.gprf[951] ),
    .X(_05397_));
 sky130_fd_sc_hd__and2_1 _11436_ (.A(net1166),
    .B(_05397_),
    .X(_01053_));
 sky130_fd_sc_hd__a22o_1 _11437_ (.A1(_04827_),
    .A2(net478),
    .B1(net275),
    .B2(\reg_module.gprf[952] ),
    .X(_05398_));
 sky130_fd_sc_hd__and2_1 _11438_ (.A(net1183),
    .B(_05398_),
    .X(_01054_));
 sky130_fd_sc_hd__a22o_1 _11439_ (.A1(_04829_),
    .A2(net477),
    .B1(net275),
    .B2(\reg_module.gprf[953] ),
    .X(_05399_));
 sky130_fd_sc_hd__and2_1 _11440_ (.A(net1180),
    .B(_05399_),
    .X(_01055_));
 sky130_fd_sc_hd__a22o_1 _11441_ (.A1(_04831_),
    .A2(net468),
    .B1(net276),
    .B2(\reg_module.gprf[954] ),
    .X(_05400_));
 sky130_fd_sc_hd__and2_1 _11442_ (.A(net1163),
    .B(_05400_),
    .X(_01056_));
 sky130_fd_sc_hd__a22o_1 _11443_ (.A1(_04833_),
    .A2(net462),
    .B1(net275),
    .B2(\reg_module.gprf[955] ),
    .X(_05401_));
 sky130_fd_sc_hd__and2_1 _11444_ (.A(net1145),
    .B(_05401_),
    .X(_01057_));
 sky130_fd_sc_hd__a22o_1 _11445_ (.A1(_04835_),
    .A2(net473),
    .B1(net275),
    .B2(\reg_module.gprf[956] ),
    .X(_05402_));
 sky130_fd_sc_hd__and2_1 _11446_ (.A(net1171),
    .B(_05402_),
    .X(_01058_));
 sky130_fd_sc_hd__a22o_1 _11447_ (.A1(_04837_),
    .A2(net475),
    .B1(net275),
    .B2(\reg_module.gprf[957] ),
    .X(_05403_));
 sky130_fd_sc_hd__and2_1 _11448_ (.A(net1177),
    .B(_05403_),
    .X(_01059_));
 sky130_fd_sc_hd__a22o_1 _11449_ (.A1(_04839_),
    .A2(net480),
    .B1(net276),
    .B2(\reg_module.gprf[958] ),
    .X(_05404_));
 sky130_fd_sc_hd__and2_1 _11450_ (.A(net1194),
    .B(_05404_),
    .X(_01060_));
 sky130_fd_sc_hd__a22o_1 _11451_ (.A1(_04841_),
    .A2(net485),
    .B1(net276),
    .B2(\reg_module.gprf[959] ),
    .X(_05405_));
 sky130_fd_sc_hd__and2_1 _11452_ (.A(net1205),
    .B(_05405_),
    .X(_01061_));
 sky130_fd_sc_hd__or2_4 _11453_ (.A(net632),
    .B(_04976_),
    .X(_05406_));
 sky130_fd_sc_hd__a22o_1 _11454_ (.A1(_04845_),
    .A2(net453),
    .B1(net270),
    .B2(\reg_module.gprf[960] ),
    .X(_05407_));
 sky130_fd_sc_hd__and2_1 _11455_ (.A(net1124),
    .B(_05407_),
    .X(_01062_));
 sky130_fd_sc_hd__a22o_1 _11456_ (.A1(_04847_),
    .A2(net457),
    .B1(net270),
    .B2(\reg_module.gprf[961] ),
    .X(_05408_));
 sky130_fd_sc_hd__and2_1 _11457_ (.A(net1132),
    .B(_05408_),
    .X(_01063_));
 sky130_fd_sc_hd__a22o_1 _11458_ (.A1(_04849_),
    .A2(net447),
    .B1(net269),
    .B2(\reg_module.gprf[962] ),
    .X(_05409_));
 sky130_fd_sc_hd__and2_1 _11459_ (.A(net1111),
    .B(_05409_),
    .X(_01064_));
 sky130_fd_sc_hd__a22o_1 _11460_ (.A1(_04851_),
    .A2(net441),
    .B1(net269),
    .B2(\reg_module.gprf[963] ),
    .X(_05410_));
 sky130_fd_sc_hd__and2_1 _11461_ (.A(net1090),
    .B(_05410_),
    .X(_01065_));
 sky130_fd_sc_hd__a22o_1 _11462_ (.A1(_04853_),
    .A2(net455),
    .B1(net270),
    .B2(\reg_module.gprf[964] ),
    .X(_05411_));
 sky130_fd_sc_hd__and2_1 _11463_ (.A(net1130),
    .B(_05411_),
    .X(_01066_));
 sky130_fd_sc_hd__a22o_1 _11464_ (.A1(_04855_),
    .A2(net452),
    .B1(net270),
    .B2(\reg_module.gprf[965] ),
    .X(_05412_));
 sky130_fd_sc_hd__and2_1 _11465_ (.A(net1120),
    .B(_05412_),
    .X(_01067_));
 sky130_fd_sc_hd__a22o_1 _11466_ (.A1(_04857_),
    .A2(net439),
    .B1(net269),
    .B2(\reg_module.gprf[966] ),
    .X(_05413_));
 sky130_fd_sc_hd__and2_1 _11467_ (.A(net1082),
    .B(_05413_),
    .X(_01068_));
 sky130_fd_sc_hd__a22o_1 _11468_ (.A1(_04859_),
    .A2(net438),
    .B1(net269),
    .B2(\reg_module.gprf[967] ),
    .X(_05414_));
 sky130_fd_sc_hd__and2_1 _11469_ (.A(net1086),
    .B(_05414_),
    .X(_01069_));
 sky130_fd_sc_hd__a22o_1 _11470_ (.A1(_04861_),
    .A2(net454),
    .B1(net270),
    .B2(\reg_module.gprf[968] ),
    .X(_05415_));
 sky130_fd_sc_hd__and2_1 _11471_ (.A(net1123),
    .B(_05415_),
    .X(_01070_));
 sky130_fd_sc_hd__a22o_1 _11472_ (.A1(_04863_),
    .A2(net435),
    .B1(net269),
    .B2(\reg_module.gprf[969] ),
    .X(_05416_));
 sky130_fd_sc_hd__and2_1 _11473_ (.A(net1075),
    .B(_05416_),
    .X(_01071_));
 sky130_fd_sc_hd__a22o_1 _11474_ (.A1(_04865_),
    .A2(net433),
    .B1(net269),
    .B2(\reg_module.gprf[970] ),
    .X(_05417_));
 sky130_fd_sc_hd__and2_1 _11475_ (.A(net1080),
    .B(_05417_),
    .X(_01072_));
 sky130_fd_sc_hd__a22o_1 _11476_ (.A1(_04867_),
    .A2(net443),
    .B1(net269),
    .B2(\reg_module.gprf[971] ),
    .X(_05418_));
 sky130_fd_sc_hd__and2_1 _11477_ (.A(net1095),
    .B(_05418_),
    .X(_01073_));
 sky130_fd_sc_hd__a22o_1 _11478_ (.A1(_04869_),
    .A2(net466),
    .B1(net271),
    .B2(\reg_module.gprf[972] ),
    .X(_05419_));
 sky130_fd_sc_hd__and2_1 _11479_ (.A(net1152),
    .B(_05419_),
    .X(_01074_));
 sky130_fd_sc_hd__a22o_1 _11480_ (.A1(_04871_),
    .A2(net443),
    .B1(net269),
    .B2(\reg_module.gprf[973] ),
    .X(_05420_));
 sky130_fd_sc_hd__and2_1 _11481_ (.A(net1098),
    .B(_05420_),
    .X(_01075_));
 sky130_fd_sc_hd__a22o_1 _11482_ (.A1(_04873_),
    .A2(net465),
    .B1(net269),
    .B2(\reg_module.gprf[974] ),
    .X(_05421_));
 sky130_fd_sc_hd__and2_1 _11483_ (.A(net1157),
    .B(_05421_),
    .X(_01076_));
 sky130_fd_sc_hd__a22o_1 _11484_ (.A1(_04875_),
    .A2(net468),
    .B1(net271),
    .B2(\reg_module.gprf[975] ),
    .X(_05422_));
 sky130_fd_sc_hd__and2_1 _11485_ (.A(net1161),
    .B(_05422_),
    .X(_01077_));
 sky130_fd_sc_hd__a22o_1 _11486_ (.A1(_04877_),
    .A2(net484),
    .B1(net272),
    .B2(\reg_module.gprf[976] ),
    .X(_05423_));
 sky130_fd_sc_hd__and2_1 _11487_ (.A(net1202),
    .B(_05423_),
    .X(_01078_));
 sky130_fd_sc_hd__a22o_1 _11488_ (.A1(_04879_),
    .A2(net462),
    .B1(net271),
    .B2(\reg_module.gprf[977] ),
    .X(_05424_));
 sky130_fd_sc_hd__and2_1 _11489_ (.A(net1147),
    .B(_05424_),
    .X(_01079_));
 sky130_fd_sc_hd__a22o_1 _11490_ (.A1(_04881_),
    .A2(net445),
    .B1(net270),
    .B2(\reg_module.gprf[978] ),
    .X(_05425_));
 sky130_fd_sc_hd__and2_1 _11491_ (.A(net1101),
    .B(_05425_),
    .X(_01080_));
 sky130_fd_sc_hd__a22o_1 _11492_ (.A1(_04883_),
    .A2(net467),
    .B1(net271),
    .B2(\reg_module.gprf[979] ),
    .X(_05426_));
 sky130_fd_sc_hd__and2_1 _11493_ (.A(net1158),
    .B(_05426_),
    .X(_01081_));
 sky130_fd_sc_hd__a22o_1 _11494_ (.A1(_04885_),
    .A2(net466),
    .B1(net269),
    .B2(\reg_module.gprf[980] ),
    .X(_05427_));
 sky130_fd_sc_hd__and2_1 _11495_ (.A(net1154),
    .B(_05427_),
    .X(_01082_));
 sky130_fd_sc_hd__a22o_1 _11496_ (.A1(_04887_),
    .A2(net486),
    .B1(net272),
    .B2(\reg_module.gprf[981] ),
    .X(_05428_));
 sky130_fd_sc_hd__and2_1 _11497_ (.A(net1207),
    .B(_05428_),
    .X(_01083_));
 sky130_fd_sc_hd__a22o_1 _11498_ (.A1(_04889_),
    .A2(net481),
    .B1(net272),
    .B2(\reg_module.gprf[982] ),
    .X(_05429_));
 sky130_fd_sc_hd__and2_1 _11499_ (.A(net1197),
    .B(_05429_),
    .X(_01084_));
 sky130_fd_sc_hd__a22o_1 _11500_ (.A1(_04891_),
    .A2(net472),
    .B1(net271),
    .B2(\reg_module.gprf[983] ),
    .X(_05430_));
 sky130_fd_sc_hd__and2_1 _11501_ (.A(net1164),
    .B(_05430_),
    .X(_01085_));
 sky130_fd_sc_hd__a22o_1 _11502_ (.A1(_04893_),
    .A2(net478),
    .B1(net271),
    .B2(\reg_module.gprf[984] ),
    .X(_05431_));
 sky130_fd_sc_hd__and2_1 _11503_ (.A(net1183),
    .B(_05431_),
    .X(_01086_));
 sky130_fd_sc_hd__a22o_1 _11504_ (.A1(_04895_),
    .A2(net477),
    .B1(net271),
    .B2(\reg_module.gprf[985] ),
    .X(_05432_));
 sky130_fd_sc_hd__and2_1 _11505_ (.A(net1180),
    .B(_05432_),
    .X(_01087_));
 sky130_fd_sc_hd__a22o_1 _11506_ (.A1(_04897_),
    .A2(net476),
    .B1(net271),
    .B2(\reg_module.gprf[986] ),
    .X(_05433_));
 sky130_fd_sc_hd__and2_1 _11507_ (.A(net1178),
    .B(_05433_),
    .X(_01088_));
 sky130_fd_sc_hd__a22o_1 _11508_ (.A1(_04899_),
    .A2(net462),
    .B1(net271),
    .B2(\reg_module.gprf[987] ),
    .X(_05434_));
 sky130_fd_sc_hd__and2_1 _11509_ (.A(net1146),
    .B(_05434_),
    .X(_01089_));
 sky130_fd_sc_hd__a22o_1 _11510_ (.A1(_04901_),
    .A2(net473),
    .B1(net271),
    .B2(\reg_module.gprf[988] ),
    .X(_05435_));
 sky130_fd_sc_hd__and2_1 _11511_ (.A(net1172),
    .B(_05435_),
    .X(_01090_));
 sky130_fd_sc_hd__a22o_1 _11512_ (.A1(_04903_),
    .A2(net475),
    .B1(net272),
    .B2(\reg_module.gprf[989] ),
    .X(_05436_));
 sky130_fd_sc_hd__and2_1 _11513_ (.A(net1177),
    .B(_05436_),
    .X(_01091_));
 sky130_fd_sc_hd__a22o_1 _11514_ (.A1(_04905_),
    .A2(net480),
    .B1(net272),
    .B2(\reg_module.gprf[990] ),
    .X(_05437_));
 sky130_fd_sc_hd__and2_1 _11515_ (.A(net1194),
    .B(_05437_),
    .X(_01092_));
 sky130_fd_sc_hd__a22o_1 _11516_ (.A1(_04907_),
    .A2(net485),
    .B1(net272),
    .B2(\reg_module.gprf[991] ),
    .X(_05438_));
 sky130_fd_sc_hd__and2_1 _11517_ (.A(net1205),
    .B(_05438_),
    .X(_01093_));
 sky130_fd_sc_hd__and2_1 _11518_ (.A(net1258),
    .B(net1125),
    .X(_01094_));
 sky130_fd_sc_hd__and2_1 _11519_ (.A(net1279),
    .B(net1133),
    .X(_01095_));
 sky130_fd_sc_hd__and2_1 _11520_ (.A(net1283),
    .B(net1111),
    .X(_01096_));
 sky130_fd_sc_hd__and2_1 _11521_ (.A(net1269),
    .B(net1090),
    .X(_01097_));
 sky130_fd_sc_hd__and2_1 _11522_ (.A(net1292),
    .B(net1131),
    .X(_01098_));
 sky130_fd_sc_hd__and2_1 _11523_ (.A(net1266),
    .B(net1123),
    .X(_01099_));
 sky130_fd_sc_hd__and2_1 _11524_ (.A(net1289),
    .B(net1082),
    .X(_01100_));
 sky130_fd_sc_hd__and2_1 _11525_ (.A(net1254),
    .B(net1093),
    .X(_01101_));
 sky130_fd_sc_hd__and2_1 _11526_ (.A(net1290),
    .B(net1134),
    .X(_01102_));
 sky130_fd_sc_hd__and2_1 _11527_ (.A(net1262),
    .B(net1075),
    .X(_01103_));
 sky130_fd_sc_hd__and2_1 _11528_ (.A(net1280),
    .B(net1073),
    .X(_01104_));
 sky130_fd_sc_hd__and2_1 _11529_ (.A(net1270),
    .B(net1095),
    .X(_01105_));
 sky130_fd_sc_hd__and2_1 _11530_ (.A(net1276),
    .B(net1153),
    .X(_01106_));
 sky130_fd_sc_hd__and2_1 _11531_ (.A(net1268),
    .B(net1097),
    .X(_01107_));
 sky130_fd_sc_hd__and2_1 _11532_ (.A(net1274),
    .B(net1117),
    .X(_01108_));
 sky130_fd_sc_hd__and2_1 _11533_ (.A(net1291),
    .B(net1156),
    .X(_01109_));
 sky130_fd_sc_hd__and2_1 _11534_ (.A(net1286),
    .B(net1202),
    .X(_01110_));
 sky130_fd_sc_hd__and2_1 _11535_ (.A(net1272),
    .B(net1145),
    .X(_01111_));
 sky130_fd_sc_hd__and2_1 _11536_ (.A(net1273),
    .B(net1101),
    .X(_01112_));
 sky130_fd_sc_hd__and2_1 _11537_ (.A(net1288),
    .B(net1158),
    .X(_01113_));
 sky130_fd_sc_hd__and2_1 _11538_ (.A(net1271),
    .B(net1154),
    .X(_01114_));
 sky130_fd_sc_hd__and2_1 _11539_ (.A(net1267),
    .B(net1207),
    .X(_01115_));
 sky130_fd_sc_hd__and2_1 _11540_ (.A(net1261),
    .B(net1197),
    .X(_01116_));
 sky130_fd_sc_hd__and2_1 _11541_ (.A(net1260),
    .B(net1164),
    .X(_01117_));
 sky130_fd_sc_hd__and2_1 _11542_ (.A(net1298),
    .B(net1183),
    .X(_01118_));
 sky130_fd_sc_hd__and2_1 _11543_ (.A(net1257),
    .B(net1180),
    .X(_01119_));
 sky130_fd_sc_hd__and2_1 _11544_ (.A(net1253),
    .B(net1178),
    .X(_01120_));
 sky130_fd_sc_hd__and2_1 _11545_ (.A(net1263),
    .B(net1146),
    .X(_01121_));
 sky130_fd_sc_hd__and2_1 _11546_ (.A(net1287),
    .B(net1172),
    .X(_01122_));
 sky130_fd_sc_hd__and2_1 _11547_ (.A(net1275),
    .B(net1177),
    .X(_01123_));
 sky130_fd_sc_hd__and2_1 _11548_ (.A(net1264),
    .B(net1193),
    .X(_01124_));
 sky130_fd_sc_hd__and2_1 _11549_ (.A(net1265),
    .B(net1206),
    .X(_01125_));
 sky130_fd_sc_hd__or2_1 _11550_ (.A(\brancher.imm12_i_s[2] ),
    .B(_01326_),
    .X(_05439_));
 sky130_fd_sc_hd__nand2_1 _11551_ (.A(\brancher.imm12_i_s[2] ),
    .B(_01326_),
    .Y(_05440_));
 sky130_fd_sc_hd__nand2_1 _11552_ (.A(_05439_),
    .B(_05440_),
    .Y(_05441_));
 sky130_fd_sc_hd__nand2_1 _11553_ (.A(\brancher.imm12_i_s[1] ),
    .B(_01302_),
    .Y(_05442_));
 sky130_fd_sc_hd__xnor2_1 _11554_ (.A(\brancher.imm12_i_s[1] ),
    .B(_01302_),
    .Y(_05443_));
 sky130_fd_sc_hd__nand2_1 _11555_ (.A(\brancher.imm12_i_s[0] ),
    .B(_01279_),
    .Y(_05444_));
 sky130_fd_sc_hd__or2_1 _11556_ (.A(_05443_),
    .B(_05444_),
    .X(_05445_));
 sky130_fd_sc_hd__o21a_1 _11557_ (.A1(_05443_),
    .A2(_05444_),
    .B1(_05442_),
    .X(_05446_));
 sky130_fd_sc_hd__nand2_4 _11558_ (.A(net836),
    .B(net956),
    .Y(_05447_));
 sky130_fd_sc_hd__a21oi_1 _11559_ (.A1(_05441_),
    .A2(_05446_),
    .B1(_05447_),
    .Y(_05448_));
 sky130_fd_sc_hd__o21ai_1 _11560_ (.A1(_05441_),
    .A2(_05446_),
    .B1(_05448_),
    .Y(_05449_));
 sky130_fd_sc_hd__or2_1 _11561_ (.A(net882),
    .B(\brancher.rPc_current_reg2[2] ),
    .X(_05450_));
 sky130_fd_sc_hd__nand2_1 _11562_ (.A(net882),
    .B(\brancher.rPc_current_reg2[2] ),
    .Y(_05451_));
 sky130_fd_sc_hd__and2_1 _11563_ (.A(net1),
    .B(net268),
    .X(_05452_));
 sky130_fd_sc_hd__nand2_2 _11564_ (.A(net1),
    .B(net268),
    .Y(_05453_));
 sky130_fd_sc_hd__nor2_2 _11565_ (.A(\alu.b_type ),
    .B(_03218_),
    .Y(_05454_));
 sky130_fd_sc_hd__nand2_2 _11566_ (.A(_01209_),
    .B(_03217_),
    .Y(_05455_));
 sky130_fd_sc_hd__nor2_2 _11567_ (.A(net201),
    .B(net630),
    .Y(_05456_));
 sky130_fd_sc_hd__nand2_1 _11568_ (.A(_05449_),
    .B(net184),
    .Y(_05457_));
 sky130_fd_sc_hd__a31o_1 _11569_ (.A1(net953),
    .A2(_05450_),
    .A3(_05451_),
    .B1(_05457_),
    .X(_05458_));
 sky130_fd_sc_hd__nand2_1 _11570_ (.A(\brancher.imm13_b[1] ),
    .B(\brancher.rPc_current_reg2[2] ),
    .Y(_05459_));
 sky130_fd_sc_hd__o21a_1 _11571_ (.A1(\brancher.imm13_b[1] ),
    .A2(\brancher.rPc_current_reg2[2] ),
    .B1(_03217_),
    .X(_05460_));
 sky130_fd_sc_hd__a31o_1 _11572_ (.A1(net176),
    .A2(_05459_),
    .A3(_05460_),
    .B1(_05458_),
    .X(_05461_));
 sky130_fd_sc_hd__o21bai_1 _11573_ (.A1(net157),
    .A2(_04046_),
    .B1_N(_05461_),
    .Y(_05462_));
 sky130_fd_sc_hd__nor2_4 _11574_ (.A(net201),
    .B(net628),
    .Y(_05463_));
 sky130_fd_sc_hd__nand2_1 _11575_ (.A(net157),
    .B(_05463_),
    .Y(_05464_));
 sky130_fd_sc_hd__o2111a_1 _11576_ (.A1(net157),
    .A2(net204),
    .B1(_05462_),
    .C1(_05464_),
    .D1(net1137),
    .X(_01126_));
 sky130_fd_sc_hd__and2_1 _11577_ (.A(\brancher.imm13_b[2] ),
    .B(\brancher.rPc_current_reg2[3] ),
    .X(_05465_));
 sky130_fd_sc_hd__nor2_1 _11578_ (.A(\brancher.imm13_b[2] ),
    .B(\brancher.rPc_current_reg2[3] ),
    .Y(_05466_));
 sky130_fd_sc_hd__nor2_1 _11579_ (.A(_05465_),
    .B(_05466_),
    .Y(_05467_));
 sky130_fd_sc_hd__xor2_1 _11580_ (.A(_05459_),
    .B(_05467_),
    .X(_05468_));
 sky130_fd_sc_hd__xor2_1 _11581_ (.A(net160),
    .B(net157),
    .X(_05469_));
 sky130_fd_sc_hd__nor2_1 _11582_ (.A(net174),
    .B(_05469_),
    .Y(_05470_));
 sky130_fd_sc_hd__a21o_1 _11583_ (.A1(net175),
    .A2(_05468_),
    .B1(net957),
    .X(_05471_));
 sky130_fd_sc_hd__nand2_1 _11584_ (.A(\brancher.imm12_i_s[3] ),
    .B(_01346_),
    .Y(_05472_));
 sky130_fd_sc_hd__or2_1 _11585_ (.A(\brancher.imm12_i_s[3] ),
    .B(_01346_),
    .X(_05473_));
 sky130_fd_sc_hd__nand2_1 _11586_ (.A(_05472_),
    .B(_05473_),
    .Y(_05474_));
 sky130_fd_sc_hd__o21a_1 _11587_ (.A1(_05441_),
    .A2(_05446_),
    .B1(_05440_),
    .X(_05475_));
 sky130_fd_sc_hd__o21ai_1 _11588_ (.A1(_05474_),
    .A2(_05475_),
    .B1(net957),
    .Y(_05476_));
 sky130_fd_sc_hd__a21o_1 _11589_ (.A1(_05474_),
    .A2(_05475_),
    .B1(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__o211ai_1 _11590_ (.A1(_05470_),
    .A2(_05471_),
    .B1(_05477_),
    .C1(net836),
    .Y(_05478_));
 sky130_fd_sc_hd__and2_1 _11591_ (.A(net861),
    .B(\brancher.rPc_current_reg2[3] ),
    .X(_05479_));
 sky130_fd_sc_hd__xor2_1 _11592_ (.A(net861),
    .B(\brancher.rPc_current_reg2[3] ),
    .X(_05480_));
 sky130_fd_sc_hd__a21oi_1 _11593_ (.A1(net882),
    .A2(\brancher.rPc_current_reg2[2] ),
    .B1(_05480_),
    .Y(_05481_));
 sky130_fd_sc_hd__and3_1 _11594_ (.A(net882),
    .B(\brancher.rPc_current_reg2[2] ),
    .C(_05480_),
    .X(_05482_));
 sky130_fd_sc_hd__o21ai_1 _11595_ (.A1(_05481_),
    .A2(_05482_),
    .B1(net953),
    .Y(_05483_));
 sky130_fd_sc_hd__and3_1 _11596_ (.A(net184),
    .B(_05478_),
    .C(_05483_),
    .X(_05484_));
 sky130_fd_sc_hd__a22o_1 _11597_ (.A1(net160),
    .A2(net201),
    .B1(_05463_),
    .B2(_05469_),
    .X(_05485_));
 sky130_fd_sc_hd__o21a_1 _11598_ (.A1(_05484_),
    .A2(_05485_),
    .B1(net1135),
    .X(_01127_));
 sky130_fd_sc_hd__or2_1 _11599_ (.A(\brancher.imm13_b[3] ),
    .B(\brancher.rPc_current_reg2[4] ),
    .X(_05486_));
 sky130_fd_sc_hd__nand2_1 _11600_ (.A(\brancher.imm13_b[3] ),
    .B(\brancher.rPc_current_reg2[4] ),
    .Y(_05487_));
 sky130_fd_sc_hd__nand2_1 _11601_ (.A(_05486_),
    .B(_05487_),
    .Y(_05488_));
 sky130_fd_sc_hd__a31o_1 _11602_ (.A1(\brancher.imm13_b[1] ),
    .A2(\brancher.rPc_current_reg2[2] ),
    .A3(_05467_),
    .B1(_05465_),
    .X(_05489_));
 sky130_fd_sc_hd__xnor2_1 _11603_ (.A(_05488_),
    .B(_05489_),
    .Y(_05490_));
 sky130_fd_sc_hd__and3_1 _11604_ (.A(net161),
    .B(net160),
    .C(net157),
    .X(_05491_));
 sky130_fd_sc_hd__a21oi_1 _11605_ (.A1(net160),
    .A2(net157),
    .B1(net161),
    .Y(_05492_));
 sky130_fd_sc_hd__nor2_1 _11606_ (.A(_05491_),
    .B(_05492_),
    .Y(_05493_));
 sky130_fd_sc_hd__mux2_1 _11607_ (.A0(_05493_),
    .A1(_05490_),
    .S(net176),
    .X(_05494_));
 sky130_fd_sc_hd__and2_1 _11608_ (.A(\brancher.imm12_i_s[4] ),
    .B(_01367_),
    .X(_05495_));
 sky130_fd_sc_hd__nor2_1 _11609_ (.A(\brancher.imm12_i_s[4] ),
    .B(_01367_),
    .Y(_05496_));
 sky130_fd_sc_hd__or2_1 _11610_ (.A(_05495_),
    .B(_05496_),
    .X(_05497_));
 sky130_fd_sc_hd__inv_2 _11611_ (.A(_05497_),
    .Y(_05498_));
 sky130_fd_sc_hd__o21ai_1 _11612_ (.A1(_05474_),
    .A2(_05475_),
    .B1(_05472_),
    .Y(_05499_));
 sky130_fd_sc_hd__and2_1 _11613_ (.A(_05498_),
    .B(_05499_),
    .X(_05500_));
 sky130_fd_sc_hd__o21ai_1 _11614_ (.A1(_05498_),
    .A2(_05499_),
    .B1(net957),
    .Y(_05501_));
 sky130_fd_sc_hd__nor2_1 _11615_ (.A(_05500_),
    .B(_05501_),
    .Y(_05502_));
 sky130_fd_sc_hd__a211o_1 _11616_ (.A1(_01208_),
    .A2(_05494_),
    .B1(_05502_),
    .C1(net952),
    .X(_05503_));
 sky130_fd_sc_hd__or2_1 _11617_ (.A(net851),
    .B(\brancher.rPc_current_reg2[4] ),
    .X(_05504_));
 sky130_fd_sc_hd__nand2_1 _11618_ (.A(net851),
    .B(\brancher.rPc_current_reg2[4] ),
    .Y(_05505_));
 sky130_fd_sc_hd__a31o_1 _11619_ (.A1(net882),
    .A2(\brancher.rPc_current_reg2[2] ),
    .A3(_05480_),
    .B1(_05479_),
    .X(_05506_));
 sky130_fd_sc_hd__and3_1 _11620_ (.A(_05504_),
    .B(_05505_),
    .C(_05506_),
    .X(_05507_));
 sky130_fd_sc_hd__a21oi_1 _11621_ (.A1(_05504_),
    .A2(_05505_),
    .B1(_05506_),
    .Y(_05508_));
 sky130_fd_sc_hd__o21ai_1 _11622_ (.A1(_05507_),
    .A2(_05508_),
    .B1(net953),
    .Y(_05509_));
 sky130_fd_sc_hd__and3_1 _11623_ (.A(net184),
    .B(_05503_),
    .C(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__a22o_1 _11624_ (.A1(net161),
    .A2(net201),
    .B1(_05463_),
    .B2(_05493_),
    .X(_05511_));
 sky130_fd_sc_hd__o21a_1 _11625_ (.A1(_05510_),
    .A2(_05511_),
    .B1(net1137),
    .X(_01128_));
 sky130_fd_sc_hd__or2_1 _11626_ (.A(\brancher.imm13_b[4] ),
    .B(\brancher.rPc_current_reg2[5] ),
    .X(_05512_));
 sky130_fd_sc_hd__nand2_1 _11627_ (.A(\brancher.imm13_b[4] ),
    .B(\brancher.rPc_current_reg2[5] ),
    .Y(_05513_));
 sky130_fd_sc_hd__nand2_1 _11628_ (.A(_05512_),
    .B(_05513_),
    .Y(_05514_));
 sky130_fd_sc_hd__a21bo_1 _11629_ (.A1(_05486_),
    .A2(_05489_),
    .B1_N(_05487_),
    .X(_05515_));
 sky130_fd_sc_hd__xnor2_1 _11630_ (.A(_05514_),
    .B(_05515_),
    .Y(_05516_));
 sky130_fd_sc_hd__and2_1 _11631_ (.A(net162),
    .B(_05491_),
    .X(_05517_));
 sky130_fd_sc_hd__nor2_1 _11632_ (.A(net162),
    .B(_05491_),
    .Y(_05518_));
 sky130_fd_sc_hd__nor2_1 _11633_ (.A(_05517_),
    .B(_05518_),
    .Y(_05519_));
 sky130_fd_sc_hd__mux2_1 _11634_ (.A0(_05519_),
    .A1(_05516_),
    .S(net174),
    .X(_05520_));
 sky130_fd_sc_hd__nor2_1 _11635_ (.A(_05495_),
    .B(_05500_),
    .Y(_05521_));
 sky130_fd_sc_hd__and2_1 _11636_ (.A(\brancher.imm12_i_s[5] ),
    .B(_01389_),
    .X(_05522_));
 sky130_fd_sc_hd__nor2_1 _11637_ (.A(\brancher.imm12_i_s[5] ),
    .B(_01389_),
    .Y(_05523_));
 sky130_fd_sc_hd__inv_2 _11638_ (.A(_05523_),
    .Y(_05524_));
 sky130_fd_sc_hd__or3_1 _11639_ (.A(_05521_),
    .B(_05522_),
    .C(_05523_),
    .X(_05525_));
 sky130_fd_sc_hd__o21ai_1 _11640_ (.A1(_05522_),
    .A2(_05523_),
    .B1(_05521_),
    .Y(_05526_));
 sky130_fd_sc_hd__a31o_1 _11641_ (.A1(net956),
    .A2(_05525_),
    .A3(_05526_),
    .B1(net952),
    .X(_05527_));
 sky130_fd_sc_hd__a21o_1 _11642_ (.A1(_01208_),
    .A2(_05520_),
    .B1(_05527_),
    .X(_05528_));
 sky130_fd_sc_hd__or2_1 _11643_ (.A(net940),
    .B(\brancher.rPc_current_reg2[5] ),
    .X(_05529_));
 sky130_fd_sc_hd__nand2_1 _11644_ (.A(net940),
    .B(\brancher.rPc_current_reg2[5] ),
    .Y(_05530_));
 sky130_fd_sc_hd__nand2_1 _11645_ (.A(_05529_),
    .B(_05530_),
    .Y(_05531_));
 sky130_fd_sc_hd__a21bo_1 _11646_ (.A1(_05504_),
    .A2(_05506_),
    .B1_N(_05505_),
    .X(_05532_));
 sky130_fd_sc_hd__xnor2_1 _11647_ (.A(_05531_),
    .B(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__o211a_1 _11648_ (.A1(net836),
    .A2(_05533_),
    .B1(_05528_),
    .C1(net184),
    .X(_05534_));
 sky130_fd_sc_hd__a22o_1 _11649_ (.A1(net162),
    .A2(net201),
    .B1(_05463_),
    .B2(_05519_),
    .X(_05535_));
 sky130_fd_sc_hd__o21a_1 _11650_ (.A1(_05534_),
    .A2(_05535_),
    .B1(net1135),
    .X(_01129_));
 sky130_fd_sc_hd__xnor2_1 _11651_ (.A(net163),
    .B(_05517_),
    .Y(_05536_));
 sky130_fd_sc_hd__and2_1 _11652_ (.A(\brancher.imm13_b[5] ),
    .B(\brancher.rPc_current_reg2[6] ),
    .X(_05537_));
 sky130_fd_sc_hd__nor2_1 _11653_ (.A(\brancher.imm13_b[5] ),
    .B(\brancher.rPc_current_reg2[6] ),
    .Y(_05538_));
 sky130_fd_sc_hd__or2_2 _11654_ (.A(_05537_),
    .B(_05538_),
    .X(_05539_));
 sky130_fd_sc_hd__a21boi_2 _11655_ (.A1(_05512_),
    .A2(_05515_),
    .B1_N(_05513_),
    .Y(_05540_));
 sky130_fd_sc_hd__xnor2_1 _11656_ (.A(_05539_),
    .B(_05540_),
    .Y(_05541_));
 sky130_fd_sc_hd__mux2_1 _11657_ (.A0(_05536_),
    .A1(_05541_),
    .S(net174),
    .X(_05542_));
 sky130_fd_sc_hd__nor2_1 _11658_ (.A(_01226_),
    .B(_01412_),
    .Y(_05543_));
 sky130_fd_sc_hd__nand2_1 _11659_ (.A(_01226_),
    .B(_01412_),
    .Y(_05544_));
 sky130_fd_sc_hd__nand2b_1 _11660_ (.A_N(_05543_),
    .B(_05544_),
    .Y(_05545_));
 sky130_fd_sc_hd__a211o_1 _11661_ (.A1(_05498_),
    .A2(_05499_),
    .B1(_05522_),
    .C1(_05495_),
    .X(_05546_));
 sky130_fd_sc_hd__nand2_1 _11662_ (.A(_05524_),
    .B(_05546_),
    .Y(_05547_));
 sky130_fd_sc_hd__xnor2_1 _11663_ (.A(_05545_),
    .B(_05547_),
    .Y(_05548_));
 sky130_fd_sc_hd__mux2_1 _11664_ (.A0(_05542_),
    .A1(_05548_),
    .S(net956),
    .X(_05549_));
 sky130_fd_sc_hd__nand2_1 _11665_ (.A(net836),
    .B(_05549_),
    .Y(_05550_));
 sky130_fd_sc_hd__a21boi_1 _11666_ (.A1(_05529_),
    .A2(_05532_),
    .B1_N(_05530_),
    .Y(_05551_));
 sky130_fd_sc_hd__nor2_1 _11667_ (.A(_05539_),
    .B(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__nand2_1 _11668_ (.A(_05539_),
    .B(_05551_),
    .Y(_05553_));
 sky130_fd_sc_hd__and2b_1 _11669_ (.A_N(_05552_),
    .B(_05553_),
    .X(_05554_));
 sky130_fd_sc_hd__o211a_1 _11670_ (.A1(net836),
    .A2(_05554_),
    .B1(_05550_),
    .C1(net184),
    .X(_05555_));
 sky130_fd_sc_hd__nor2_1 _11671_ (.A(net628),
    .B(_05536_),
    .Y(_05556_));
 sky130_fd_sc_hd__mux2_1 _11672_ (.A0(net163),
    .A1(_05556_),
    .S(net204),
    .X(_05557_));
 sky130_fd_sc_hd__o21a_1 _11673_ (.A1(_05555_),
    .A2(_05557_),
    .B1(net1135),
    .X(_01130_));
 sky130_fd_sc_hd__and2_1 _11674_ (.A(\brancher.imm13_b[6] ),
    .B(\brancher.rPc_current_reg2[7] ),
    .X(_05558_));
 sky130_fd_sc_hd__or2_1 _11675_ (.A(\brancher.imm13_b[6] ),
    .B(\brancher.rPc_current_reg2[7] ),
    .X(_05559_));
 sky130_fd_sc_hd__and2b_1 _11676_ (.A_N(_05558_),
    .B(_05559_),
    .X(_05560_));
 sky130_fd_sc_hd__inv_2 _11677_ (.A(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__o21ba_1 _11678_ (.A1(_05539_),
    .A2(_05540_),
    .B1_N(_05537_),
    .X(_05562_));
 sky130_fd_sc_hd__xnor2_1 _11679_ (.A(_05560_),
    .B(_05562_),
    .Y(_05563_));
 sky130_fd_sc_hd__and3_1 _11680_ (.A(net164),
    .B(net163),
    .C(_05517_),
    .X(_05564_));
 sky130_fd_sc_hd__a21oi_1 _11681_ (.A1(net163),
    .A2(_05517_),
    .B1(net164),
    .Y(_05565_));
 sky130_fd_sc_hd__nor2_1 _11682_ (.A(_05564_),
    .B(_05565_),
    .Y(_05566_));
 sky130_fd_sc_hd__mux2_1 _11683_ (.A0(_05566_),
    .A1(_05563_),
    .S(net174),
    .X(_05567_));
 sky130_fd_sc_hd__nor2_1 _11684_ (.A(_01225_),
    .B(_01437_),
    .Y(_05568_));
 sky130_fd_sc_hd__nand2_1 _11685_ (.A(_01225_),
    .B(_01437_),
    .Y(_05569_));
 sky130_fd_sc_hd__nand2b_1 _11686_ (.A_N(_05568_),
    .B(_05569_),
    .Y(_05570_));
 sky130_fd_sc_hd__a31o_1 _11687_ (.A1(_05524_),
    .A2(_05544_),
    .A3(_05546_),
    .B1(_05543_),
    .X(_05571_));
 sky130_fd_sc_hd__xnor2_1 _11688_ (.A(_05570_),
    .B(_05571_),
    .Y(_05572_));
 sky130_fd_sc_hd__and3_1 _11689_ (.A(net836),
    .B(net956),
    .C(_05572_),
    .X(_05573_));
 sky130_fd_sc_hd__o21ai_1 _11690_ (.A1(_05537_),
    .A2(_05552_),
    .B1(_05560_),
    .Y(_05574_));
 sky130_fd_sc_hd__or3_1 _11691_ (.A(_05537_),
    .B(_05552_),
    .C(_05560_),
    .X(_05575_));
 sky130_fd_sc_hd__and3_1 _11692_ (.A(net952),
    .B(_05574_),
    .C(_05575_),
    .X(_05576_));
 sky130_fd_sc_hd__a211o_1 _11693_ (.A1(_03217_),
    .A2(_05567_),
    .B1(_05573_),
    .C1(_05576_),
    .X(_05577_));
 sky130_fd_sc_hd__mux2_1 _11694_ (.A0(net164),
    .A1(_05577_),
    .S(net204),
    .X(_05578_));
 sky130_fd_sc_hd__and2_1 _11695_ (.A(net1135),
    .B(_05578_),
    .X(_01131_));
 sky130_fd_sc_hd__and2_1 _11696_ (.A(net165),
    .B(_05564_),
    .X(_05579_));
 sky130_fd_sc_hd__inv_2 _11697_ (.A(_05579_),
    .Y(_05580_));
 sky130_fd_sc_hd__or2_1 _11698_ (.A(net165),
    .B(_05564_),
    .X(_05581_));
 sky130_fd_sc_hd__nand2_1 _11699_ (.A(_05580_),
    .B(_05581_),
    .Y(_05582_));
 sky130_fd_sc_hd__and2_1 _11700_ (.A(\brancher.imm13_b[7] ),
    .B(\brancher.rPc_current_reg2[8] ),
    .X(_05583_));
 sky130_fd_sc_hd__nand2_1 _11701_ (.A(\brancher.imm13_b[7] ),
    .B(\brancher.rPc_current_reg2[8] ),
    .Y(_05584_));
 sky130_fd_sc_hd__nor2_1 _11702_ (.A(\brancher.imm13_b[7] ),
    .B(\brancher.rPc_current_reg2[8] ),
    .Y(_05585_));
 sky130_fd_sc_hd__nor2_1 _11703_ (.A(_05583_),
    .B(_05585_),
    .Y(_05586_));
 sky130_fd_sc_hd__a31oi_2 _11704_ (.A1(\brancher.imm13_b[5] ),
    .A2(\brancher.rPc_current_reg2[6] ),
    .A3(_05559_),
    .B1(_05558_),
    .Y(_05587_));
 sky130_fd_sc_hd__o31ai_2 _11705_ (.A1(_05539_),
    .A2(_05540_),
    .A3(_05561_),
    .B1(_05587_),
    .Y(_05588_));
 sky130_fd_sc_hd__xnor2_1 _11706_ (.A(_05586_),
    .B(_05588_),
    .Y(_05589_));
 sky130_fd_sc_hd__mux2_1 _11707_ (.A0(_05582_),
    .A1(_05589_),
    .S(net174),
    .X(_05590_));
 sky130_fd_sc_hd__and2_1 _11708_ (.A(\brancher.imm12_i_s[8] ),
    .B(_01460_),
    .X(_05591_));
 sky130_fd_sc_hd__inv_2 _11709_ (.A(_05591_),
    .Y(_05592_));
 sky130_fd_sc_hd__nor2_1 _11710_ (.A(\brancher.imm12_i_s[8] ),
    .B(_01460_),
    .Y(_05593_));
 sky130_fd_sc_hd__or2_1 _11711_ (.A(_05591_),
    .B(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__a21oi_1 _11712_ (.A1(_05569_),
    .A2(_05571_),
    .B1(_05568_),
    .Y(_05595_));
 sky130_fd_sc_hd__nor2_1 _11713_ (.A(_05594_),
    .B(_05595_),
    .Y(_05596_));
 sky130_fd_sc_hd__a21o_1 _11714_ (.A1(_05594_),
    .A2(_05595_),
    .B1(_01208_),
    .X(_05597_));
 sky130_fd_sc_hd__o221a_1 _11715_ (.A1(net956),
    .A2(_05590_),
    .B1(_05596_),
    .B2(_05597_),
    .C1(net836),
    .X(_05598_));
 sky130_fd_sc_hd__o31a_1 _11716_ (.A1(_05539_),
    .A2(_05551_),
    .A3(_05561_),
    .B1(_05587_),
    .X(_05599_));
 sky130_fd_sc_hd__xor2_1 _11717_ (.A(_05586_),
    .B(_05599_),
    .X(_05600_));
 sky130_fd_sc_hd__a21oi_1 _11718_ (.A1(net952),
    .A2(_05600_),
    .B1(_05598_),
    .Y(_05601_));
 sky130_fd_sc_hd__a32o_1 _11719_ (.A1(_05463_),
    .A2(_05580_),
    .A3(_05581_),
    .B1(net201),
    .B2(net165),
    .X(_05602_));
 sky130_fd_sc_hd__a21o_1 _11720_ (.A1(net184),
    .A2(_05601_),
    .B1(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__and2_1 _11721_ (.A(net1135),
    .B(_05603_),
    .X(_01132_));
 sky130_fd_sc_hd__nand2_1 _11722_ (.A(net166),
    .B(net201),
    .Y(_05604_));
 sky130_fd_sc_hd__nor2_1 _11723_ (.A(\brancher.imm13_b[8] ),
    .B(\brancher.rPc_current_reg2[9] ),
    .Y(_05605_));
 sky130_fd_sc_hd__nand2_1 _11724_ (.A(\brancher.imm13_b[8] ),
    .B(\brancher.rPc_current_reg2[9] ),
    .Y(_05606_));
 sky130_fd_sc_hd__nand2b_2 _11725_ (.A_N(_05605_),
    .B(_05606_),
    .Y(_05607_));
 sky130_fd_sc_hd__inv_2 _11726_ (.A(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__a21oi_1 _11727_ (.A1(_05586_),
    .A2(_05588_),
    .B1(_05583_),
    .Y(_05609_));
 sky130_fd_sc_hd__xnor2_1 _11728_ (.A(_05607_),
    .B(_05609_),
    .Y(_05610_));
 sky130_fd_sc_hd__xnor2_1 _11729_ (.A(net166),
    .B(_05579_),
    .Y(_05611_));
 sky130_fd_sc_hd__mux2_1 _11730_ (.A0(_05611_),
    .A1(_05610_),
    .S(net174),
    .X(_05612_));
 sky130_fd_sc_hd__nor2_1 _11731_ (.A(_05591_),
    .B(_05596_),
    .Y(_05613_));
 sky130_fd_sc_hd__nand2_1 _11732_ (.A(_01224_),
    .B(_01485_),
    .Y(_05614_));
 sky130_fd_sc_hd__inv_2 _11733_ (.A(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__or2_1 _11734_ (.A(_01224_),
    .B(_01485_),
    .X(_05616_));
 sky130_fd_sc_hd__nand2_1 _11735_ (.A(_05614_),
    .B(_05616_),
    .Y(_05617_));
 sky130_fd_sc_hd__xnor2_1 _11736_ (.A(_05613_),
    .B(_05617_),
    .Y(_05618_));
 sky130_fd_sc_hd__o21a_1 _11737_ (.A1(_05585_),
    .A2(_05599_),
    .B1(_05584_),
    .X(_05619_));
 sky130_fd_sc_hd__xnor2_1 _11738_ (.A(_05607_),
    .B(_05619_),
    .Y(_05620_));
 sky130_fd_sc_hd__o22a_1 _11739_ (.A1(_05447_),
    .A2(_05618_),
    .B1(_05620_),
    .B2(net836),
    .X(_05621_));
 sky130_fd_sc_hd__o211a_1 _11740_ (.A1(_03218_),
    .A2(_05612_),
    .B1(_05621_),
    .C1(net628),
    .X(_05622_));
 sky130_fd_sc_hd__a211o_1 _11741_ (.A1(net630),
    .A2(_05611_),
    .B1(_05622_),
    .C1(net201),
    .X(_05623_));
 sky130_fd_sc_hd__a21boi_1 _11742_ (.A1(_05604_),
    .A2(_05623_),
    .B1_N(net1135),
    .Y(_01133_));
 sky130_fd_sc_hd__and3_1 _11743_ (.A(net136),
    .B(net166),
    .C(_05579_),
    .X(_05624_));
 sky130_fd_sc_hd__a21oi_1 _11744_ (.A1(net166),
    .A2(_05579_),
    .B1(net136),
    .Y(_05625_));
 sky130_fd_sc_hd__nor2_1 _11745_ (.A(_05624_),
    .B(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__and2_1 _11746_ (.A(\brancher.imm13_b[9] ),
    .B(\brancher.rPc_current_reg2[10] ),
    .X(_05627_));
 sky130_fd_sc_hd__nand2_1 _11747_ (.A(\brancher.imm13_b[9] ),
    .B(\brancher.rPc_current_reg2[10] ),
    .Y(_05628_));
 sky130_fd_sc_hd__or2_1 _11748_ (.A(\brancher.imm13_b[9] ),
    .B(\brancher.rPc_current_reg2[10] ),
    .X(_05629_));
 sky130_fd_sc_hd__nand2_1 _11749_ (.A(_05628_),
    .B(_05629_),
    .Y(_05630_));
 sky130_fd_sc_hd__a21oi_1 _11750_ (.A1(_05584_),
    .A2(_05606_),
    .B1(_05605_),
    .Y(_05631_));
 sky130_fd_sc_hd__a21o_1 _11751_ (.A1(_05584_),
    .A2(_05606_),
    .B1(_05605_),
    .X(_05632_));
 sky130_fd_sc_hd__a31o_1 _11752_ (.A1(_05586_),
    .A2(_05588_),
    .A3(_05608_),
    .B1(_05631_),
    .X(_05633_));
 sky130_fd_sc_hd__nand2b_1 _11753_ (.A_N(_05630_),
    .B(_05633_),
    .Y(_05634_));
 sky130_fd_sc_hd__xnor2_1 _11754_ (.A(_05630_),
    .B(_05633_),
    .Y(_05635_));
 sky130_fd_sc_hd__mux2_1 _11755_ (.A0(_05626_),
    .A1(_05635_),
    .S(net174),
    .X(_05636_));
 sky130_fd_sc_hd__or2_1 _11756_ (.A(_01223_),
    .B(_01509_),
    .X(_05637_));
 sky130_fd_sc_hd__nand2_1 _11757_ (.A(_01223_),
    .B(_01509_),
    .Y(_05638_));
 sky130_fd_sc_hd__nand2_1 _11758_ (.A(_05637_),
    .B(_05638_),
    .Y(_05639_));
 sky130_fd_sc_hd__o211a_1 _11759_ (.A1(_05594_),
    .A2(_05595_),
    .B1(_05616_),
    .C1(_05592_),
    .X(_05640_));
 sky130_fd_sc_hd__or2_1 _11760_ (.A(_05615_),
    .B(_05640_),
    .X(_05641_));
 sky130_fd_sc_hd__xor2_1 _11761_ (.A(_05639_),
    .B(_05641_),
    .X(_05642_));
 sky130_fd_sc_hd__mux2_1 _11762_ (.A0(_05636_),
    .A1(_05642_),
    .S(net956),
    .X(_05643_));
 sky130_fd_sc_hd__o41a_1 _11763_ (.A1(_05583_),
    .A2(_05585_),
    .A3(_05599_),
    .A4(_05607_),
    .B1(_05632_),
    .X(_05644_));
 sky130_fd_sc_hd__nor2_1 _11764_ (.A(_05630_),
    .B(_05644_),
    .Y(_05645_));
 sky130_fd_sc_hd__and2_1 _11765_ (.A(_05630_),
    .B(_05644_),
    .X(_05646_));
 sky130_fd_sc_hd__nor2_1 _11766_ (.A(_05645_),
    .B(_05646_),
    .Y(_05647_));
 sky130_fd_sc_hd__mux2_1 _11767_ (.A0(_05643_),
    .A1(_05647_),
    .S(net952),
    .X(_05648_));
 sky130_fd_sc_hd__a22o_1 _11768_ (.A1(net136),
    .A2(net201),
    .B1(_05463_),
    .B2(_05626_),
    .X(_05649_));
 sky130_fd_sc_hd__a21oi_1 _11769_ (.A1(net184),
    .A2(_05648_),
    .B1(_05649_),
    .Y(_05650_));
 sky130_fd_sc_hd__and2b_1 _11770_ (.A_N(_05650_),
    .B(net1135),
    .X(_01134_));
 sky130_fd_sc_hd__and2_1 _11771_ (.A(net137),
    .B(_05624_),
    .X(_05651_));
 sky130_fd_sc_hd__nor2_1 _11772_ (.A(net137),
    .B(_05624_),
    .Y(_05652_));
 sky130_fd_sc_hd__or2_1 _11773_ (.A(\brancher.imm13_b[10] ),
    .B(\brancher.rPc_current_reg2[11] ),
    .X(_05653_));
 sky130_fd_sc_hd__inv_2 _11774_ (.A(_05653_),
    .Y(_05654_));
 sky130_fd_sc_hd__nand2_1 _11775_ (.A(\brancher.imm13_b[10] ),
    .B(\brancher.rPc_current_reg2[11] ),
    .Y(_05655_));
 sky130_fd_sc_hd__and2_1 _11776_ (.A(_05653_),
    .B(_05655_),
    .X(_05656_));
 sky130_fd_sc_hd__and3_1 _11777_ (.A(_05628_),
    .B(_05634_),
    .C(_05656_),
    .X(_05657_));
 sky130_fd_sc_hd__a21oi_1 _11778_ (.A1(_05628_),
    .A2(_05634_),
    .B1(_05656_),
    .Y(_05658_));
 sky130_fd_sc_hd__or3b_1 _11779_ (.A(_05657_),
    .B(_05658_),
    .C_N(net174),
    .X(_05659_));
 sky130_fd_sc_hd__o21bai_1 _11780_ (.A1(_05651_),
    .A2(_05652_),
    .B1_N(net174),
    .Y(_05660_));
 sky130_fd_sc_hd__o21a_1 _11781_ (.A1(_05639_),
    .A2(_05641_),
    .B1(_05637_),
    .X(_05661_));
 sky130_fd_sc_hd__nand2_1 _11782_ (.A(net944),
    .B(_01534_),
    .Y(_05662_));
 sky130_fd_sc_hd__inv_2 _11783_ (.A(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__nor2_1 _11784_ (.A(net944),
    .B(_01534_),
    .Y(_05664_));
 sky130_fd_sc_hd__o21ai_1 _11785_ (.A1(_05663_),
    .A2(_05664_),
    .B1(_05661_),
    .Y(_05665_));
 sky130_fd_sc_hd__o31a_1 _11786_ (.A1(_05661_),
    .A2(_05663_),
    .A3(_05664_),
    .B1(net956),
    .X(_05666_));
 sky130_fd_sc_hd__a32o_1 _11787_ (.A1(_01208_),
    .A2(_05659_),
    .A3(_05660_),
    .B1(_05665_),
    .B2(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__o21ai_1 _11788_ (.A1(_05627_),
    .A2(_05645_),
    .B1(_05656_),
    .Y(_05668_));
 sky130_fd_sc_hd__o31a_1 _11789_ (.A1(_05627_),
    .A2(_05645_),
    .A3(_05656_),
    .B1(net952),
    .X(_05669_));
 sky130_fd_sc_hd__a22o_1 _11790_ (.A1(net836),
    .A2(_05667_),
    .B1(_05668_),
    .B2(_05669_),
    .X(_05670_));
 sky130_fd_sc_hd__mux2_1 _11791_ (.A0(net137),
    .A1(_05670_),
    .S(net204),
    .X(_05671_));
 sky130_fd_sc_hd__and2_1 _11792_ (.A(net1136),
    .B(_05671_),
    .X(_01135_));
 sky130_fd_sc_hd__or2_1 _11793_ (.A(\brancher.imm13_b[11] ),
    .B(\brancher.rPc_current_reg2[12] ),
    .X(_05672_));
 sky130_fd_sc_hd__nand2_1 _11794_ (.A(\brancher.imm13_b[11] ),
    .B(\brancher.rPc_current_reg2[12] ),
    .Y(_05673_));
 sky130_fd_sc_hd__nand2_1 _11795_ (.A(_05672_),
    .B(_05673_),
    .Y(_05674_));
 sky130_fd_sc_hd__a31o_1 _11796_ (.A1(_05628_),
    .A2(_05634_),
    .A3(_05655_),
    .B1(_05654_),
    .X(_05675_));
 sky130_fd_sc_hd__xnor2_1 _11797_ (.A(_05674_),
    .B(_05675_),
    .Y(_05676_));
 sky130_fd_sc_hd__xnor2_1 _11798_ (.A(net138),
    .B(_05651_),
    .Y(_05677_));
 sky130_fd_sc_hd__xnor2_1 _11799_ (.A(net944),
    .B(_01558_),
    .Y(_05678_));
 sky130_fd_sc_hd__o311a_1 _11800_ (.A1(_05615_),
    .A2(_05639_),
    .A3(_05640_),
    .B1(_05662_),
    .C1(_05637_),
    .X(_05679_));
 sky130_fd_sc_hd__o21ai_1 _11801_ (.A1(_05664_),
    .A2(_05679_),
    .B1(_05678_),
    .Y(_05680_));
 sky130_fd_sc_hd__or3_1 _11802_ (.A(_05664_),
    .B(_05678_),
    .C(_05679_),
    .X(_05681_));
 sky130_fd_sc_hd__xor2_1 _11803_ (.A(net918),
    .B(\brancher.rPc_current_reg2[12] ),
    .X(_05682_));
 sky130_fd_sc_hd__o211ai_1 _11804_ (.A1(_05630_),
    .A2(_05644_),
    .B1(_05655_),
    .C1(_05628_),
    .Y(_05683_));
 sky130_fd_sc_hd__nand2_1 _11805_ (.A(_05653_),
    .B(_05683_),
    .Y(_05684_));
 sky130_fd_sc_hd__xor2_1 _11806_ (.A(_05682_),
    .B(_05684_),
    .X(_05685_));
 sky130_fd_sc_hd__nand2_1 _11807_ (.A(net952),
    .B(_05685_),
    .Y(_05686_));
 sky130_fd_sc_hd__mux2_1 _11808_ (.A0(_05677_),
    .A1(_05676_),
    .S(net174),
    .X(_05687_));
 sky130_fd_sc_hd__a31o_1 _11809_ (.A1(net957),
    .A2(_05680_),
    .A3(_05681_),
    .B1(net952),
    .X(_05688_));
 sky130_fd_sc_hd__o21bai_1 _11810_ (.A1(net957),
    .A2(_05687_),
    .B1_N(_05688_),
    .Y(_05689_));
 sky130_fd_sc_hd__and3_1 _11811_ (.A(net628),
    .B(_05686_),
    .C(_05689_),
    .X(_05690_));
 sky130_fd_sc_hd__o21ai_1 _11812_ (.A1(net628),
    .A2(_05677_),
    .B1(net204),
    .Y(_05691_));
 sky130_fd_sc_hd__o221a_1 _11813_ (.A1(net138),
    .A2(net204),
    .B1(_05690_),
    .B2(_05691_),
    .C1(net1136),
    .X(_01136_));
 sky130_fd_sc_hd__and3_1 _11814_ (.A(net139),
    .B(net138),
    .C(_05651_),
    .X(_05692_));
 sky130_fd_sc_hd__a21oi_1 _11815_ (.A1(net138),
    .A2(_05651_),
    .B1(net139),
    .Y(_05693_));
 sky130_fd_sc_hd__nor2_1 _11816_ (.A(_05692_),
    .B(_05693_),
    .Y(_05694_));
 sky130_fd_sc_hd__o21ai_1 _11817_ (.A1(_05674_),
    .A2(_05675_),
    .B1(_05673_),
    .Y(_05695_));
 sky130_fd_sc_hd__or2_1 _11818_ (.A(net840),
    .B(\brancher.rPc_current_reg2[13] ),
    .X(_05696_));
 sky130_fd_sc_hd__nand2_1 _11819_ (.A(net840),
    .B(\brancher.rPc_current_reg2[13] ),
    .Y(_05697_));
 sky130_fd_sc_hd__nand2_1 _11820_ (.A(_05696_),
    .B(_05697_),
    .Y(_05698_));
 sky130_fd_sc_hd__xnor2_1 _11821_ (.A(_05695_),
    .B(_05698_),
    .Y(_05699_));
 sky130_fd_sc_hd__mux2_1 _11822_ (.A0(_05694_),
    .A1(_05699_),
    .S(net175),
    .X(_05700_));
 sky130_fd_sc_hd__xnor2_1 _11823_ (.A(net944),
    .B(_01580_),
    .Y(_05701_));
 sky130_fd_sc_hd__a21bo_1 _11824_ (.A1(net944),
    .A2(_01558_),
    .B1_N(_05681_),
    .X(_05702_));
 sky130_fd_sc_hd__xnor2_1 _11825_ (.A(_05701_),
    .B(_05702_),
    .Y(_05703_));
 sky130_fd_sc_hd__mux2_1 _11826_ (.A0(_05700_),
    .A1(_05703_),
    .S(net957),
    .X(_05704_));
 sky130_fd_sc_hd__a32o_1 _11827_ (.A1(_05653_),
    .A2(_05682_),
    .A3(_05683_),
    .B1(\brancher.rPc_current_reg2[12] ),
    .B2(net918),
    .X(_05705_));
 sky130_fd_sc_hd__or2_1 _11828_ (.A(net847),
    .B(\brancher.rPc_current_reg2[13] ),
    .X(_05706_));
 sky130_fd_sc_hd__nand2_1 _11829_ (.A(net847),
    .B(\brancher.rPc_current_reg2[13] ),
    .Y(_05707_));
 sky130_fd_sc_hd__a21oi_1 _11830_ (.A1(_05706_),
    .A2(_05707_),
    .B1(_05705_),
    .Y(_05708_));
 sky130_fd_sc_hd__a31o_1 _11831_ (.A1(_05705_),
    .A2(_05706_),
    .A3(_05707_),
    .B1(net836),
    .X(_05709_));
 sky130_fd_sc_hd__a2bb2o_1 _11832_ (.A1_N(_05708_),
    .A2_N(_05709_),
    .B1(net837),
    .B2(_05704_),
    .X(_05710_));
 sky130_fd_sc_hd__mux2_1 _11833_ (.A0(net139),
    .A1(_05710_),
    .S(net204),
    .X(_05711_));
 sky130_fd_sc_hd__and2_1 _11834_ (.A(net1136),
    .B(_05711_),
    .X(_01137_));
 sky130_fd_sc_hd__nand2_1 _11835_ (.A(net840),
    .B(\brancher.rPc_current_reg2[14] ),
    .Y(_05712_));
 sky130_fd_sc_hd__or2_1 _11836_ (.A(\brancher.imm13_b[12] ),
    .B(\brancher.rPc_current_reg2[14] ),
    .X(_05713_));
 sky130_fd_sc_hd__nand2_1 _11837_ (.A(_05712_),
    .B(_05713_),
    .Y(_05714_));
 sky130_fd_sc_hd__a21bo_1 _11838_ (.A1(_05695_),
    .A2(_05696_),
    .B1_N(_05697_),
    .X(_05715_));
 sky130_fd_sc_hd__nand2b_1 _11839_ (.A_N(_05714_),
    .B(_05715_),
    .Y(_05716_));
 sky130_fd_sc_hd__xor2_1 _11840_ (.A(_05714_),
    .B(_05715_),
    .X(_05717_));
 sky130_fd_sc_hd__and2_1 _11841_ (.A(net140),
    .B(_05692_),
    .X(_05718_));
 sky130_fd_sc_hd__nor2_1 _11842_ (.A(net140),
    .B(_05692_),
    .Y(_05719_));
 sky130_fd_sc_hd__or2_1 _11843_ (.A(_05718_),
    .B(_05719_),
    .X(_05720_));
 sky130_fd_sc_hd__inv_2 _11844_ (.A(_05720_),
    .Y(_05721_));
 sky130_fd_sc_hd__and2_1 _11845_ (.A(net944),
    .B(_01602_),
    .X(_05722_));
 sky130_fd_sc_hd__nor2_1 _11846_ (.A(net945),
    .B(_01602_),
    .Y(_05723_));
 sky130_fd_sc_hd__or2_1 _11847_ (.A(_05722_),
    .B(_05723_),
    .X(_05724_));
 sky130_fd_sc_hd__or2_1 _11848_ (.A(_05681_),
    .B(_05701_),
    .X(_05725_));
 sky130_fd_sc_hd__o21ai_1 _11849_ (.A1(_01558_),
    .A2(_01580_),
    .B1(net944),
    .Y(_05726_));
 sky130_fd_sc_hd__inv_2 _11850_ (.A(_05726_),
    .Y(_05727_));
 sky130_fd_sc_hd__and3_1 _11851_ (.A(_05724_),
    .B(_05725_),
    .C(_05726_),
    .X(_05728_));
 sky130_fd_sc_hd__a21oi_1 _11852_ (.A1(_05725_),
    .A2(_05726_),
    .B1(_05724_),
    .Y(_05729_));
 sky130_fd_sc_hd__xor2_1 _11853_ (.A(net845),
    .B(\brancher.rPc_current_reg2[14] ),
    .X(_05730_));
 sky130_fd_sc_hd__a21bo_1 _11854_ (.A1(_05705_),
    .A2(_05706_),
    .B1_N(_05707_),
    .X(_05731_));
 sky130_fd_sc_hd__and2_1 _11855_ (.A(_05730_),
    .B(_05731_),
    .X(_05732_));
 sky130_fd_sc_hd__nor2_1 _11856_ (.A(_05730_),
    .B(_05731_),
    .Y(_05733_));
 sky130_fd_sc_hd__o21ai_1 _11857_ (.A1(_05732_),
    .A2(_05733_),
    .B1(net953),
    .Y(_05734_));
 sky130_fd_sc_hd__mux2_1 _11858_ (.A0(_05720_),
    .A1(_05717_),
    .S(net175),
    .X(_05735_));
 sky130_fd_sc_hd__o31a_1 _11859_ (.A1(_01208_),
    .A2(_05728_),
    .A3(_05729_),
    .B1(net837),
    .X(_05736_));
 sky130_fd_sc_hd__o21ai_1 _11860_ (.A1(net956),
    .A2(_05735_),
    .B1(_05736_),
    .Y(_05737_));
 sky130_fd_sc_hd__and3_1 _11861_ (.A(_05456_),
    .B(_05734_),
    .C(_05737_),
    .X(_05738_));
 sky130_fd_sc_hd__a22o_1 _11862_ (.A1(net140),
    .A2(net201),
    .B1(_05463_),
    .B2(_05721_),
    .X(_05739_));
 sky130_fd_sc_hd__o21a_1 _11863_ (.A1(_05738_),
    .A2(_05739_),
    .B1(net1136),
    .X(_01138_));
 sky130_fd_sc_hd__xor2_1 _11864_ (.A(net141),
    .B(_05718_),
    .X(_05740_));
 sky130_fd_sc_hd__xnor2_1 _11865_ (.A(net840),
    .B(\brancher.rPc_current_reg2[15] ),
    .Y(_05741_));
 sky130_fd_sc_hd__nand2_1 _11866_ (.A(_05712_),
    .B(_05716_),
    .Y(_05742_));
 sky130_fd_sc_hd__xnor2_1 _11867_ (.A(_05741_),
    .B(_05742_),
    .Y(_05743_));
 sky130_fd_sc_hd__mux2_1 _11868_ (.A0(_05740_),
    .A1(_05743_),
    .S(net175),
    .X(_05744_));
 sky130_fd_sc_hd__xnor2_1 _11869_ (.A(net945),
    .B(_01624_),
    .Y(_05745_));
 sky130_fd_sc_hd__or2_1 _11870_ (.A(_05722_),
    .B(_05729_),
    .X(_05746_));
 sky130_fd_sc_hd__xnor2_1 _11871_ (.A(_05745_),
    .B(_05746_),
    .Y(_05747_));
 sky130_fd_sc_hd__mux2_1 _11872_ (.A0(_05744_),
    .A1(_05747_),
    .S(net957),
    .X(_05748_));
 sky130_fd_sc_hd__a21o_1 _11873_ (.A1(net845),
    .A2(\brancher.rPc_current_reg2[14] ),
    .B1(_05732_),
    .X(_05749_));
 sky130_fd_sc_hd__or2_1 _11874_ (.A(net943),
    .B(\brancher.rPc_current_reg2[15] ),
    .X(_05750_));
 sky130_fd_sc_hd__nand2_1 _11875_ (.A(net943),
    .B(\brancher.rPc_current_reg2[15] ),
    .Y(_05751_));
 sky130_fd_sc_hd__a21oi_1 _11876_ (.A1(_05750_),
    .A2(_05751_),
    .B1(_05749_),
    .Y(_05752_));
 sky130_fd_sc_hd__a31o_1 _11877_ (.A1(_05749_),
    .A2(_05750_),
    .A3(_05751_),
    .B1(net837),
    .X(_05753_));
 sky130_fd_sc_hd__a2bb2o_1 _11878_ (.A1_N(_05752_),
    .A2_N(_05753_),
    .B1(net837),
    .B2(_05748_),
    .X(_05754_));
 sky130_fd_sc_hd__mux2_1 _11879_ (.A0(net141),
    .A1(_05754_),
    .S(net204),
    .X(_05755_));
 sky130_fd_sc_hd__and2_1 _11880_ (.A(net1136),
    .B(_05755_),
    .X(_01139_));
 sky130_fd_sc_hd__xnor2_1 _11881_ (.A(net840),
    .B(\brancher.rPc_current_reg2[16] ),
    .Y(_05756_));
 sky130_fd_sc_hd__or2_1 _11882_ (.A(_05716_),
    .B(_05741_),
    .X(_05757_));
 sky130_fd_sc_hd__o21ai_1 _11883_ (.A1(\brancher.rPc_current_reg2[14] ),
    .A2(\brancher.rPc_current_reg2[15] ),
    .B1(net840),
    .Y(_05758_));
 sky130_fd_sc_hd__a21oi_1 _11884_ (.A1(_05757_),
    .A2(_05758_),
    .B1(_05756_),
    .Y(_05759_));
 sky130_fd_sc_hd__and3_1 _11885_ (.A(_05756_),
    .B(_05757_),
    .C(_05758_),
    .X(_05760_));
 sky130_fd_sc_hd__or2_1 _11886_ (.A(_05759_),
    .B(_05760_),
    .X(_05761_));
 sky130_fd_sc_hd__and3_1 _11887_ (.A(net142),
    .B(net141),
    .C(_05718_),
    .X(_05762_));
 sky130_fd_sc_hd__a21oi_1 _11888_ (.A1(net141),
    .A2(_05718_),
    .B1(net142),
    .Y(_05763_));
 sky130_fd_sc_hd__or2_1 _11889_ (.A(_05762_),
    .B(_05763_),
    .X(_05764_));
 sky130_fd_sc_hd__mux2_1 _11890_ (.A0(_05764_),
    .A1(_05761_),
    .S(net175),
    .X(_05765_));
 sky130_fd_sc_hd__nor2_1 _11891_ (.A(net956),
    .B(_05765_),
    .Y(_05766_));
 sky130_fd_sc_hd__or2_1 _11892_ (.A(_05724_),
    .B(_05745_),
    .X(_05767_));
 sky130_fd_sc_hd__a211oi_1 _11893_ (.A1(net945),
    .A2(_01624_),
    .B1(_05722_),
    .C1(_05727_),
    .Y(_05768_));
 sky130_fd_sc_hd__o31a_1 _11894_ (.A1(_05681_),
    .A2(_05701_),
    .A3(_05767_),
    .B1(_05768_),
    .X(_05769_));
 sky130_fd_sc_hd__nand2_1 _11895_ (.A(net945),
    .B(_01644_),
    .Y(_05770_));
 sky130_fd_sc_hd__or2_1 _11896_ (.A(net945),
    .B(_01644_),
    .X(_05771_));
 sky130_fd_sc_hd__nand2_1 _11897_ (.A(_05770_),
    .B(_05771_),
    .Y(_05772_));
 sky130_fd_sc_hd__or2_1 _11898_ (.A(_05769_),
    .B(_05772_),
    .X(_05773_));
 sky130_fd_sc_hd__nand2_1 _11899_ (.A(_05769_),
    .B(_05772_),
    .Y(_05774_));
 sky130_fd_sc_hd__a311o_1 _11900_ (.A1(net960),
    .A2(_05773_),
    .A3(_05774_),
    .B1(_05766_),
    .C1(net954),
    .X(_05775_));
 sky130_fd_sc_hd__nor2_1 _11901_ (.A(net1064),
    .B(\brancher.rPc_current_reg2[16] ),
    .Y(_05776_));
 sky130_fd_sc_hd__and2_1 _11902_ (.A(net1064),
    .B(\brancher.rPc_current_reg2[16] ),
    .X(_05777_));
 sky130_fd_sc_hd__nor2_1 _11903_ (.A(_05776_),
    .B(_05777_),
    .Y(_05778_));
 sky130_fd_sc_hd__a221o_1 _11904_ (.A1(net845),
    .A2(\brancher.rPc_current_reg2[14] ),
    .B1(\brancher.rPc_current_reg2[15] ),
    .B2(net943),
    .C1(_05732_),
    .X(_05779_));
 sky130_fd_sc_hd__and2_1 _11905_ (.A(_05750_),
    .B(_05779_),
    .X(_05780_));
 sky130_fd_sc_hd__xor2_1 _11906_ (.A(_05778_),
    .B(_05780_),
    .X(_05781_));
 sky130_fd_sc_hd__o211a_1 _11907_ (.A1(net837),
    .A2(_05781_),
    .B1(_05775_),
    .C1(_05456_),
    .X(_05782_));
 sky130_fd_sc_hd__nor2_1 _11908_ (.A(net628),
    .B(_05764_),
    .Y(_05783_));
 sky130_fd_sc_hd__mux2_1 _11909_ (.A0(net142),
    .A1(_05783_),
    .S(net204),
    .X(_05784_));
 sky130_fd_sc_hd__o21a_1 _11910_ (.A1(_05782_),
    .A2(_05784_),
    .B1(net1188),
    .X(_01140_));
 sky130_fd_sc_hd__xnor2_1 _11911_ (.A(net840),
    .B(\brancher.rPc_current_reg2[17] ),
    .Y(_05785_));
 sky130_fd_sc_hd__a21oi_1 _11912_ (.A1(net840),
    .A2(\brancher.rPc_current_reg2[16] ),
    .B1(_05759_),
    .Y(_05786_));
 sky130_fd_sc_hd__xnor2_1 _11913_ (.A(_05785_),
    .B(_05786_),
    .Y(_05787_));
 sky130_fd_sc_hd__and2_1 _11914_ (.A(net143),
    .B(_05762_),
    .X(_05788_));
 sky130_fd_sc_hd__nor2_1 _11915_ (.A(net143),
    .B(_05762_),
    .Y(_05789_));
 sky130_fd_sc_hd__or2_1 _11916_ (.A(_05788_),
    .B(_05789_),
    .X(_05790_));
 sky130_fd_sc_hd__mux2_1 _11917_ (.A0(_05790_),
    .A1(_05787_),
    .S(net175),
    .X(_05791_));
 sky130_fd_sc_hd__xnor2_1 _11918_ (.A(net812),
    .B(_01666_),
    .Y(_05792_));
 sky130_fd_sc_hd__and3_1 _11919_ (.A(_05770_),
    .B(_05773_),
    .C(_05792_),
    .X(_05793_));
 sky130_fd_sc_hd__a21oi_1 _11920_ (.A1(_05770_),
    .A2(_05773_),
    .B1(_05792_),
    .Y(_05794_));
 sky130_fd_sc_hd__or3_1 _11921_ (.A(_05447_),
    .B(_05793_),
    .C(_05794_),
    .X(_05795_));
 sky130_fd_sc_hd__a31oi_2 _11922_ (.A1(_05750_),
    .A2(_05778_),
    .A3(_05779_),
    .B1(_05777_),
    .Y(_05796_));
 sky130_fd_sc_hd__nor2_1 _11923_ (.A(net1030),
    .B(\brancher.rPc_current_reg2[17] ),
    .Y(_05797_));
 sky130_fd_sc_hd__and2_1 _11924_ (.A(net1030),
    .B(\brancher.rPc_current_reg2[17] ),
    .X(_05798_));
 sky130_fd_sc_hd__nor3_1 _11925_ (.A(_05796_),
    .B(_05797_),
    .C(_05798_),
    .Y(_05799_));
 sky130_fd_sc_hd__o21a_1 _11926_ (.A1(_05797_),
    .A2(_05798_),
    .B1(_05796_),
    .X(_05800_));
 sky130_fd_sc_hd__o311a_1 _11927_ (.A1(net838),
    .A2(_05799_),
    .A3(_05800_),
    .B1(net629),
    .C1(_05795_),
    .X(_05801_));
 sky130_fd_sc_hd__o21ai_1 _11928_ (.A1(_03218_),
    .A2(_05791_),
    .B1(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__a21oi_1 _11929_ (.A1(net630),
    .A2(_05790_),
    .B1(net200),
    .Y(_05803_));
 sky130_fd_sc_hd__a22o_1 _11930_ (.A1(net143),
    .A2(net200),
    .B1(_05802_),
    .B2(_05803_),
    .X(_05804_));
 sky130_fd_sc_hd__and2_1 _11931_ (.A(net1188),
    .B(_05804_),
    .X(_01141_));
 sky130_fd_sc_hd__and2_1 _11932_ (.A(net844),
    .B(\brancher.rPc_current_reg2[18] ),
    .X(_05805_));
 sky130_fd_sc_hd__nor2_1 _11933_ (.A(net844),
    .B(\brancher.rPc_current_reg2[18] ),
    .Y(_05806_));
 sky130_fd_sc_hd__or2_1 _11934_ (.A(_05805_),
    .B(_05806_),
    .X(_05807_));
 sky130_fd_sc_hd__or3_1 _11935_ (.A(_05756_),
    .B(_05757_),
    .C(_05785_),
    .X(_05808_));
 sky130_fd_sc_hd__o21ai_1 _11936_ (.A1(\brancher.rPc_current_reg2[16] ),
    .A2(\brancher.rPc_current_reg2[17] ),
    .B1(net840),
    .Y(_05809_));
 sky130_fd_sc_hd__and3_1 _11937_ (.A(_05758_),
    .B(_05808_),
    .C(_05809_),
    .X(_05810_));
 sky130_fd_sc_hd__xnor2_1 _11938_ (.A(_05807_),
    .B(_05810_),
    .Y(_05811_));
 sky130_fd_sc_hd__nand2_1 _11939_ (.A(net144),
    .B(_05788_),
    .Y(_05812_));
 sky130_fd_sc_hd__or2_1 _11940_ (.A(net144),
    .B(_05788_),
    .X(_05813_));
 sky130_fd_sc_hd__nand2_1 _11941_ (.A(_05812_),
    .B(_05813_),
    .Y(_05814_));
 sky130_fd_sc_hd__and2_1 _11942_ (.A(net945),
    .B(_01689_),
    .X(_05815_));
 sky130_fd_sc_hd__nor2_1 _11943_ (.A(net945),
    .B(_01689_),
    .Y(_05816_));
 sky130_fd_sc_hd__or2_1 _11944_ (.A(_05815_),
    .B(_05816_),
    .X(_05817_));
 sky130_fd_sc_hd__or2_1 _11945_ (.A(_05773_),
    .B(_05792_),
    .X(_05818_));
 sky130_fd_sc_hd__o21ai_1 _11946_ (.A1(net812),
    .A2(_01666_),
    .B1(_05770_),
    .Y(_05819_));
 sky130_fd_sc_hd__inv_2 _11947_ (.A(_05819_),
    .Y(_05820_));
 sky130_fd_sc_hd__and3_1 _11948_ (.A(_05817_),
    .B(_05818_),
    .C(_05820_),
    .X(_05821_));
 sky130_fd_sc_hd__a21oi_1 _11949_ (.A1(_05818_),
    .A2(_05820_),
    .B1(_05817_),
    .Y(_05822_));
 sky130_fd_sc_hd__or2_1 _11950_ (.A(net997),
    .B(\brancher.rPc_current_reg2[18] ),
    .X(_05823_));
 sky130_fd_sc_hd__nand2_1 _11951_ (.A(net997),
    .B(\brancher.rPc_current_reg2[18] ),
    .Y(_05824_));
 sky130_fd_sc_hd__nand2_1 _11952_ (.A(_05823_),
    .B(_05824_),
    .Y(_05825_));
 sky130_fd_sc_hd__o21ba_1 _11953_ (.A1(_05796_),
    .A2(_05797_),
    .B1_N(_05798_),
    .X(_05826_));
 sky130_fd_sc_hd__xnor2_1 _11954_ (.A(_05825_),
    .B(_05826_),
    .Y(_05827_));
 sky130_fd_sc_hd__nand2_1 _11955_ (.A(net954),
    .B(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__mux2_1 _11956_ (.A0(_05814_),
    .A1(_05811_),
    .S(net178),
    .X(_05829_));
 sky130_fd_sc_hd__or2_1 _11957_ (.A(net960),
    .B(_05829_),
    .X(_05830_));
 sky130_fd_sc_hd__o311ai_1 _11958_ (.A1(_01208_),
    .A2(_05821_),
    .A3(_05822_),
    .B1(_05830_),
    .C1(net838),
    .Y(_05831_));
 sky130_fd_sc_hd__nor2_1 _11959_ (.A(net629),
    .B(_05814_),
    .Y(_05832_));
 sky130_fd_sc_hd__a311o_1 _11960_ (.A1(net629),
    .A2(_05828_),
    .A3(_05831_),
    .B1(_05832_),
    .C1(net200),
    .X(_05833_));
 sky130_fd_sc_hd__o211a_1 _11961_ (.A1(net144),
    .A2(net203),
    .B1(_05833_),
    .C1(net1188),
    .X(_01142_));
 sky130_fd_sc_hd__nor2_1 _11962_ (.A(_01206_),
    .B(net203),
    .Y(_05834_));
 sky130_fd_sc_hd__xnor2_1 _11963_ (.A(net844),
    .B(\brancher.rPc_current_reg2[19] ),
    .Y(_05835_));
 sky130_fd_sc_hd__o21ba_1 _11964_ (.A1(_05806_),
    .A2(_05810_),
    .B1_N(_05805_),
    .X(_05836_));
 sky130_fd_sc_hd__xor2_1 _11965_ (.A(_05835_),
    .B(_05836_),
    .X(_05837_));
 sky130_fd_sc_hd__nor2_1 _11966_ (.A(_01206_),
    .B(_05812_),
    .Y(_05838_));
 sky130_fd_sc_hd__and2_1 _11967_ (.A(_01206_),
    .B(_05812_),
    .X(_05839_));
 sky130_fd_sc_hd__nor2_1 _11968_ (.A(_05838_),
    .B(_05839_),
    .Y(_05840_));
 sky130_fd_sc_hd__mux2_1 _11969_ (.A0(_05840_),
    .A1(_05837_),
    .S(net178),
    .X(_05841_));
 sky130_fd_sc_hd__o21a_1 _11970_ (.A1(_05825_),
    .A2(_05826_),
    .B1(_05824_),
    .X(_05842_));
 sky130_fd_sc_hd__and2_1 _11971_ (.A(net990),
    .B(\brancher.rPc_current_reg2[19] ),
    .X(_05843_));
 sky130_fd_sc_hd__nor2_1 _11972_ (.A(net990),
    .B(\brancher.rPc_current_reg2[19] ),
    .Y(_05844_));
 sky130_fd_sc_hd__or3_1 _11973_ (.A(_05842_),
    .B(_05843_),
    .C(_05844_),
    .X(_05845_));
 sky130_fd_sc_hd__o21ai_1 _11974_ (.A1(_05843_),
    .A2(_05844_),
    .B1(_05842_),
    .Y(_05846_));
 sky130_fd_sc_hd__xnor2_1 _11975_ (.A(net947),
    .B(_01709_),
    .Y(_05847_));
 sky130_fd_sc_hd__nor2_1 _11976_ (.A(_05815_),
    .B(_05822_),
    .Y(_05848_));
 sky130_fd_sc_hd__a21oi_1 _11977_ (.A1(_05847_),
    .A2(_05848_),
    .B1(_05447_),
    .Y(_05849_));
 sky130_fd_sc_hd__o21a_1 _11978_ (.A1(_05847_),
    .A2(_05848_),
    .B1(_05849_),
    .X(_05850_));
 sky130_fd_sc_hd__a311o_1 _11979_ (.A1(net954),
    .A2(_05845_),
    .A3(_05846_),
    .B1(_05850_),
    .C1(net630),
    .X(_05851_));
 sky130_fd_sc_hd__a21o_1 _11980_ (.A1(_03217_),
    .A2(_05841_),
    .B1(_05851_),
    .X(_05852_));
 sky130_fd_sc_hd__o211a_1 _11981_ (.A1(net629),
    .A2(_05840_),
    .B1(_05852_),
    .C1(net203),
    .X(_05853_));
 sky130_fd_sc_hd__o21a_1 _11982_ (.A1(_05834_),
    .A2(_05853_),
    .B1(net1188),
    .X(_01143_));
 sky130_fd_sc_hd__nand2_1 _11983_ (.A(net844),
    .B(\brancher.rPc_current_reg2[20] ),
    .Y(_05854_));
 sky130_fd_sc_hd__or2_1 _11984_ (.A(net844),
    .B(\brancher.rPc_current_reg2[20] ),
    .X(_05855_));
 sky130_fd_sc_hd__nand2_1 _11985_ (.A(_05854_),
    .B(_05855_),
    .Y(_05856_));
 sky130_fd_sc_hd__or3_1 _11986_ (.A(_05807_),
    .B(_05810_),
    .C(_05835_),
    .X(_05857_));
 sky130_fd_sc_hd__o21ai_1 _11987_ (.A1(\brancher.rPc_current_reg2[18] ),
    .A2(\brancher.rPc_current_reg2[19] ),
    .B1(net844),
    .Y(_05858_));
 sky130_fd_sc_hd__nand2_1 _11988_ (.A(_05857_),
    .B(_05858_),
    .Y(_05859_));
 sky130_fd_sc_hd__xnor2_1 _11989_ (.A(_05856_),
    .B(_05859_),
    .Y(_05860_));
 sky130_fd_sc_hd__and2_1 _11990_ (.A(net147),
    .B(_05838_),
    .X(_05861_));
 sky130_fd_sc_hd__nor2_1 _11991_ (.A(net147),
    .B(_05838_),
    .Y(_05862_));
 sky130_fd_sc_hd__nor2_1 _11992_ (.A(_05861_),
    .B(_05862_),
    .Y(_05863_));
 sky130_fd_sc_hd__mux2_1 _11993_ (.A0(_05863_),
    .A1(_05860_),
    .S(net178),
    .X(_05864_));
 sky130_fd_sc_hd__nor2_1 _11994_ (.A(net812),
    .B(_01732_),
    .Y(_05865_));
 sky130_fd_sc_hd__inv_2 _11995_ (.A(_05865_),
    .Y(_05866_));
 sky130_fd_sc_hd__nand2_1 _11996_ (.A(net812),
    .B(_01732_),
    .Y(_05867_));
 sky130_fd_sc_hd__nand2_1 _11997_ (.A(_05866_),
    .B(_05867_),
    .Y(_05868_));
 sky130_fd_sc_hd__or2_1 _11998_ (.A(_05817_),
    .B(_05847_),
    .X(_05869_));
 sky130_fd_sc_hd__nor4_1 _11999_ (.A(_05769_),
    .B(_05772_),
    .C(_05792_),
    .D(_05869_),
    .Y(_05870_));
 sky130_fd_sc_hd__a211oi_1 _12000_ (.A1(net947),
    .A2(_01709_),
    .B1(_05815_),
    .C1(_05819_),
    .Y(_05871_));
 sky130_fd_sc_hd__and2b_1 _12001_ (.A_N(net180),
    .B(_05871_),
    .X(_05872_));
 sky130_fd_sc_hd__or2_1 _12002_ (.A(_05868_),
    .B(_05872_),
    .X(_05873_));
 sky130_fd_sc_hd__nand2_1 _12003_ (.A(_05868_),
    .B(_05872_),
    .Y(_05874_));
 sky130_fd_sc_hd__a31o_1 _12004_ (.A1(net960),
    .A2(_05873_),
    .A3(_05874_),
    .B1(net954),
    .X(_05875_));
 sky130_fd_sc_hd__a21o_1 _12005_ (.A1(_01208_),
    .A2(_05864_),
    .B1(_05875_),
    .X(_05876_));
 sky130_fd_sc_hd__or2_1 _12006_ (.A(net1069),
    .B(\brancher.rPc_current_reg2[20] ),
    .X(_05877_));
 sky130_fd_sc_hd__nand2_1 _12007_ (.A(net1069),
    .B(\brancher.rPc_current_reg2[20] ),
    .Y(_05878_));
 sky130_fd_sc_hd__nand2_1 _12008_ (.A(_05877_),
    .B(_05878_),
    .Y(_05879_));
 sky130_fd_sc_hd__nor2_1 _12009_ (.A(_05842_),
    .B(_05844_),
    .Y(_05880_));
 sky130_fd_sc_hd__nor2_1 _12010_ (.A(_05843_),
    .B(_05880_),
    .Y(_05881_));
 sky130_fd_sc_hd__xnor2_1 _12011_ (.A(_05879_),
    .B(_05881_),
    .Y(_05882_));
 sky130_fd_sc_hd__nand2_1 _12012_ (.A(net954),
    .B(_05882_),
    .Y(_05883_));
 sky130_fd_sc_hd__and3_1 _12013_ (.A(_05456_),
    .B(_05876_),
    .C(_05883_),
    .X(_05884_));
 sky130_fd_sc_hd__a22o_1 _12014_ (.A1(net147),
    .A2(net200),
    .B1(_05463_),
    .B2(_05863_),
    .X(_05885_));
 sky130_fd_sc_hd__o21a_1 _12015_ (.A1(_05884_),
    .A2(_05885_),
    .B1(net1188),
    .X(_01144_));
 sky130_fd_sc_hd__nand2_1 _12016_ (.A(net148),
    .B(net200),
    .Y(_05886_));
 sky130_fd_sc_hd__nand2_1 _12017_ (.A(net844),
    .B(\brancher.rPc_current_reg2[21] ),
    .Y(_05887_));
 sky130_fd_sc_hd__or2_1 _12018_ (.A(net844),
    .B(\brancher.rPc_current_reg2[21] ),
    .X(_05888_));
 sky130_fd_sc_hd__nand2_1 _12019_ (.A(_05887_),
    .B(_05888_),
    .Y(_05889_));
 sky130_fd_sc_hd__a21bo_1 _12020_ (.A1(_05855_),
    .A2(_05859_),
    .B1_N(_05854_),
    .X(_05890_));
 sky130_fd_sc_hd__xor2_1 _12021_ (.A(_05889_),
    .B(_05890_),
    .X(_05891_));
 sky130_fd_sc_hd__xnor2_1 _12022_ (.A(net148),
    .B(_05861_),
    .Y(_05892_));
 sky130_fd_sc_hd__mux2_1 _12023_ (.A0(_05892_),
    .A1(_05891_),
    .S(net178),
    .X(_05893_));
 sky130_fd_sc_hd__nand2_1 _12024_ (.A(net947),
    .B(_01754_),
    .Y(_05894_));
 sky130_fd_sc_hd__and2_1 _12025_ (.A(_05866_),
    .B(_05873_),
    .X(_05895_));
 sky130_fd_sc_hd__nor2_1 _12026_ (.A(net947),
    .B(_01754_),
    .Y(_05896_));
 sky130_fd_sc_hd__inv_2 _12027_ (.A(_05896_),
    .Y(_05897_));
 sky130_fd_sc_hd__nand2_1 _12028_ (.A(_05894_),
    .B(_05897_),
    .Y(_05898_));
 sky130_fd_sc_hd__xnor2_1 _12029_ (.A(_05895_),
    .B(_05898_),
    .Y(_05899_));
 sky130_fd_sc_hd__o21a_1 _12030_ (.A1(_05879_),
    .A2(_05881_),
    .B1(_05878_),
    .X(_05900_));
 sky130_fd_sc_hd__and2_1 _12031_ (.A(_05889_),
    .B(_05900_),
    .X(_05901_));
 sky130_fd_sc_hd__nor2_1 _12032_ (.A(_05889_),
    .B(_05900_),
    .Y(_05902_));
 sky130_fd_sc_hd__o32a_1 _12033_ (.A1(net838),
    .A2(_05901_),
    .A3(_05902_),
    .B1(_05447_),
    .B2(_05899_),
    .X(_05903_));
 sky130_fd_sc_hd__o211a_1 _12034_ (.A1(_03218_),
    .A2(_05893_),
    .B1(_05903_),
    .C1(net628),
    .X(_05904_));
 sky130_fd_sc_hd__a211o_1 _12035_ (.A1(net630),
    .A2(_05892_),
    .B1(_05904_),
    .C1(net200),
    .X(_05905_));
 sky130_fd_sc_hd__a21boi_1 _12036_ (.A1(_05886_),
    .A2(_05905_),
    .B1_N(net1188),
    .Y(_01145_));
 sky130_fd_sc_hd__and2_1 _12037_ (.A(net149),
    .B(net200),
    .X(_05906_));
 sky130_fd_sc_hd__and3_1 _12038_ (.A(net149),
    .B(net148),
    .C(_05861_),
    .X(_05907_));
 sky130_fd_sc_hd__a21oi_1 _12039_ (.A1(net148),
    .A2(_05861_),
    .B1(net149),
    .Y(_05908_));
 sky130_fd_sc_hd__nor2_1 _12040_ (.A(_05907_),
    .B(_05908_),
    .Y(_05909_));
 sky130_fd_sc_hd__or2_1 _12041_ (.A(net841),
    .B(\brancher.rPc_current_reg2[22] ),
    .X(_05910_));
 sky130_fd_sc_hd__nand2_1 _12042_ (.A(net841),
    .B(\brancher.rPc_current_reg2[22] ),
    .Y(_05911_));
 sky130_fd_sc_hd__and2_1 _12043_ (.A(_05910_),
    .B(_05911_),
    .X(_05912_));
 sky130_fd_sc_hd__nand2_1 _12044_ (.A(_05910_),
    .B(_05911_),
    .Y(_05913_));
 sky130_fd_sc_hd__and3_1 _12045_ (.A(_05854_),
    .B(_05858_),
    .C(_05887_),
    .X(_05914_));
 sky130_fd_sc_hd__o31a_1 _12046_ (.A1(_05856_),
    .A2(_05857_),
    .A3(_05889_),
    .B1(_05914_),
    .X(_05915_));
 sky130_fd_sc_hd__or2_1 _12047_ (.A(_05913_),
    .B(_05915_),
    .X(_05916_));
 sky130_fd_sc_hd__nand2_1 _12048_ (.A(_05913_),
    .B(_05915_),
    .Y(_05917_));
 sky130_fd_sc_hd__nand2_1 _12049_ (.A(net947),
    .B(_01776_),
    .Y(_05918_));
 sky130_fd_sc_hd__or2_1 _12050_ (.A(net947),
    .B(_01776_),
    .X(_05919_));
 sky130_fd_sc_hd__nand2_1 _12051_ (.A(_05918_),
    .B(_05919_),
    .Y(_05920_));
 sky130_fd_sc_hd__a31o_1 _12052_ (.A1(_05866_),
    .A2(_05873_),
    .A3(_05894_),
    .B1(_05896_),
    .X(_05921_));
 sky130_fd_sc_hd__and2b_1 _12053_ (.A_N(net177),
    .B(_05909_),
    .X(_05922_));
 sky130_fd_sc_hd__a311o_1 _12054_ (.A1(net177),
    .A2(_05916_),
    .A3(_05917_),
    .B1(_05922_),
    .C1(net958),
    .X(_05923_));
 sky130_fd_sc_hd__xnor2_1 _12055_ (.A(_05920_),
    .B(_05921_),
    .Y(_05924_));
 sky130_fd_sc_hd__nand2_1 _12056_ (.A(net958),
    .B(_05924_),
    .Y(_05925_));
 sky130_fd_sc_hd__a21boi_1 _12057_ (.A1(_05887_),
    .A2(_05900_),
    .B1_N(_05888_),
    .Y(_05926_));
 sky130_fd_sc_hd__or2_1 _12058_ (.A(_05912_),
    .B(_05926_),
    .X(_05927_));
 sky130_fd_sc_hd__nand2_1 _12059_ (.A(_05912_),
    .B(_05926_),
    .Y(_05928_));
 sky130_fd_sc_hd__a31o_1 _12060_ (.A1(net954),
    .A2(_05927_),
    .A3(_05928_),
    .B1(net630),
    .X(_05929_));
 sky130_fd_sc_hd__a31o_1 _12061_ (.A1(net839),
    .A2(_05923_),
    .A3(_05925_),
    .B1(_05929_),
    .X(_05930_));
 sky130_fd_sc_hd__o211a_1 _12062_ (.A1(net628),
    .A2(_05909_),
    .B1(_05930_),
    .C1(net202),
    .X(_05931_));
 sky130_fd_sc_hd__o21a_1 _12063_ (.A1(_05906_),
    .A2(_05931_),
    .B1(net1188),
    .X(_01146_));
 sky130_fd_sc_hd__xnor2_2 _12064_ (.A(net841),
    .B(\brancher.rPc_current_reg2[23] ),
    .Y(_05932_));
 sky130_fd_sc_hd__o21ai_1 _12065_ (.A1(_05913_),
    .A2(_05915_),
    .B1(_05911_),
    .Y(_05933_));
 sky130_fd_sc_hd__xnor2_1 _12066_ (.A(_05932_),
    .B(_05933_),
    .Y(_05934_));
 sky130_fd_sc_hd__and2_1 _12067_ (.A(net150),
    .B(_05907_),
    .X(_05935_));
 sky130_fd_sc_hd__nor2_1 _12068_ (.A(net150),
    .B(_05907_),
    .Y(_05936_));
 sky130_fd_sc_hd__nor2_1 _12069_ (.A(_05935_),
    .B(_05936_),
    .Y(_05937_));
 sky130_fd_sc_hd__a21oi_1 _12070_ (.A1(_05911_),
    .A2(_05928_),
    .B1(_05932_),
    .Y(_05938_));
 sky130_fd_sc_hd__a31o_1 _12071_ (.A1(_05911_),
    .A2(_05928_),
    .A3(_05932_),
    .B1(net838),
    .X(_05939_));
 sky130_fd_sc_hd__nor2_1 _12072_ (.A(_05938_),
    .B(_05939_),
    .Y(_05940_));
 sky130_fd_sc_hd__xnor2_1 _12073_ (.A(net812),
    .B(_01798_),
    .Y(_05941_));
 sky130_fd_sc_hd__o21ai_1 _12074_ (.A1(_05920_),
    .A2(_05921_),
    .B1(_05918_),
    .Y(_05942_));
 sky130_fd_sc_hd__mux2_1 _12075_ (.A0(_05937_),
    .A1(_05934_),
    .S(net177),
    .X(_05943_));
 sky130_fd_sc_hd__xnor2_1 _12076_ (.A(_05941_),
    .B(_05942_),
    .Y(_05944_));
 sky130_fd_sc_hd__mux2_1 _12077_ (.A0(_05943_),
    .A1(_05944_),
    .S(net958),
    .X(_05945_));
 sky130_fd_sc_hd__a211o_1 _12078_ (.A1(net838),
    .A2(_05945_),
    .B1(_05940_),
    .C1(net630),
    .X(_05946_));
 sky130_fd_sc_hd__o21a_1 _12079_ (.A1(net628),
    .A2(_05937_),
    .B1(net202),
    .X(_05947_));
 sky130_fd_sc_hd__a22o_1 _12080_ (.A1(net150),
    .A2(net200),
    .B1(_05946_),
    .B2(_05947_),
    .X(_05948_));
 sky130_fd_sc_hd__and2_1 _12081_ (.A(net1188),
    .B(_05948_),
    .X(_01147_));
 sky130_fd_sc_hd__nand2_1 _12082_ (.A(net843),
    .B(\brancher.rPc_current_reg2[24] ),
    .Y(_05949_));
 sky130_fd_sc_hd__or2_1 _12083_ (.A(net843),
    .B(\brancher.rPc_current_reg2[24] ),
    .X(_05950_));
 sky130_fd_sc_hd__nand2_2 _12084_ (.A(_05949_),
    .B(_05950_),
    .Y(_05951_));
 sky130_fd_sc_hd__o21ai_1 _12085_ (.A1(\brancher.rPc_current_reg2[22] ),
    .A2(\brancher.rPc_current_reg2[23] ),
    .B1(net841),
    .Y(_05952_));
 sky130_fd_sc_hd__o31a_1 _12086_ (.A1(_05913_),
    .A2(_05915_),
    .A3(_05932_),
    .B1(_05952_),
    .X(_05953_));
 sky130_fd_sc_hd__xnor2_1 _12087_ (.A(_05951_),
    .B(_05953_),
    .Y(_05954_));
 sky130_fd_sc_hd__nand2_1 _12088_ (.A(net151),
    .B(_05935_),
    .Y(_05955_));
 sky130_fd_sc_hd__or2_1 _12089_ (.A(net151),
    .B(_05935_),
    .X(_05956_));
 sky130_fd_sc_hd__nand2_1 _12090_ (.A(_05955_),
    .B(_05956_),
    .Y(_05957_));
 sky130_fd_sc_hd__mux2_1 _12091_ (.A0(_05957_),
    .A1(_05954_),
    .S(net177),
    .X(_05958_));
 sky130_fd_sc_hd__and2_1 _12092_ (.A(net946),
    .B(_01820_),
    .X(_05959_));
 sky130_fd_sc_hd__nor2_1 _12093_ (.A(net946),
    .B(_01820_),
    .Y(_05960_));
 sky130_fd_sc_hd__or2_1 _12094_ (.A(_05959_),
    .B(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__nor4_1 _12095_ (.A(_05868_),
    .B(_05898_),
    .C(_05920_),
    .D(_05941_),
    .Y(_05962_));
 sky130_fd_sc_hd__nand2_1 _12096_ (.A(net180),
    .B(_05962_),
    .Y(_05963_));
 sky130_fd_sc_hd__o211a_1 _12097_ (.A1(net812),
    .A2(_01798_),
    .B1(_05866_),
    .C1(_05894_),
    .X(_05964_));
 sky130_fd_sc_hd__and3_1 _12098_ (.A(_05871_),
    .B(_05918_),
    .C(_05964_),
    .X(_05965_));
 sky130_fd_sc_hd__a21o_1 _12099_ (.A1(_05963_),
    .A2(_05965_),
    .B1(_05961_),
    .X(_05966_));
 sky130_fd_sc_hd__nand2_1 _12100_ (.A(net959),
    .B(_05966_),
    .Y(_05967_));
 sky130_fd_sc_hd__a31o_1 _12101_ (.A1(_05961_),
    .A2(_05963_),
    .A3(_05965_),
    .B1(_05967_),
    .X(_05968_));
 sky130_fd_sc_hd__o211a_1 _12102_ (.A1(net958),
    .A2(_05958_),
    .B1(_05968_),
    .C1(net838),
    .X(_05969_));
 sky130_fd_sc_hd__o21a_1 _12103_ (.A1(_05928_),
    .A2(_05932_),
    .B1(_05952_),
    .X(_05970_));
 sky130_fd_sc_hd__xnor2_1 _12104_ (.A(_05951_),
    .B(_05970_),
    .Y(_05971_));
 sky130_fd_sc_hd__a211o_1 _12105_ (.A1(net955),
    .A2(_05971_),
    .B1(_05969_),
    .C1(net630),
    .X(_05972_));
 sky130_fd_sc_hd__o211ai_1 _12106_ (.A1(net628),
    .A2(_05957_),
    .B1(_05972_),
    .C1(net202),
    .Y(_05973_));
 sky130_fd_sc_hd__o211a_1 _12107_ (.A1(net151),
    .A2(net202),
    .B1(_05973_),
    .C1(net1190),
    .X(_01148_));
 sky130_fd_sc_hd__or2_1 _12108_ (.A(net841),
    .B(\brancher.rPc_current_reg2[25] ),
    .X(_05974_));
 sky130_fd_sc_hd__nand2_1 _12109_ (.A(net841),
    .B(\brancher.rPc_current_reg2[25] ),
    .Y(_05975_));
 sky130_fd_sc_hd__and2_1 _12110_ (.A(_05974_),
    .B(_05975_),
    .X(_05976_));
 sky130_fd_sc_hd__o21a_1 _12111_ (.A1(_05951_),
    .A2(_05953_),
    .B1(_05949_),
    .X(_05977_));
 sky130_fd_sc_hd__xnor2_1 _12112_ (.A(_05976_),
    .B(_05977_),
    .Y(_05978_));
 sky130_fd_sc_hd__xnor2_1 _12113_ (.A(net152),
    .B(_05955_),
    .Y(_05979_));
 sky130_fd_sc_hd__o21ai_1 _12114_ (.A1(_05951_),
    .A2(_05970_),
    .B1(_05949_),
    .Y(_05980_));
 sky130_fd_sc_hd__nand2_1 _12115_ (.A(_05976_),
    .B(_05980_),
    .Y(_05981_));
 sky130_fd_sc_hd__o21a_1 _12116_ (.A1(_05976_),
    .A2(_05980_),
    .B1(net955),
    .X(_05982_));
 sky130_fd_sc_hd__xnor2_1 _12117_ (.A(net812),
    .B(_01842_),
    .Y(_05983_));
 sky130_fd_sc_hd__and2b_1 _12118_ (.A_N(_05959_),
    .B(_05966_),
    .X(_05984_));
 sky130_fd_sc_hd__mux2_1 _12119_ (.A0(_05979_),
    .A1(_05978_),
    .S(net178),
    .X(_05985_));
 sky130_fd_sc_hd__xnor2_1 _12120_ (.A(_05983_),
    .B(_05984_),
    .Y(_05986_));
 sky130_fd_sc_hd__nand2_1 _12121_ (.A(net958),
    .B(_05986_),
    .Y(_05987_));
 sky130_fd_sc_hd__o211a_1 _12122_ (.A1(net958),
    .A2(_05985_),
    .B1(_05987_),
    .C1(net838),
    .X(_05988_));
 sky130_fd_sc_hd__a211o_1 _12123_ (.A1(_05981_),
    .A2(_05982_),
    .B1(_05988_),
    .C1(net630),
    .X(_05989_));
 sky130_fd_sc_hd__o21a_1 _12124_ (.A1(net629),
    .A2(_05979_),
    .B1(net202),
    .X(_05990_));
 sky130_fd_sc_hd__a22o_1 _12125_ (.A1(net152),
    .A2(net200),
    .B1(_05989_),
    .B2(_05990_),
    .X(_05991_));
 sky130_fd_sc_hd__and2_1 _12126_ (.A(net1190),
    .B(_05991_),
    .X(_01149_));
 sky130_fd_sc_hd__and2_1 _12127_ (.A(net841),
    .B(\brancher.rPc_current_reg2[26] ),
    .X(_05992_));
 sky130_fd_sc_hd__nor2_1 _12128_ (.A(net841),
    .B(\brancher.rPc_current_reg2[26] ),
    .Y(_05993_));
 sky130_fd_sc_hd__or2_1 _12129_ (.A(_05992_),
    .B(_05993_),
    .X(_05994_));
 sky130_fd_sc_hd__nor4b_1 _12130_ (.A(_05913_),
    .B(_05932_),
    .C(_05951_),
    .D_N(_05976_),
    .Y(_05995_));
 sky130_fd_sc_hd__or4b_1 _12131_ (.A(_05856_),
    .B(_05857_),
    .C(_05889_),
    .D_N(net432),
    .X(_05996_));
 sky130_fd_sc_hd__and3_1 _12132_ (.A(_05949_),
    .B(_05952_),
    .C(_05975_),
    .X(_05997_));
 sky130_fd_sc_hd__and3_1 _12133_ (.A(_05914_),
    .B(_05996_),
    .C(_05997_),
    .X(_05998_));
 sky130_fd_sc_hd__a31oi_2 _12134_ (.A1(_05914_),
    .A2(_05996_),
    .A3(_05997_),
    .B1(_05994_),
    .Y(_05999_));
 sky130_fd_sc_hd__and4_1 _12135_ (.A(net153),
    .B(net152),
    .C(net151),
    .D(_05935_),
    .X(_06000_));
 sky130_fd_sc_hd__a31o_1 _12136_ (.A1(net152),
    .A2(net151),
    .A3(_05935_),
    .B1(net153),
    .X(_06001_));
 sky130_fd_sc_hd__nand2b_1 _12137_ (.A_N(_06000_),
    .B(_06001_),
    .Y(_06002_));
 sky130_fd_sc_hd__xnor2_1 _12138_ (.A(net946),
    .B(_01863_),
    .Y(_06003_));
 sky130_fd_sc_hd__or2_1 _12139_ (.A(_05966_),
    .B(_05983_),
    .X(_06004_));
 sky130_fd_sc_hd__o21ba_1 _12140_ (.A1(net812),
    .A2(_01842_),
    .B1_N(_05959_),
    .X(_06005_));
 sky130_fd_sc_hd__a21oi_1 _12141_ (.A1(_06004_),
    .A2(_06005_),
    .B1(_06003_),
    .Y(_06006_));
 sky130_fd_sc_hd__and3_1 _12142_ (.A(_06003_),
    .B(_06004_),
    .C(_06005_),
    .X(_06007_));
 sky130_fd_sc_hd__a21bo_1 _12143_ (.A1(_05994_),
    .A2(_05998_),
    .B1_N(net177),
    .X(_06008_));
 sky130_fd_sc_hd__o221ai_1 _12144_ (.A1(net177),
    .A2(_06002_),
    .B1(_06008_),
    .B2(_05999_),
    .C1(_01208_),
    .Y(_06009_));
 sky130_fd_sc_hd__o21ai_1 _12145_ (.A1(_06006_),
    .A2(_06007_),
    .B1(net958),
    .Y(_06010_));
 sky130_fd_sc_hd__a21boi_1 _12146_ (.A1(_05926_),
    .A2(_05995_),
    .B1_N(_05997_),
    .Y(_06011_));
 sky130_fd_sc_hd__nand2_1 _12147_ (.A(_05994_),
    .B(_06011_),
    .Y(_06012_));
 sky130_fd_sc_hd__or2_1 _12148_ (.A(_05994_),
    .B(_06011_),
    .X(_06013_));
 sky130_fd_sc_hd__a31o_1 _12149_ (.A1(net955),
    .A2(_06012_),
    .A3(_06013_),
    .B1(net630),
    .X(_06014_));
 sky130_fd_sc_hd__a31o_1 _12150_ (.A1(net838),
    .A2(_06009_),
    .A3(_06010_),
    .B1(_06014_),
    .X(_06015_));
 sky130_fd_sc_hd__a21oi_1 _12151_ (.A1(_05454_),
    .A2(_06002_),
    .B1(net200),
    .Y(_06016_));
 sky130_fd_sc_hd__a22o_1 _12152_ (.A1(net153),
    .A2(_05453_),
    .B1(_06015_),
    .B2(_06016_),
    .X(_06017_));
 sky130_fd_sc_hd__and2_1 _12153_ (.A(net1190),
    .B(_06017_),
    .X(_01150_));
 sky130_fd_sc_hd__xor2_2 _12154_ (.A(net841),
    .B(\brancher.rPc_current_reg2[27] ),
    .X(_06018_));
 sky130_fd_sc_hd__or3_1 _12155_ (.A(_05992_),
    .B(_05999_),
    .C(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__o21ai_1 _12156_ (.A1(_05992_),
    .A2(_05999_),
    .B1(_06018_),
    .Y(_06020_));
 sky130_fd_sc_hd__xnor2_1 _12157_ (.A(net154),
    .B(_06000_),
    .Y(_06021_));
 sky130_fd_sc_hd__nor2_1 _12158_ (.A(net177),
    .B(_06021_),
    .Y(_06022_));
 sky130_fd_sc_hd__a311o_1 _12159_ (.A1(net177),
    .A2(_06019_),
    .A3(_06020_),
    .B1(_06022_),
    .C1(net958),
    .X(_06023_));
 sky130_fd_sc_hd__xnor2_1 _12160_ (.A(net946),
    .B(_01884_),
    .Y(_06024_));
 sky130_fd_sc_hd__a21oi_1 _12161_ (.A1(net946),
    .A2(_01863_),
    .B1(_06006_),
    .Y(_06025_));
 sky130_fd_sc_hd__xnor2_1 _12162_ (.A(_06024_),
    .B(_06025_),
    .Y(_06026_));
 sky130_fd_sc_hd__a21oi_1 _12163_ (.A1(net958),
    .A2(_06026_),
    .B1(net955),
    .Y(_06027_));
 sky130_fd_sc_hd__nand2b_1 _12164_ (.A_N(_05992_),
    .B(_06013_),
    .Y(_06028_));
 sky130_fd_sc_hd__xor2_1 _12165_ (.A(_06018_),
    .B(_06028_),
    .X(_06029_));
 sky130_fd_sc_hd__a22o_1 _12166_ (.A1(_06023_),
    .A2(_06027_),
    .B1(_06029_),
    .B2(net954),
    .X(_06030_));
 sky130_fd_sc_hd__mux2_1 _12167_ (.A0(net154),
    .A1(_06030_),
    .S(net202),
    .X(_06031_));
 sky130_fd_sc_hd__and2_1 _12168_ (.A(net1190),
    .B(_06031_),
    .X(_01151_));
 sky130_fd_sc_hd__and3_1 _12169_ (.A(net155),
    .B(net154),
    .C(_06000_),
    .X(_06032_));
 sky130_fd_sc_hd__a21oi_1 _12170_ (.A1(net154),
    .A2(_06000_),
    .B1(net155),
    .Y(_06033_));
 sky130_fd_sc_hd__nand2_1 _12171_ (.A(net842),
    .B(\brancher.rPc_current_reg2[28] ),
    .Y(_06034_));
 sky130_fd_sc_hd__or2_1 _12172_ (.A(net842),
    .B(\brancher.rPc_current_reg2[28] ),
    .X(_06035_));
 sky130_fd_sc_hd__nand2_1 _12173_ (.A(_06034_),
    .B(_06035_),
    .Y(_06036_));
 sky130_fd_sc_hd__o21ai_1 _12174_ (.A1(\brancher.rPc_current_reg2[26] ),
    .A2(\brancher.rPc_current_reg2[27] ),
    .B1(net841),
    .Y(_06037_));
 sky130_fd_sc_hd__nand2_1 _12175_ (.A(_05999_),
    .B(_06018_),
    .Y(_06038_));
 sky130_fd_sc_hd__and2_1 _12176_ (.A(_06037_),
    .B(_06038_),
    .X(_06039_));
 sky130_fd_sc_hd__xnor2_1 _12177_ (.A(_06036_),
    .B(_06039_),
    .Y(_06040_));
 sky130_fd_sc_hd__and2_1 _12178_ (.A(net177),
    .B(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__o21ba_1 _12179_ (.A1(_06032_),
    .A2(_06033_),
    .B1_N(net177),
    .X(_06042_));
 sky130_fd_sc_hd__or2_1 _12180_ (.A(_01219_),
    .B(_01906_),
    .X(_06043_));
 sky130_fd_sc_hd__nand2_1 _12181_ (.A(_01219_),
    .B(_01906_),
    .Y(_06044_));
 sky130_fd_sc_hd__nand2_1 _12182_ (.A(_06043_),
    .B(_06044_),
    .Y(_06045_));
 sky130_fd_sc_hd__or2_1 _12183_ (.A(_06003_),
    .B(_06024_),
    .X(_06046_));
 sky130_fd_sc_hd__a2111o_1 _12184_ (.A1(_05963_),
    .A2(_05965_),
    .B1(_05983_),
    .C1(_06046_),
    .D1(_05961_),
    .X(_06047_));
 sky130_fd_sc_hd__o21ai_1 _12185_ (.A1(_01863_),
    .A2(_01884_),
    .B1(net946),
    .Y(_06048_));
 sky130_fd_sc_hd__and4_1 _12186_ (.A(_06005_),
    .B(_06045_),
    .C(_06047_),
    .D(_06048_),
    .X(_06049_));
 sky130_fd_sc_hd__a31o_1 _12187_ (.A1(_06005_),
    .A2(_06047_),
    .A3(_06048_),
    .B1(_06045_),
    .X(_06050_));
 sky130_fd_sc_hd__nand2_1 _12188_ (.A(net959),
    .B(_06050_),
    .Y(_06051_));
 sky130_fd_sc_hd__o32a_1 _12189_ (.A1(net959),
    .A2(_06041_),
    .A3(_06042_),
    .B1(_06049_),
    .B2(_06051_),
    .X(_06052_));
 sky130_fd_sc_hd__or3b_1 _12190_ (.A(_05994_),
    .B(_06011_),
    .C_N(_06018_),
    .X(_06053_));
 sky130_fd_sc_hd__a21oi_1 _12191_ (.A1(_06037_),
    .A2(_06053_),
    .B1(_06036_),
    .Y(_06054_));
 sky130_fd_sc_hd__a31o_1 _12192_ (.A1(_06036_),
    .A2(_06037_),
    .A3(_06053_),
    .B1(net839),
    .X(_06055_));
 sky130_fd_sc_hd__o22a_1 _12193_ (.A1(net955),
    .A2(_06052_),
    .B1(_06054_),
    .B2(_06055_),
    .X(_06056_));
 sky130_fd_sc_hd__mux2_1 _12194_ (.A0(_01204_),
    .A1(_06056_),
    .S(net202),
    .X(_06057_));
 sky130_fd_sc_hd__and2b_1 _12195_ (.A_N(_06057_),
    .B(net1191),
    .X(_01152_));
 sky130_fd_sc_hd__nor2_1 _12196_ (.A(_01203_),
    .B(net202),
    .Y(_06058_));
 sky130_fd_sc_hd__nand2_1 _12197_ (.A(net842),
    .B(\brancher.rPc_current_reg2[29] ),
    .Y(_06059_));
 sky130_fd_sc_hd__or2_1 _12198_ (.A(net842),
    .B(\brancher.rPc_current_reg2[29] ),
    .X(_06060_));
 sky130_fd_sc_hd__nand2_1 _12199_ (.A(_06059_),
    .B(_06060_),
    .Y(_06061_));
 sky130_fd_sc_hd__o21ai_1 _12200_ (.A1(_06036_),
    .A2(_06039_),
    .B1(_06034_),
    .Y(_06062_));
 sky130_fd_sc_hd__xnor2_1 _12201_ (.A(_06061_),
    .B(_06062_),
    .Y(_06063_));
 sky130_fd_sc_hd__xnor2_1 _12202_ (.A(_01203_),
    .B(_06032_),
    .Y(_06064_));
 sky130_fd_sc_hd__mux2_1 _12203_ (.A0(_06064_),
    .A1(_06063_),
    .S(net178),
    .X(_06065_));
 sky130_fd_sc_hd__and2_1 _12204_ (.A(net946),
    .B(_01928_),
    .X(_06066_));
 sky130_fd_sc_hd__nand2_1 _12205_ (.A(net946),
    .B(_01928_),
    .Y(_06067_));
 sky130_fd_sc_hd__nor2_1 _12206_ (.A(net946),
    .B(_01928_),
    .Y(_06068_));
 sky130_fd_sc_hd__o211ai_1 _12207_ (.A1(_06066_),
    .A2(_06068_),
    .B1(_06043_),
    .C1(_06050_),
    .Y(_06069_));
 sky130_fd_sc_hd__a21o_1 _12208_ (.A1(_06043_),
    .A2(_06050_),
    .B1(_06068_),
    .X(_06070_));
 sky130_fd_sc_hd__o2111a_1 _12209_ (.A1(_06066_),
    .A2(_06070_),
    .B1(_06069_),
    .C1(net838),
    .D1(net959),
    .X(_06071_));
 sky130_fd_sc_hd__a21o_1 _12210_ (.A1(net842),
    .A2(\brancher.rPc_current_reg2[28] ),
    .B1(_06054_),
    .X(_06072_));
 sky130_fd_sc_hd__xnor2_1 _12211_ (.A(_06061_),
    .B(_06072_),
    .Y(_06073_));
 sky130_fd_sc_hd__a21o_1 _12212_ (.A1(net954),
    .A2(_06073_),
    .B1(_05454_),
    .X(_06074_));
 sky130_fd_sc_hd__a211o_1 _12213_ (.A1(_03217_),
    .A2(_06065_),
    .B1(_06071_),
    .C1(_06074_),
    .X(_06075_));
 sky130_fd_sc_hd__o211a_1 _12214_ (.A1(net629),
    .A2(_06064_),
    .B1(_06075_),
    .C1(net202),
    .X(_06076_));
 sky130_fd_sc_hd__o21a_1 _12215_ (.A1(_06058_),
    .A2(_06076_),
    .B1(net1209),
    .X(_01153_));
 sky130_fd_sc_hd__and2_1 _12216_ (.A(net842),
    .B(\brancher.rPc_current_reg2[30] ),
    .X(_06077_));
 sky130_fd_sc_hd__nand2_1 _12217_ (.A(net842),
    .B(\brancher.rPc_current_reg2[30] ),
    .Y(_06078_));
 sky130_fd_sc_hd__nor2_1 _12218_ (.A(net842),
    .B(\brancher.rPc_current_reg2[30] ),
    .Y(_06079_));
 sky130_fd_sc_hd__nor2_1 _12219_ (.A(_06077_),
    .B(_06079_),
    .Y(_06080_));
 sky130_fd_sc_hd__and3_1 _12220_ (.A(_06034_),
    .B(_06037_),
    .C(_06059_),
    .X(_06081_));
 sky130_fd_sc_hd__or2_1 _12221_ (.A(_06036_),
    .B(_06061_),
    .X(_06082_));
 sky130_fd_sc_hd__o21ai_1 _12222_ (.A1(_06038_),
    .A2(_06082_),
    .B1(_06081_),
    .Y(_06083_));
 sky130_fd_sc_hd__xor2_1 _12223_ (.A(_06080_),
    .B(_06083_),
    .X(_06084_));
 sky130_fd_sc_hd__and3_1 _12224_ (.A(net158),
    .B(net156),
    .C(_06032_),
    .X(_06085_));
 sky130_fd_sc_hd__a21o_1 _12225_ (.A1(net156),
    .A2(_06032_),
    .B1(net158),
    .X(_06086_));
 sky130_fd_sc_hd__and2b_1 _12226_ (.A_N(_06085_),
    .B(_06086_),
    .X(_06087_));
 sky130_fd_sc_hd__mux2_1 _12227_ (.A0(_06087_),
    .A1(_06084_),
    .S(net178),
    .X(_06088_));
 sky130_fd_sc_hd__xnor2_1 _12228_ (.A(net946),
    .B(_01947_),
    .Y(_06089_));
 sky130_fd_sc_hd__and3_1 _12229_ (.A(_06067_),
    .B(_06070_),
    .C(_06089_),
    .X(_06090_));
 sky130_fd_sc_hd__a21oi_1 _12230_ (.A1(_06067_),
    .A2(_06070_),
    .B1(_06089_),
    .Y(_06091_));
 sky130_fd_sc_hd__o21ai_1 _12231_ (.A1(_06090_),
    .A2(_06091_),
    .B1(net958),
    .Y(_06092_));
 sky130_fd_sc_hd__o211a_1 _12232_ (.A1(net959),
    .A2(_06088_),
    .B1(_06092_),
    .C1(net838),
    .X(_06093_));
 sky130_fd_sc_hd__o21a_1 _12233_ (.A1(_06053_),
    .A2(_06082_),
    .B1(_06081_),
    .X(_06094_));
 sky130_fd_sc_hd__xnor2_1 _12234_ (.A(_06080_),
    .B(_06094_),
    .Y(_06095_));
 sky130_fd_sc_hd__a21o_1 _12235_ (.A1(net954),
    .A2(_06095_),
    .B1(_06093_),
    .X(_06096_));
 sky130_fd_sc_hd__mux2_1 _12236_ (.A0(net158),
    .A1(_06096_),
    .S(net202),
    .X(_06097_));
 sky130_fd_sc_hd__and2_1 _12237_ (.A(net1209),
    .B(_06097_),
    .X(_01154_));
 sky130_fd_sc_hd__xnor2_1 _12238_ (.A(net159),
    .B(_06085_),
    .Y(_06098_));
 sky130_fd_sc_hd__a21o_1 _12239_ (.A1(_06080_),
    .A2(_06083_),
    .B1(_06077_),
    .X(_06099_));
 sky130_fd_sc_hd__xor2_1 _12240_ (.A(net843),
    .B(\brancher.rPc_current_reg2[31] ),
    .X(_06100_));
 sky130_fd_sc_hd__xnor2_1 _12241_ (.A(_06099_),
    .B(_06100_),
    .Y(_06101_));
 sky130_fd_sc_hd__mux2_1 _12242_ (.A0(_06098_),
    .A1(_06101_),
    .S(_04045_),
    .X(_06102_));
 sky130_fd_sc_hd__a21oi_1 _12243_ (.A1(net947),
    .A2(_01947_),
    .B1(_06091_),
    .Y(_06103_));
 sky130_fd_sc_hd__xnor2_1 _12244_ (.A(_01219_),
    .B(_01969_),
    .Y(_06104_));
 sky130_fd_sc_hd__xnor2_1 _12245_ (.A(_06103_),
    .B(_06104_),
    .Y(_06105_));
 sky130_fd_sc_hd__mux2_1 _12246_ (.A0(_06102_),
    .A1(_06105_),
    .S(net960),
    .X(_06106_));
 sky130_fd_sc_hd__o21ai_1 _12247_ (.A1(_06079_),
    .A2(_06094_),
    .B1(_06078_),
    .Y(_06107_));
 sky130_fd_sc_hd__o21ai_1 _12248_ (.A1(_06100_),
    .A2(_06107_),
    .B1(net954),
    .Y(_06108_));
 sky130_fd_sc_hd__a21o_1 _12249_ (.A1(_06100_),
    .A2(_06107_),
    .B1(_06108_),
    .X(_06109_));
 sky130_fd_sc_hd__o21ai_1 _12250_ (.A1(\brancher.op_jal ),
    .A2(_06106_),
    .B1(_06109_),
    .Y(_06110_));
 sky130_fd_sc_hd__mux2_1 _12251_ (.A0(net159),
    .A1(_06110_),
    .S(net203),
    .X(_06111_));
 sky130_fd_sc_hd__and2_1 _12252_ (.A(net1200),
    .B(_06111_),
    .X(_01155_));
 sky130_fd_sc_hd__nand2_1 _12253_ (.A(_04046_),
    .B(net184),
    .Y(_06112_));
 sky130_fd_sc_hd__o211a_1 _12254_ (.A1(net953),
    .A2(net176),
    .B1(_05447_),
    .C1(net184),
    .X(_06113_));
 sky130_fd_sc_hd__a22o_1 _12255_ (.A1(net135),
    .A2(_06112_),
    .B1(_06113_),
    .B2(\brancher.rPc_current_reg2[0] ),
    .X(_06114_));
 sky130_fd_sc_hd__and2_1 _12256_ (.A(net1137),
    .B(_06114_),
    .X(_01156_));
 sky130_fd_sc_hd__a21oi_1 _12257_ (.A1(_05443_),
    .A2(_05444_),
    .B1(_05447_),
    .Y(_06115_));
 sky130_fd_sc_hd__and3_1 _12258_ (.A(_05445_),
    .B(net184),
    .C(_06115_),
    .X(_06116_));
 sky130_fd_sc_hd__a221o_1 _12259_ (.A1(net146),
    .A2(_06112_),
    .B1(_06113_),
    .B2(\brancher.rPc_current_reg2[1] ),
    .C1(_06116_),
    .X(_06117_));
 sky130_fd_sc_hd__and2_1 _12260_ (.A(net1137),
    .B(_06117_),
    .X(_01157_));
 sky130_fd_sc_hd__and2_1 _12261_ (.A(net1137),
    .B(_04046_),
    .X(_01158_));
 sky130_fd_sc_hd__a22o_1 _12262_ (.A1(\brancher.imm13_b[1] ),
    .A2(net256),
    .B1(net169),
    .B2(_04105_),
    .X(_01159_));
 sky130_fd_sc_hd__a22o_1 _12263_ (.A1(net1232),
    .A2(net256),
    .B1(net169),
    .B2(_04110_),
    .X(_01160_));
 sky130_fd_sc_hd__a21o_1 _12264_ (.A1(net1242),
    .A2(net255),
    .B1(_04115_),
    .X(_01161_));
 sky130_fd_sc_hd__a22o_1 _12265_ (.A1(\brancher.imm13_b[4] ),
    .A2(net256),
    .B1(net169),
    .B2(_04120_),
    .X(_01162_));
 sky130_fd_sc_hd__a21o_1 _12266_ (.A1(\brancher.imm13_b[5] ),
    .A2(net250),
    .B1(_04124_),
    .X(_01163_));
 sky130_fd_sc_hd__a21o_1 _12267_ (.A1(net1448),
    .A2(net250),
    .B1(_04126_),
    .X(_01164_));
 sky130_fd_sc_hd__a21o_1 _12268_ (.A1(\brancher.imm13_b[7] ),
    .A2(net250),
    .B1(_04128_),
    .X(_01165_));
 sky130_fd_sc_hd__a21o_1 _12269_ (.A1(net1449),
    .A2(net252),
    .B1(_04130_),
    .X(_01166_));
 sky130_fd_sc_hd__a21o_1 _12270_ (.A1(net1450),
    .A2(net252),
    .B1(_04132_),
    .X(_01167_));
 sky130_fd_sc_hd__a21o_1 _12271_ (.A1(\brancher.imm13_b[10] ),
    .A2(net259),
    .B1(_04134_),
    .X(_01168_));
 sky130_fd_sc_hd__a22o_1 _12272_ (.A1(\brancher.imm13_b[11] ),
    .A2(net256),
    .B1(net170),
    .B2(_04100_),
    .X(_01169_));
 sky130_fd_sc_hd__a21o_1 _12273_ (.A1(net840),
    .A2(net252),
    .B1(_04136_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _12274_ (.A0(net135),
    .A1(net1439),
    .S(net258),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _12275_ (.A0(net146),
    .A1(net1347),
    .S(net258),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _12276_ (.A0(net157),
    .A1(net1323),
    .S(net255),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _12277_ (.A0(net160),
    .A1(net1343),
    .S(net255),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _12278_ (.A0(net161),
    .A1(net1324),
    .S(net255),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _12279_ (.A0(net162),
    .A1(net1326),
    .S(net250),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _12280_ (.A0(net163),
    .A1(net1309),
    .S(net250),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _12281_ (.A0(net164),
    .A1(net1349),
    .S(net250),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _12282_ (.A0(net165),
    .A1(net1328),
    .S(net251),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _12283_ (.A0(net166),
    .A1(net1303),
    .S(net252),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _12284_ (.A0(net136),
    .A1(net1319),
    .S(net252),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _12285_ (.A0(net137),
    .A1(net1314),
    .S(net252),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _12286_ (.A0(net138),
    .A1(net1311),
    .S(net253),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _12287_ (.A0(net139),
    .A1(net1296),
    .S(net253),
    .X(_01184_));
 sky130_fd_sc_hd__mux2_1 _12288_ (.A0(net140),
    .A1(net1294),
    .S(net253),
    .X(_01185_));
 sky130_fd_sc_hd__mux2_1 _12289_ (.A0(net141),
    .A1(net1299),
    .S(net260),
    .X(_01186_));
 sky130_fd_sc_hd__mux2_1 _12290_ (.A0(net142),
    .A1(net1300),
    .S(net260),
    .X(_01187_));
 sky130_fd_sc_hd__mux2_1 _12291_ (.A0(net143),
    .A1(net1295),
    .S(net260),
    .X(_01188_));
 sky130_fd_sc_hd__mux2_1 _12292_ (.A0(net144),
    .A1(net1313),
    .S(net260),
    .X(_01189_));
 sky130_fd_sc_hd__mux2_1 _12293_ (.A0(net145),
    .A1(net1306),
    .S(net260),
    .X(_01190_));
 sky130_fd_sc_hd__mux2_1 _12294_ (.A0(net147),
    .A1(net1341),
    .S(net260),
    .X(_01191_));
 sky130_fd_sc_hd__mux2_1 _12295_ (.A0(net148),
    .A1(net1345),
    .S(net261),
    .X(_01192_));
 sky130_fd_sc_hd__mux2_1 _12296_ (.A0(net149),
    .A1(net1317),
    .S(net261),
    .X(_01193_));
 sky130_fd_sc_hd__mux2_1 _12297_ (.A0(net150),
    .A1(net1308),
    .S(net261),
    .X(_01194_));
 sky130_fd_sc_hd__mux2_1 _12298_ (.A0(net151),
    .A1(net1336),
    .S(net262),
    .X(_01195_));
 sky130_fd_sc_hd__mux2_1 _12299_ (.A0(net152),
    .A1(net1338),
    .S(net262),
    .X(_01196_));
 sky130_fd_sc_hd__mux2_1 _12300_ (.A0(net153),
    .A1(net1433),
    .S(net261),
    .X(_01197_));
 sky130_fd_sc_hd__mux2_1 _12301_ (.A0(net154),
    .A1(net1344),
    .S(net262),
    .X(_01198_));
 sky130_fd_sc_hd__mux2_1 _12302_ (.A0(net155),
    .A1(net1330),
    .S(net261),
    .X(_01199_));
 sky130_fd_sc_hd__mux2_1 _12303_ (.A0(net1340),
    .A1(net1332),
    .S(net263),
    .X(_01200_));
 sky130_fd_sc_hd__mux2_1 _12304_ (.A0(net158),
    .A1(net1255),
    .S(net263),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _12305_ (.A0(net159),
    .A1(net1251),
    .S(net263),
    .X(_01202_));
 sky130_fd_sc_hd__dfxtp_1 _12306_ (.CLK(clknet_leaf_40_clk),
    .D(_00034_),
    .Q(\brancher.imm21_j[19] ));
 sky130_fd_sc_hd__dfxtp_2 _12307_ (.CLK(clknet_leaf_40_clk),
    .D(_00035_),
    .Q(\brancher.imm21_j[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12308_ (.CLK(clknet_leaf_40_clk),
    .D(_00036_),
    .Q(\brancher.imm21_j[16] ));
 sky130_fd_sc_hd__dfxtp_2 _12309_ (.CLK(clknet_leaf_40_clk),
    .D(_00037_),
    .Q(\brancher.imm21_j[17] ));
 sky130_fd_sc_hd__dfxtp_2 _12310_ (.CLK(clknet_leaf_40_clk),
    .D(_00038_),
    .Q(\brancher.imm21_j[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12311_ (.CLK(clknet_leaf_33_clk),
    .D(net1259),
    .Q(rOp_memLd));
 sky130_fd_sc_hd__dfxtp_1 _12312_ (.CLK(clknet_leaf_33_clk),
    .D(net1213),
    .Q(rOp_memLd2));
 sky130_fd_sc_hd__dfxtp_2 _12313_ (.CLK(clknet_leaf_42_clk),
    .D(_00039_),
    .Q(\alu.r_type ));
 sky130_fd_sc_hd__dfxtp_1 _12314_ (.CLK(clknet_leaf_33_clk),
    .D(net1228),
    .Q(rRegWrEn2));
 sky130_fd_sc_hd__dfxtp_1 _12315_ (.CLK(clknet_leaf_45_clk),
    .D(_00002_),
    .Q(\rWrData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12316_ (.CLK(clknet_leaf_41_clk),
    .D(_00013_),
    .Q(\rWrData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12317_ (.CLK(clknet_leaf_45_clk),
    .D(_00024_),
    .Q(\rWrData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12318_ (.CLK(clknet_leaf_41_clk),
    .D(_00027_),
    .Q(\rWrData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12319_ (.CLK(clknet_leaf_45_clk),
    .D(_00028_),
    .Q(\rWrData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12320_ (.CLK(clknet_leaf_23_clk),
    .D(_00029_),
    .Q(\rWrData[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12321_ (.CLK(clknet_leaf_21_clk),
    .D(_00030_),
    .Q(\rWrData[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12322_ (.CLK(clknet_leaf_21_clk),
    .D(_00031_),
    .Q(\rWrData[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12323_ (.CLK(clknet_leaf_24_clk),
    .D(_00032_),
    .Q(\rWrData[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12324_ (.CLK(clknet_leaf_21_clk),
    .D(_00033_),
    .Q(\rWrData[9] ));
 sky130_fd_sc_hd__dfxtp_2 _12325_ (.CLK(clknet_leaf_18_clk),
    .D(_00003_),
    .Q(\rWrData[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12326_ (.CLK(clknet_leaf_18_clk),
    .D(_00004_),
    .Q(\rWrData[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12327_ (.CLK(clknet_leaf_18_clk),
    .D(_00005_),
    .Q(\rWrData[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12328_ (.CLK(clknet_leaf_17_clk),
    .D(_00006_),
    .Q(\rWrData[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12329_ (.CLK(clknet_leaf_19_clk),
    .D(_00007_),
    .Q(\rWrData[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12330_ (.CLK(clknet_leaf_50_clk),
    .D(_00008_),
    .Q(\rWrData[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12331_ (.CLK(clknet_leaf_52_clk),
    .D(_00009_),
    .Q(\rWrData[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12332_ (.CLK(clknet_leaf_76_clk),
    .D(_00010_),
    .Q(\rWrData[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12333_ (.CLK(clknet_leaf_76_clk),
    .D(_00011_),
    .Q(\rWrData[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12334_ (.CLK(clknet_leaf_76_clk),
    .D(_00012_),
    .Q(\rWrData[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12335_ (.CLK(clknet_leaf_76_clk),
    .D(_00014_),
    .Q(\rWrData[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12336_ (.CLK(clknet_leaf_61_clk),
    .D(_00015_),
    .Q(\rWrData[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12337_ (.CLK(clknet_leaf_71_clk),
    .D(_00016_),
    .Q(\rWrData[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12338_ (.CLK(clknet_leaf_78_clk),
    .D(_00017_),
    .Q(\rWrData[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12339_ (.CLK(clknet_leaf_82_clk),
    .D(_00018_),
    .Q(\rWrData[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12340_ (.CLK(clknet_leaf_70_clk),
    .D(_00019_),
    .Q(\rWrData[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12341_ (.CLK(clknet_leaf_73_clk),
    .D(_00020_),
    .Q(\rWrData[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12342_ (.CLK(clknet_leaf_78_clk),
    .D(_00021_),
    .Q(\rWrData[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12343_ (.CLK(clknet_leaf_82_clk),
    .D(_00022_),
    .Q(\rWrData[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12344_ (.CLK(clknet_leaf_82_clk),
    .D(_00023_),
    .Q(\rWrData[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12345_ (.CLK(clknet_leaf_61_clk),
    .D(_00025_),
    .Q(\rWrData[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12346_ (.CLK(clknet_leaf_61_clk),
    .D(_00026_),
    .Q(\rWrData[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12347_ (.CLK(clknet_leaf_46_clk),
    .D(net1229),
    .Q(\rWrDataWB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12348_ (.CLK(clknet_leaf_41_clk),
    .D(net1216),
    .Q(\rWrDataWB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12349_ (.CLK(clknet_leaf_45_clk),
    .D(net1218),
    .Q(\rWrDataWB[2] ));
 sky130_fd_sc_hd__dfxtp_2 _12350_ (.CLK(clknet_leaf_24_clk),
    .D(net1248),
    .Q(\rWrDataWB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12351_ (.CLK(clknet_leaf_41_clk),
    .D(net1234),
    .Q(\rWrDataWB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12352_ (.CLK(clknet_leaf_26_clk),
    .D(net1241),
    .Q(\rWrDataWB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12353_ (.CLK(clknet_leaf_26_clk),
    .D(net1243),
    .Q(\rWrDataWB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12354_ (.CLK(clknet_leaf_26_clk),
    .D(net1239),
    .Q(\rWrDataWB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12355_ (.CLK(clknet_leaf_24_clk),
    .D(net1225),
    .Q(\rWrDataWB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12356_ (.CLK(clknet_leaf_16_clk),
    .D(net1223),
    .Q(\rWrDataWB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12357_ (.CLK(clknet_leaf_12_clk),
    .D(net1247),
    .Q(\rWrDataWB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12358_ (.CLK(clknet_leaf_118_clk),
    .D(net1238),
    .Q(\rWrDataWB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12359_ (.CLK(clknet_leaf_18_clk),
    .D(net1214),
    .Q(\rWrDataWB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12360_ (.CLK(clknet_leaf_17_clk),
    .D(net1222),
    .Q(\rWrDataWB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12361_ (.CLK(clknet_leaf_50_clk),
    .D(net1219),
    .Q(\rWrDataWB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12362_ (.CLK(clknet_leaf_76_clk),
    .D(net1227),
    .Q(\rWrDataWB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12363_ (.CLK(clknet_leaf_53_clk),
    .D(net1215),
    .Q(\rWrDataWB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12364_ (.CLK(clknet_leaf_76_clk),
    .D(net1246),
    .Q(\rWrDataWB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12365_ (.CLK(clknet_leaf_104_clk),
    .D(net1240),
    .Q(\rWrDataWB[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12366_ (.CLK(clknet_leaf_109_clk),
    .D(net1224),
    .Q(\rWrDataWB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12367_ (.CLK(clknet_leaf_111_clk),
    .D(net1226),
    .Q(\rWrDataWB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12368_ (.CLK(clknet_leaf_61_clk),
    .D(net1221),
    .Q(\rWrDataWB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12369_ (.CLK(clknet_leaf_71_clk),
    .D(net1220),
    .Q(\rWrDataWB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12370_ (.CLK(clknet_leaf_82_clk),
    .D(net1322),
    .Q(\rWrDataWB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12371_ (.CLK(clknet_leaf_81_clk),
    .D(net1211),
    .Q(\rWrDataWB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12372_ (.CLK(clknet_leaf_68_clk),
    .D(net1217),
    .Q(\rWrDataWB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12373_ (.CLK(clknet_leaf_74_clk),
    .D(net1233),
    .Q(\rWrDataWB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12374_ (.CLK(clknet_leaf_80_clk),
    .D(net1236),
    .Q(\rWrDataWB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12375_ (.CLK(clknet_leaf_83_clk),
    .D(net1212),
    .Q(\rWrDataWB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12376_ (.CLK(clknet_leaf_82_clk),
    .D(net1230),
    .Q(\rWrDataWB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12377_ (.CLK(clknet_leaf_82_clk),
    .D(net1321),
    .Q(\rWrDataWB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12378_ (.CLK(clknet_leaf_62_clk),
    .D(net1231),
    .Q(\rWrDataWB[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12379_ (.CLK(clknet_leaf_33_clk),
    .D(net1250),
    .Q(\rReg_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12380_ (.CLK(clknet_leaf_41_clk),
    .D(net1249),
    .Q(\rReg_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12381_ (.CLK(clknet_leaf_41_clk),
    .D(net1232),
    .Q(\rReg_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12382_ (.CLK(clknet_leaf_41_clk),
    .D(net1242),
    .Q(\rReg_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12383_ (.CLK(clknet_leaf_33_clk),
    .D(net1252),
    .Q(\rReg_d[4] ));
 sky130_fd_sc_hd__dfxtp_2 _12384_ (.CLK(clknet_leaf_33_clk),
    .D(net1235),
    .Q(\rReg_d2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12385_ (.CLK(clknet_leaf_33_clk),
    .D(net1245),
    .Q(\rReg_d2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12386_ (.CLK(clknet_leaf_33_clk),
    .D(net1256),
    .Q(\rReg_d2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12387_ (.CLK(clknet_leaf_33_clk),
    .D(net1244),
    .Q(\rReg_d2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12388_ (.CLK(clknet_leaf_33_clk),
    .D(net1237),
    .Q(\rReg_d2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12389_ (.CLK(clknet_leaf_24_clk),
    .D(_00000_),
    .Q(rHazardStallRs1));
 sky130_fd_sc_hd__dfxtp_1 _12390_ (.CLK(clknet_leaf_24_clk),
    .D(_00001_),
    .Q(rHazardStallRs2));
 sky130_fd_sc_hd__dfxtp_1 _12391_ (.CLK(clknet_leaf_41_clk),
    .D(_00040_),
    .Q(rRegWrEn));
 sky130_fd_sc_hd__dfxtp_1 _12392_ (.CLK(clknet_leaf_43_clk),
    .D(net257),
    .Q(\dec.rStall ));
 sky130_fd_sc_hd__dfxtp_1 _12393_ (.CLK(clknet_leaf_43_clk),
    .D(net34),
    .Q(\dec.rInstrustion[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12394_ (.CLK(clknet_leaf_43_clk),
    .D(net45),
    .Q(\dec.rInstrustion[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12395_ (.CLK(clknet_leaf_39_clk),
    .D(net56),
    .Q(\dec.rInstrustion[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12396_ (.CLK(clknet_leaf_43_clk),
    .D(net59),
    .Q(\dec.rInstrustion[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12397_ (.CLK(clknet_leaf_44_clk),
    .D(net60),
    .Q(\dec.rInstrustion[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12398_ (.CLK(clknet_leaf_44_clk),
    .D(net61),
    .Q(\dec.rInstrustion[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12399_ (.CLK(clknet_leaf_44_clk),
    .D(net62),
    .Q(\dec.rInstrustion[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12400_ (.CLK(clknet_leaf_39_clk),
    .D(net63),
    .Q(\dec.rInstrustion[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12401_ (.CLK(clknet_leaf_39_clk),
    .D(net64),
    .Q(\dec.rInstrustion[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12402_ (.CLK(clknet_leaf_39_clk),
    .D(net65),
    .Q(\dec.rInstrustion[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12403_ (.CLK(clknet_leaf_31_clk),
    .D(net35),
    .Q(\dec.rInstrustion[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12404_ (.CLK(clknet_leaf_38_clk),
    .D(net36),
    .Q(\dec.rInstrustion[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12405_ (.CLK(clknet_leaf_44_clk),
    .D(net37),
    .Q(\dec.rInstrustion[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12406_ (.CLK(clknet_leaf_44_clk),
    .D(net38),
    .Q(\dec.rInstrustion[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12407_ (.CLK(clknet_leaf_44_clk),
    .D(net39),
    .Q(\dec.rInstrustion[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12408_ (.CLK(clknet_leaf_38_clk),
    .D(net40),
    .Q(\dec.rInstrustion[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12409_ (.CLK(clknet_leaf_38_clk),
    .D(net41),
    .Q(\dec.rInstrustion[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12410_ (.CLK(clknet_leaf_38_clk),
    .D(net42),
    .Q(\dec.rInstrustion[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12411_ (.CLK(clknet_leaf_38_clk),
    .D(net43),
    .Q(\dec.rInstrustion[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12412_ (.CLK(clknet_leaf_38_clk),
    .D(net44),
    .Q(\dec.rInstrustion[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12413_ (.CLK(clknet_leaf_38_clk),
    .D(net46),
    .Q(\dec.rInstrustion[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12414_ (.CLK(clknet_leaf_39_clk),
    .D(net47),
    .Q(\dec.rInstrustion[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12415_ (.CLK(clknet_leaf_43_clk),
    .D(net48),
    .Q(\dec.rInstrustion[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12416_ (.CLK(clknet_leaf_36_clk),
    .D(net49),
    .Q(\dec.rInstrustion[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12417_ (.CLK(clknet_leaf_39_clk),
    .D(net50),
    .Q(\dec.rInstrustion[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12418_ (.CLK(clknet_leaf_30_clk),
    .D(net51),
    .Q(\dec.rInstrustion[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12419_ (.CLK(clknet_leaf_30_clk),
    .D(net52),
    .Q(\dec.rInstrustion[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12420_ (.CLK(clknet_leaf_30_clk),
    .D(net53),
    .Q(\dec.rInstrustion[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12421_ (.CLK(clknet_leaf_30_clk),
    .D(net54),
    .Q(\dec.rInstrustion[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12422_ (.CLK(clknet_leaf_30_clk),
    .D(net55),
    .Q(\dec.rInstrustion[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12423_ (.CLK(clknet_leaf_44_clk),
    .D(net57),
    .Q(\dec.rInstrustion[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12424_ (.CLK(clknet_leaf_30_clk),
    .D(net58),
    .Q(\dec.rInstrustion[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12425_ (.CLK(clknet_leaf_44_clk),
    .D(_00041_),
    .Q(\alu.op_consShf ));
 sky130_fd_sc_hd__dfxtp_1 _12426_ (.CLK(clknet_leaf_43_clk),
    .D(_00042_),
    .Q(\dec.op_memSt ));
 sky130_fd_sc_hd__dfxtp_1 _12427_ (.CLK(clknet_leaf_44_clk),
    .D(_00043_),
    .Q(\dec.op_intRegImm ));
 sky130_fd_sc_hd__dfxtp_2 _12428_ (.CLK(clknet_leaf_43_clk),
    .D(_00044_),
    .Q(\dec.op_memLd ));
 sky130_fd_sc_hd__dfxtp_2 _12429_ (.CLK(clknet_leaf_42_clk),
    .D(_00045_),
    .Q(\brancher.op_jalr ));
 sky130_fd_sc_hd__dfxtp_4 _12430_ (.CLK(clknet_leaf_43_clk),
    .D(_00046_),
    .Q(\brancher.op_jal ));
 sky130_fd_sc_hd__dfxtp_1 _12431_ (.CLK(clknet_leaf_42_clk),
    .D(_00047_),
    .Q(\dec.op_auipc ));
 sky130_fd_sc_hd__dfxtp_1 _12432_ (.CLK(clknet_leaf_42_clk),
    .D(_00048_),
    .Q(\dec.op_lui ));
 sky130_fd_sc_hd__dfxtp_2 _12433_ (.CLK(clknet_leaf_39_clk),
    .D(_00049_),
    .Q(\brancher.imm12_i_s[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12434_ (.CLK(clknet_leaf_42_clk),
    .D(_00050_),
    .Q(\brancher.imm12_i_s[1] ));
 sky130_fd_sc_hd__dfxtp_2 _12435_ (.CLK(clknet_leaf_42_clk),
    .D(_00051_),
    .Q(\brancher.imm12_i_s[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12436_ (.CLK(clknet_leaf_40_clk),
    .D(_00052_),
    .Q(\brancher.imm12_i_s[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12437_ (.CLK(clknet_leaf_40_clk),
    .D(_00053_),
    .Q(\brancher.imm12_i_s[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12438_ (.CLK(clknet_leaf_25_clk),
    .D(_00054_),
    .Q(\brancher.imm12_i_s[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12439_ (.CLK(clknet_leaf_23_clk),
    .D(_00055_),
    .Q(\brancher.imm12_i_s[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12440_ (.CLK(clknet_leaf_25_clk),
    .D(_00056_),
    .Q(\brancher.imm12_i_s[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12441_ (.CLK(clknet_leaf_24_clk),
    .D(_00057_),
    .Q(\brancher.imm12_i_s[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12442_ (.CLK(clknet_leaf_23_clk),
    .D(_00058_),
    .Q(\brancher.imm12_i_s[9] ));
 sky130_fd_sc_hd__dfxtp_2 _12443_ (.CLK(clknet_leaf_42_clk),
    .D(_00059_),
    .Q(\brancher.imm12_i_s[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12444_ (.CLK(clknet_leaf_23_clk),
    .D(_00060_),
    .Q(\brancher.imm12_i_s[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12445_ (.CLK(clknet_leaf_44_clk),
    .D(_00061_),
    .Q(\brancher.funct3[2] ));
 sky130_fd_sc_hd__dfxtp_2 _12446_ (.CLK(clknet_leaf_40_clk),
    .D(_00062_),
    .Q(\brancher.imm21_j[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12447_ (.CLK(clknet_leaf_39_clk),
    .D(_00063_),
    .Q(\brancher.imm21_j[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12448_ (.CLK(clknet_leaf_43_clk),
    .D(_00064_),
    .Q(\brancher.imm21_j[1] ));
 sky130_fd_sc_hd__dfxtp_4 _12449_ (.CLK(clknet_leaf_42_clk),
    .D(_00065_),
    .Q(\brancher.imm21_j[2] ));
 sky130_fd_sc_hd__dfxtp_2 _12450_ (.CLK(clknet_leaf_40_clk),
    .D(_00066_),
    .Q(\brancher.imm21_j[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12451_ (.CLK(clknet_leaf_44_clk),
    .D(_00067_),
    .Q(\brancher.funct3[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12452_ (.CLK(clknet_leaf_44_clk),
    .D(_00068_),
    .Q(\brancher.funct3[1] ));
 sky130_fd_sc_hd__dfxtp_4 _12453_ (.CLK(clknet_leaf_42_clk),
    .D(_00069_),
    .Q(\alu.b_type ));
 sky130_fd_sc_hd__dfxtp_1 _12454_ (.CLK(clknet_leaf_42_clk),
    .D(net1278),
    .Q(\brancher.rPc_current_reg2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12455_ (.CLK(clknet_leaf_42_clk),
    .D(net1285),
    .Q(\brancher.rPc_current_reg2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12456_ (.CLK(clknet_leaf_45_clk),
    .D(_00072_),
    .Q(\brancher.rPc_current_reg2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12457_ (.CLK(clknet_leaf_41_clk),
    .D(_00073_),
    .Q(\brancher.rPc_current_reg2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12458_ (.CLK(clknet_leaf_45_clk),
    .D(net1325),
    .Q(\brancher.rPc_current_reg2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12459_ (.CLK(clknet_leaf_24_clk),
    .D(net1327),
    .Q(\brancher.rPc_current_reg2[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12460_ (.CLK(clknet_leaf_22_clk),
    .D(net1310),
    .Q(\brancher.rPc_current_reg2[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12461_ (.CLK(clknet_leaf_23_clk),
    .D(net1282),
    .Q(\brancher.rPc_current_reg2[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12462_ (.CLK(clknet_leaf_23_clk),
    .D(net1329),
    .Q(\brancher.rPc_current_reg2[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12463_ (.CLK(clknet_leaf_23_clk),
    .D(net1304),
    .Q(\brancher.rPc_current_reg2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12464_ (.CLK(clknet_leaf_20_clk),
    .D(net1320),
    .Q(\brancher.rPc_current_reg2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12465_ (.CLK(clknet_leaf_20_clk),
    .D(net1302),
    .Q(\brancher.rPc_current_reg2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12466_ (.CLK(clknet_leaf_49_clk),
    .D(net1312),
    .Q(\brancher.rPc_current_reg2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12467_ (.CLK(clknet_leaf_48_clk),
    .D(net1297),
    .Q(\brancher.rPc_current_reg2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12468_ (.CLK(clknet_leaf_49_clk),
    .D(_00084_),
    .Q(\brancher.rPc_current_reg2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12469_ (.CLK(clknet_leaf_49_clk),
    .D(_00085_),
    .Q(\brancher.rPc_current_reg2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12470_ (.CLK(clknet_leaf_51_clk),
    .D(_00086_),
    .Q(\brancher.rPc_current_reg2[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12471_ (.CLK(clknet_leaf_51_clk),
    .D(_00087_),
    .Q(\brancher.rPc_current_reg2[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12472_ (.CLK(clknet_leaf_51_clk),
    .D(_00088_),
    .Q(\brancher.rPc_current_reg2[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12473_ (.CLK(clknet_leaf_51_clk),
    .D(_00089_),
    .Q(\brancher.rPc_current_reg2[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12474_ (.CLK(clknet_leaf_51_clk),
    .D(net1342),
    .Q(\brancher.rPc_current_reg2[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12475_ (.CLK(clknet_leaf_75_clk),
    .D(net1335),
    .Q(\brancher.rPc_current_reg2[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12476_ (.CLK(clknet_leaf_73_clk),
    .D(net1318),
    .Q(\brancher.rPc_current_reg2[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12477_ (.CLK(clknet_leaf_73_clk),
    .D(_00093_),
    .Q(\brancher.rPc_current_reg2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12478_ (.CLK(clknet_leaf_73_clk),
    .D(net1337),
    .Q(\brancher.rPc_current_reg2[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12479_ (.CLK(clknet_leaf_73_clk),
    .D(net1316),
    .Q(\brancher.rPc_current_reg2[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12480_ (.CLK(clknet_leaf_72_clk),
    .D(_00096_),
    .Q(\brancher.rPc_current_reg2[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12481_ (.CLK(clknet_leaf_73_clk),
    .D(_00097_),
    .Q(\brancher.rPc_current_reg2[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12482_ (.CLK(clknet_leaf_72_clk),
    .D(net1331),
    .Q(\brancher.rPc_current_reg2[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12483_ (.CLK(clknet_leaf_72_clk),
    .D(net1333),
    .Q(\brancher.rPc_current_reg2[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12484_ (.CLK(clknet_leaf_72_clk),
    .D(_00100_),
    .Q(\brancher.rPc_current_reg2[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12485_ (.CLK(clknet_leaf_72_clk),
    .D(_00101_),
    .Q(\brancher.rPc_current_reg2[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12486_ (.CLK(clknet_leaf_10_clk),
    .D(_00102_),
    .Q(\reg_module.gprf[0] ));
 sky130_fd_sc_hd__dfxtp_1 _12487_ (.CLK(clknet_leaf_36_clk),
    .D(_00103_),
    .Q(\reg_module.gprf[1] ));
 sky130_fd_sc_hd__dfxtp_1 _12488_ (.CLK(clknet_leaf_117_clk),
    .D(_00104_),
    .Q(\reg_module.gprf[2] ));
 sky130_fd_sc_hd__dfxtp_1 _12489_ (.CLK(clknet_leaf_3_clk),
    .D(_00105_),
    .Q(\reg_module.gprf[3] ));
 sky130_fd_sc_hd__dfxtp_1 _12490_ (.CLK(clknet_leaf_31_clk),
    .D(_00106_),
    .Q(\reg_module.gprf[4] ));
 sky130_fd_sc_hd__dfxtp_1 _12491_ (.CLK(clknet_leaf_8_clk),
    .D(_00107_),
    .Q(\reg_module.gprf[5] ));
 sky130_fd_sc_hd__dfxtp_1 _12492_ (.CLK(clknet_leaf_1_clk),
    .D(_00108_),
    .Q(\reg_module.gprf[6] ));
 sky130_fd_sc_hd__dfxtp_1 _12493_ (.CLK(clknet_leaf_6_clk),
    .D(_00109_),
    .Q(\reg_module.gprf[7] ));
 sky130_fd_sc_hd__dfxtp_1 _12494_ (.CLK(clknet_leaf_29_clk),
    .D(_00110_),
    .Q(\reg_module.gprf[8] ));
 sky130_fd_sc_hd__dfxtp_1 _12495_ (.CLK(clknet_leaf_124_clk),
    .D(_00111_),
    .Q(\reg_module.gprf[9] ));
 sky130_fd_sc_hd__dfxtp_1 _12496_ (.CLK(clknet_leaf_130_clk),
    .D(_00112_),
    .Q(\reg_module.gprf[10] ));
 sky130_fd_sc_hd__dfxtp_1 _12497_ (.CLK(clknet_leaf_122_clk),
    .D(_00113_),
    .Q(\reg_module.gprf[11] ));
 sky130_fd_sc_hd__dfxtp_1 _12498_ (.CLK(clknet_leaf_119_clk),
    .D(_00114_),
    .Q(\reg_module.gprf[12] ));
 sky130_fd_sc_hd__dfxtp_1 _12499_ (.CLK(clknet_leaf_126_clk),
    .D(_00115_),
    .Q(\reg_module.gprf[13] ));
 sky130_fd_sc_hd__dfxtp_1 _12500_ (.CLK(clknet_leaf_18_clk),
    .D(_00116_),
    .Q(\reg_module.gprf[14] ));
 sky130_fd_sc_hd__dfxtp_1 _12501_ (.CLK(clknet_leaf_109_clk),
    .D(_00117_),
    .Q(\reg_module.gprf[15] ));
 sky130_fd_sc_hd__dfxtp_1 _12502_ (.CLK(clknet_leaf_55_clk),
    .D(_00118_),
    .Q(\reg_module.gprf[16] ));
 sky130_fd_sc_hd__dfxtp_1 _12503_ (.CLK(clknet_leaf_103_clk),
    .D(_00119_),
    .Q(\reg_module.gprf[17] ));
 sky130_fd_sc_hd__dfxtp_1 _12504_ (.CLK(clknet_leaf_121_clk),
    .D(_00120_),
    .Q(\reg_module.gprf[18] ));
 sky130_fd_sc_hd__dfxtp_1 _12505_ (.CLK(clknet_leaf_107_clk),
    .D(_00121_),
    .Q(\reg_module.gprf[19] ));
 sky130_fd_sc_hd__dfxtp_1 _12506_ (.CLK(clknet_leaf_115_clk),
    .D(_00122_),
    .Q(\reg_module.gprf[20] ));
 sky130_fd_sc_hd__dfxtp_1 _12507_ (.CLK(clknet_leaf_58_clk),
    .D(_00123_),
    .Q(\reg_module.gprf[21] ));
 sky130_fd_sc_hd__dfxtp_1 _12508_ (.CLK(clknet_leaf_64_clk),
    .D(_00124_),
    .Q(\reg_module.gprf[22] ));
 sky130_fd_sc_hd__dfxtp_1 _12509_ (.CLK(clknet_leaf_96_clk),
    .D(_00125_),
    .Q(\reg_module.gprf[23] ));
 sky130_fd_sc_hd__dfxtp_1 _12510_ (.CLK(clknet_leaf_83_clk),
    .D(_00126_),
    .Q(\reg_module.gprf[24] ));
 sky130_fd_sc_hd__dfxtp_1 _12511_ (.CLK(clknet_leaf_90_clk),
    .D(_00127_),
    .Q(\reg_module.gprf[25] ));
 sky130_fd_sc_hd__dfxtp_1 _12512_ (.CLK(clknet_leaf_108_clk),
    .D(_00128_),
    .Q(\reg_module.gprf[26] ));
 sky130_fd_sc_hd__dfxtp_1 _12513_ (.CLK(clknet_leaf_96_clk),
    .D(_00129_),
    .Q(\reg_module.gprf[27] ));
 sky130_fd_sc_hd__dfxtp_1 _12514_ (.CLK(clknet_leaf_94_clk),
    .D(_00130_),
    .Q(\reg_module.gprf[28] ));
 sky130_fd_sc_hd__dfxtp_1 _12515_ (.CLK(clknet_leaf_80_clk),
    .D(_00131_),
    .Q(\reg_module.gprf[29] ));
 sky130_fd_sc_hd__dfxtp_1 _12516_ (.CLK(clknet_leaf_67_clk),
    .D(_00132_),
    .Q(\reg_module.gprf[30] ));
 sky130_fd_sc_hd__dfxtp_1 _12517_ (.CLK(clknet_leaf_60_clk),
    .D(_00133_),
    .Q(\reg_module.gprf[31] ));
 sky130_fd_sc_hd__dfxtp_1 _12518_ (.CLK(clknet_leaf_10_clk),
    .D(_00134_),
    .Q(\reg_module.gprf[32] ));
 sky130_fd_sc_hd__dfxtp_1 _12519_ (.CLK(clknet_leaf_36_clk),
    .D(_00135_),
    .Q(\reg_module.gprf[33] ));
 sky130_fd_sc_hd__dfxtp_1 _12520_ (.CLK(clknet_leaf_117_clk),
    .D(_00136_),
    .Q(\reg_module.gprf[34] ));
 sky130_fd_sc_hd__dfxtp_1 _12521_ (.CLK(clknet_leaf_3_clk),
    .D(_00137_),
    .Q(\reg_module.gprf[35] ));
 sky130_fd_sc_hd__dfxtp_1 _12522_ (.CLK(clknet_leaf_30_clk),
    .D(_00138_),
    .Q(\reg_module.gprf[36] ));
 sky130_fd_sc_hd__dfxtp_1 _12523_ (.CLK(clknet_leaf_8_clk),
    .D(_00139_),
    .Q(\reg_module.gprf[37] ));
 sky130_fd_sc_hd__dfxtp_1 _12524_ (.CLK(clknet_leaf_1_clk),
    .D(_00140_),
    .Q(\reg_module.gprf[38] ));
 sky130_fd_sc_hd__dfxtp_1 _12525_ (.CLK(clknet_leaf_6_clk),
    .D(_00141_),
    .Q(\reg_module.gprf[39] ));
 sky130_fd_sc_hd__dfxtp_1 _12526_ (.CLK(clknet_leaf_29_clk),
    .D(_00142_),
    .Q(\reg_module.gprf[40] ));
 sky130_fd_sc_hd__dfxtp_1 _12527_ (.CLK(clknet_leaf_125_clk),
    .D(_00143_),
    .Q(\reg_module.gprf[41] ));
 sky130_fd_sc_hd__dfxtp_1 _12528_ (.CLK(clknet_leaf_128_clk),
    .D(_00144_),
    .Q(\reg_module.gprf[42] ));
 sky130_fd_sc_hd__dfxtp_1 _12529_ (.CLK(clknet_leaf_122_clk),
    .D(_00145_),
    .Q(\reg_module.gprf[43] ));
 sky130_fd_sc_hd__dfxtp_1 _12530_ (.CLK(clknet_leaf_120_clk),
    .D(_00146_),
    .Q(\reg_module.gprf[44] ));
 sky130_fd_sc_hd__dfxtp_1 _12531_ (.CLK(clknet_leaf_126_clk),
    .D(_00147_),
    .Q(\reg_module.gprf[45] ));
 sky130_fd_sc_hd__dfxtp_1 _12532_ (.CLK(clknet_leaf_18_clk),
    .D(_00148_),
    .Q(\reg_module.gprf[46] ));
 sky130_fd_sc_hd__dfxtp_1 _12533_ (.CLK(clknet_leaf_110_clk),
    .D(_00149_),
    .Q(\reg_module.gprf[47] ));
 sky130_fd_sc_hd__dfxtp_1 _12534_ (.CLK(clknet_leaf_54_clk),
    .D(_00150_),
    .Q(\reg_module.gprf[48] ));
 sky130_fd_sc_hd__dfxtp_1 _12535_ (.CLK(clknet_leaf_103_clk),
    .D(_00151_),
    .Q(\reg_module.gprf[49] ));
 sky130_fd_sc_hd__dfxtp_1 _12536_ (.CLK(clknet_leaf_120_clk),
    .D(_00152_),
    .Q(\reg_module.gprf[50] ));
 sky130_fd_sc_hd__dfxtp_1 _12537_ (.CLK(clknet_leaf_98_clk),
    .D(_00153_),
    .Q(\reg_module.gprf[51] ));
 sky130_fd_sc_hd__dfxtp_1 _12538_ (.CLK(clknet_leaf_116_clk),
    .D(_00154_),
    .Q(\reg_module.gprf[52] ));
 sky130_fd_sc_hd__dfxtp_1 _12539_ (.CLK(clknet_leaf_60_clk),
    .D(_00155_),
    .Q(\reg_module.gprf[53] ));
 sky130_fd_sc_hd__dfxtp_1 _12540_ (.CLK(clknet_leaf_68_clk),
    .D(_00156_),
    .Q(\reg_module.gprf[54] ));
 sky130_fd_sc_hd__dfxtp_1 _12541_ (.CLK(clknet_leaf_96_clk),
    .D(_00157_),
    .Q(\reg_module.gprf[55] ));
 sky130_fd_sc_hd__dfxtp_1 _12542_ (.CLK(clknet_leaf_88_clk),
    .D(_00158_),
    .Q(\reg_module.gprf[56] ));
 sky130_fd_sc_hd__dfxtp_1 _12543_ (.CLK(clknet_leaf_90_clk),
    .D(_00159_),
    .Q(\reg_module.gprf[57] ));
 sky130_fd_sc_hd__dfxtp_1 _12544_ (.CLK(clknet_leaf_108_clk),
    .D(_00160_),
    .Q(\reg_module.gprf[58] ));
 sky130_fd_sc_hd__dfxtp_1 _12545_ (.CLK(clknet_leaf_99_clk),
    .D(_00161_),
    .Q(\reg_module.gprf[59] ));
 sky130_fd_sc_hd__dfxtp_1 _12546_ (.CLK(clknet_leaf_94_clk),
    .D(_00162_),
    .Q(\reg_module.gprf[60] ));
 sky130_fd_sc_hd__dfxtp_1 _12547_ (.CLK(clknet_leaf_107_clk),
    .D(_00163_),
    .Q(\reg_module.gprf[61] ));
 sky130_fd_sc_hd__dfxtp_1 _12548_ (.CLK(clknet_leaf_68_clk),
    .D(_00164_),
    .Q(\reg_module.gprf[62] ));
 sky130_fd_sc_hd__dfxtp_1 _12549_ (.CLK(clknet_leaf_61_clk),
    .D(_00165_),
    .Q(\reg_module.gprf[63] ));
 sky130_fd_sc_hd__dfxtp_1 _12550_ (.CLK(clknet_leaf_10_clk),
    .D(_00166_),
    .Q(\reg_module.gprf[64] ));
 sky130_fd_sc_hd__dfxtp_1 _12551_ (.CLK(clknet_leaf_36_clk),
    .D(_00167_),
    .Q(\reg_module.gprf[65] ));
 sky130_fd_sc_hd__dfxtp_1 _12552_ (.CLK(clknet_leaf_117_clk),
    .D(_00168_),
    .Q(\reg_module.gprf[66] ));
 sky130_fd_sc_hd__dfxtp_1 _12553_ (.CLK(clknet_leaf_2_clk),
    .D(_00169_),
    .Q(\reg_module.gprf[67] ));
 sky130_fd_sc_hd__dfxtp_1 _12554_ (.CLK(clknet_leaf_31_clk),
    .D(_00170_),
    .Q(\reg_module.gprf[68] ));
 sky130_fd_sc_hd__dfxtp_1 _12555_ (.CLK(clknet_leaf_8_clk),
    .D(_00171_),
    .Q(\reg_module.gprf[69] ));
 sky130_fd_sc_hd__dfxtp_1 _12556_ (.CLK(clknet_leaf_1_clk),
    .D(_00172_),
    .Q(\reg_module.gprf[70] ));
 sky130_fd_sc_hd__dfxtp_1 _12557_ (.CLK(clknet_leaf_6_clk),
    .D(_00173_),
    .Q(\reg_module.gprf[71] ));
 sky130_fd_sc_hd__dfxtp_1 _12558_ (.CLK(clknet_leaf_28_clk),
    .D(_00174_),
    .Q(\reg_module.gprf[72] ));
 sky130_fd_sc_hd__dfxtp_1 _12559_ (.CLK(clknet_leaf_125_clk),
    .D(_00175_),
    .Q(\reg_module.gprf[73] ));
 sky130_fd_sc_hd__dfxtp_1 _12560_ (.CLK(clknet_leaf_128_clk),
    .D(_00176_),
    .Q(\reg_module.gprf[74] ));
 sky130_fd_sc_hd__dfxtp_1 _12561_ (.CLK(clknet_leaf_122_clk),
    .D(_00177_),
    .Q(\reg_module.gprf[75] ));
 sky130_fd_sc_hd__dfxtp_1 _12562_ (.CLK(clknet_leaf_120_clk),
    .D(_00178_),
    .Q(\reg_module.gprf[76] ));
 sky130_fd_sc_hd__dfxtp_1 _12563_ (.CLK(clknet_leaf_126_clk),
    .D(_00179_),
    .Q(\reg_module.gprf[77] ));
 sky130_fd_sc_hd__dfxtp_1 _12564_ (.CLK(clknet_leaf_113_clk),
    .D(_00180_),
    .Q(\reg_module.gprf[78] ));
 sky130_fd_sc_hd__dfxtp_1 _12565_ (.CLK(clknet_leaf_110_clk),
    .D(_00181_),
    .Q(\reg_module.gprf[79] ));
 sky130_fd_sc_hd__dfxtp_1 _12566_ (.CLK(clknet_leaf_55_clk),
    .D(_00182_),
    .Q(\reg_module.gprf[80] ));
 sky130_fd_sc_hd__dfxtp_1 _12567_ (.CLK(clknet_leaf_103_clk),
    .D(_00183_),
    .Q(\reg_module.gprf[81] ));
 sky130_fd_sc_hd__dfxtp_1 _12568_ (.CLK(clknet_leaf_120_clk),
    .D(_00184_),
    .Q(\reg_module.gprf[82] ));
 sky130_fd_sc_hd__dfxtp_1 _12569_ (.CLK(clknet_leaf_98_clk),
    .D(_00185_),
    .Q(\reg_module.gprf[83] ));
 sky130_fd_sc_hd__dfxtp_1 _12570_ (.CLK(clknet_leaf_116_clk),
    .D(_00186_),
    .Q(\reg_module.gprf[84] ));
 sky130_fd_sc_hd__dfxtp_1 _12571_ (.CLK(clknet_leaf_58_clk),
    .D(_00187_),
    .Q(\reg_module.gprf[85] ));
 sky130_fd_sc_hd__dfxtp_1 _12572_ (.CLK(clknet_leaf_65_clk),
    .D(_00188_),
    .Q(\reg_module.gprf[86] ));
 sky130_fd_sc_hd__dfxtp_1 _12573_ (.CLK(clknet_leaf_96_clk),
    .D(_00189_),
    .Q(\reg_module.gprf[87] ));
 sky130_fd_sc_hd__dfxtp_1 _12574_ (.CLK(clknet_leaf_85_clk),
    .D(_00190_),
    .Q(\reg_module.gprf[88] ));
 sky130_fd_sc_hd__dfxtp_1 _12575_ (.CLK(clknet_leaf_90_clk),
    .D(_00191_),
    .Q(\reg_module.gprf[89] ));
 sky130_fd_sc_hd__dfxtp_1 _12576_ (.CLK(clknet_leaf_108_clk),
    .D(_00192_),
    .Q(\reg_module.gprf[90] ));
 sky130_fd_sc_hd__dfxtp_1 _12577_ (.CLK(clknet_leaf_98_clk),
    .D(_00193_),
    .Q(\reg_module.gprf[91] ));
 sky130_fd_sc_hd__dfxtp_1 _12578_ (.CLK(clknet_leaf_94_clk),
    .D(_00194_),
    .Q(\reg_module.gprf[92] ));
 sky130_fd_sc_hd__dfxtp_1 _12579_ (.CLK(clknet_leaf_80_clk),
    .D(_00195_),
    .Q(\reg_module.gprf[93] ));
 sky130_fd_sc_hd__dfxtp_1 _12580_ (.CLK(clknet_leaf_67_clk),
    .D(_00196_),
    .Q(\reg_module.gprf[94] ));
 sky130_fd_sc_hd__dfxtp_1 _12581_ (.CLK(clknet_leaf_60_clk),
    .D(_00197_),
    .Q(\reg_module.gprf[95] ));
 sky130_fd_sc_hd__dfxtp_1 _12582_ (.CLK(clknet_leaf_11_clk),
    .D(_00198_),
    .Q(\reg_module.gprf[96] ));
 sky130_fd_sc_hd__dfxtp_1 _12583_ (.CLK(clknet_leaf_34_clk),
    .D(_00199_),
    .Q(\reg_module.gprf[97] ));
 sky130_fd_sc_hd__dfxtp_1 _12584_ (.CLK(clknet_leaf_116_clk),
    .D(_00200_),
    .Q(\reg_module.gprf[98] ));
 sky130_fd_sc_hd__dfxtp_1 _12585_ (.CLK(clknet_leaf_3_clk),
    .D(_00201_),
    .Q(\reg_module.gprf[99] ));
 sky130_fd_sc_hd__dfxtp_1 _12586_ (.CLK(clknet_leaf_31_clk),
    .D(_00202_),
    .Q(\reg_module.gprf[100] ));
 sky130_fd_sc_hd__dfxtp_1 _12587_ (.CLK(clknet_leaf_8_clk),
    .D(_00203_),
    .Q(\reg_module.gprf[101] ));
 sky130_fd_sc_hd__dfxtp_1 _12588_ (.CLK(clknet_leaf_0_clk),
    .D(_00204_),
    .Q(\reg_module.gprf[102] ));
 sky130_fd_sc_hd__dfxtp_1 _12589_ (.CLK(clknet_leaf_5_clk),
    .D(_00205_),
    .Q(\reg_module.gprf[103] ));
 sky130_fd_sc_hd__dfxtp_1 _12590_ (.CLK(clknet_leaf_29_clk),
    .D(_00206_),
    .Q(\reg_module.gprf[104] ));
 sky130_fd_sc_hd__dfxtp_1 _12591_ (.CLK(clknet_leaf_123_clk),
    .D(_00207_),
    .Q(\reg_module.gprf[105] ));
 sky130_fd_sc_hd__dfxtp_1 _12592_ (.CLK(clknet_leaf_128_clk),
    .D(_00208_),
    .Q(\reg_module.gprf[106] ));
 sky130_fd_sc_hd__dfxtp_1 _12593_ (.CLK(clknet_leaf_121_clk),
    .D(_00209_),
    .Q(\reg_module.gprf[107] ));
 sky130_fd_sc_hd__dfxtp_1 _12594_ (.CLK(clknet_leaf_120_clk),
    .D(_00210_),
    .Q(\reg_module.gprf[108] ));
 sky130_fd_sc_hd__dfxtp_1 _12595_ (.CLK(clknet_leaf_126_clk),
    .D(_00211_),
    .Q(\reg_module.gprf[109] ));
 sky130_fd_sc_hd__dfxtp_1 _12596_ (.CLK(clknet_leaf_113_clk),
    .D(_00212_),
    .Q(\reg_module.gprf[110] ));
 sky130_fd_sc_hd__dfxtp_1 _12597_ (.CLK(clknet_leaf_108_clk),
    .D(_00213_),
    .Q(\reg_module.gprf[111] ));
 sky130_fd_sc_hd__dfxtp_1 _12598_ (.CLK(clknet_leaf_55_clk),
    .D(_00214_),
    .Q(\reg_module.gprf[112] ));
 sky130_fd_sc_hd__dfxtp_1 _12599_ (.CLK(clknet_leaf_101_clk),
    .D(_00215_),
    .Q(\reg_module.gprf[113] ));
 sky130_fd_sc_hd__dfxtp_1 _12600_ (.CLK(clknet_leaf_121_clk),
    .D(_00216_),
    .Q(\reg_module.gprf[114] ));
 sky130_fd_sc_hd__dfxtp_1 _12601_ (.CLK(clknet_leaf_98_clk),
    .D(_00217_),
    .Q(\reg_module.gprf[115] ));
 sky130_fd_sc_hd__dfxtp_1 _12602_ (.CLK(clknet_leaf_115_clk),
    .D(_00218_),
    .Q(\reg_module.gprf[116] ));
 sky130_fd_sc_hd__dfxtp_1 _12603_ (.CLK(clknet_leaf_58_clk),
    .D(_00219_),
    .Q(\reg_module.gprf[117] ));
 sky130_fd_sc_hd__dfxtp_1 _12604_ (.CLK(clknet_leaf_65_clk),
    .D(_00220_),
    .Q(\reg_module.gprf[118] ));
 sky130_fd_sc_hd__dfxtp_1 _12605_ (.CLK(clknet_leaf_96_clk),
    .D(_00221_),
    .Q(\reg_module.gprf[119] ));
 sky130_fd_sc_hd__dfxtp_1 _12606_ (.CLK(clknet_leaf_85_clk),
    .D(_00222_),
    .Q(\reg_module.gprf[120] ));
 sky130_fd_sc_hd__dfxtp_1 _12607_ (.CLK(clknet_leaf_90_clk),
    .D(_00223_),
    .Q(\reg_module.gprf[121] ));
 sky130_fd_sc_hd__dfxtp_1 _12608_ (.CLK(clknet_leaf_79_clk),
    .D(_00224_),
    .Q(\reg_module.gprf[122] ));
 sky130_fd_sc_hd__dfxtp_1 _12609_ (.CLK(clknet_leaf_96_clk),
    .D(_00225_),
    .Q(\reg_module.gprf[123] ));
 sky130_fd_sc_hd__dfxtp_1 _12610_ (.CLK(clknet_leaf_93_clk),
    .D(_00226_),
    .Q(\reg_module.gprf[124] ));
 sky130_fd_sc_hd__dfxtp_1 _12611_ (.CLK(clknet_leaf_80_clk),
    .D(_00227_),
    .Q(\reg_module.gprf[125] ));
 sky130_fd_sc_hd__dfxtp_1 _12612_ (.CLK(clknet_leaf_83_clk),
    .D(_00228_),
    .Q(\reg_module.gprf[126] ));
 sky130_fd_sc_hd__dfxtp_1 _12613_ (.CLK(clknet_leaf_63_clk),
    .D(_00229_),
    .Q(\reg_module.gprf[127] ));
 sky130_fd_sc_hd__dfxtp_1 _12614_ (.CLK(clknet_leaf_12_clk),
    .D(_00230_),
    .Q(\reg_module.gprf[128] ));
 sky130_fd_sc_hd__dfxtp_1 _12615_ (.CLK(clknet_leaf_35_clk),
    .D(_00231_),
    .Q(\reg_module.gprf[129] ));
 sky130_fd_sc_hd__dfxtp_1 _12616_ (.CLK(clknet_leaf_14_clk),
    .D(_00232_),
    .Q(\reg_module.gprf[130] ));
 sky130_fd_sc_hd__dfxtp_1 _12617_ (.CLK(clknet_leaf_3_clk),
    .D(_00233_),
    .Q(\reg_module.gprf[131] ));
 sky130_fd_sc_hd__dfxtp_1 _12618_ (.CLK(clknet_leaf_35_clk),
    .D(_00234_),
    .Q(\reg_module.gprf[132] ));
 sky130_fd_sc_hd__dfxtp_1 _12619_ (.CLK(clknet_leaf_28_clk),
    .D(_00235_),
    .Q(\reg_module.gprf[133] ));
 sky130_fd_sc_hd__dfxtp_1 _12620_ (.CLK(clknet_leaf_0_clk),
    .D(_00236_),
    .Q(\reg_module.gprf[134] ));
 sky130_fd_sc_hd__dfxtp_1 _12621_ (.CLK(clknet_leaf_6_clk),
    .D(_00237_),
    .Q(\reg_module.gprf[135] ));
 sky130_fd_sc_hd__dfxtp_1 _12622_ (.CLK(clknet_leaf_29_clk),
    .D(_00238_),
    .Q(\reg_module.gprf[136] ));
 sky130_fd_sc_hd__dfxtp_1 _12623_ (.CLK(clknet_leaf_126_clk),
    .D(_00239_),
    .Q(\reg_module.gprf[137] ));
 sky130_fd_sc_hd__dfxtp_1 _12624_ (.CLK(clknet_leaf_131_clk),
    .D(_00240_),
    .Q(\reg_module.gprf[138] ));
 sky130_fd_sc_hd__dfxtp_1 _12625_ (.CLK(clknet_leaf_120_clk),
    .D(_00241_),
    .Q(\reg_module.gprf[139] ));
 sky130_fd_sc_hd__dfxtp_1 _12626_ (.CLK(clknet_leaf_118_clk),
    .D(_00242_),
    .Q(\reg_module.gprf[140] ));
 sky130_fd_sc_hd__dfxtp_1 _12627_ (.CLK(clknet_leaf_117_clk),
    .D(_00243_),
    .Q(\reg_module.gprf[141] ));
 sky130_fd_sc_hd__dfxtp_1 _12628_ (.CLK(clknet_leaf_17_clk),
    .D(_00244_),
    .Q(\reg_module.gprf[142] ));
 sky130_fd_sc_hd__dfxtp_1 _12629_ (.CLK(clknet_leaf_110_clk),
    .D(_00245_),
    .Q(\reg_module.gprf[143] ));
 sky130_fd_sc_hd__dfxtp_1 _12630_ (.CLK(clknet_leaf_54_clk),
    .D(_00246_),
    .Q(\reg_module.gprf[144] ));
 sky130_fd_sc_hd__dfxtp_1 _12631_ (.CLK(clknet_leaf_104_clk),
    .D(_00247_),
    .Q(\reg_module.gprf[145] ));
 sky130_fd_sc_hd__dfxtp_1 _12632_ (.CLK(clknet_leaf_103_clk),
    .D(_00248_),
    .Q(\reg_module.gprf[146] ));
 sky130_fd_sc_hd__dfxtp_1 _12633_ (.CLK(clknet_leaf_106_clk),
    .D(_00249_),
    .Q(\reg_module.gprf[147] ));
 sky130_fd_sc_hd__dfxtp_1 _12634_ (.CLK(clknet_leaf_116_clk),
    .D(_00250_),
    .Q(\reg_module.gprf[148] ));
 sky130_fd_sc_hd__dfxtp_1 _12635_ (.CLK(clknet_leaf_60_clk),
    .D(_00251_),
    .Q(\reg_module.gprf[149] ));
 sky130_fd_sc_hd__dfxtp_1 _12636_ (.CLK(clknet_leaf_68_clk),
    .D(_00252_),
    .Q(\reg_module.gprf[150] ));
 sky130_fd_sc_hd__dfxtp_1 _12637_ (.CLK(clknet_leaf_97_clk),
    .D(_00253_),
    .Q(\reg_module.gprf[151] ));
 sky130_fd_sc_hd__dfxtp_1 _12638_ (.CLK(clknet_leaf_87_clk),
    .D(_00254_),
    .Q(\reg_module.gprf[152] ));
 sky130_fd_sc_hd__dfxtp_1 _12639_ (.CLK(clknet_leaf_87_clk),
    .D(_00255_),
    .Q(\reg_module.gprf[153] ));
 sky130_fd_sc_hd__dfxtp_1 _12640_ (.CLK(clknet_leaf_79_clk),
    .D(_00256_),
    .Q(\reg_module.gprf[154] ));
 sky130_fd_sc_hd__dfxtp_1 _12641_ (.CLK(clknet_leaf_99_clk),
    .D(_00257_),
    .Q(\reg_module.gprf[155] ));
 sky130_fd_sc_hd__dfxtp_1 _12642_ (.CLK(clknet_leaf_92_clk),
    .D(_00258_),
    .Q(\reg_module.gprf[156] ));
 sky130_fd_sc_hd__dfxtp_1 _12643_ (.CLK(clknet_leaf_107_clk),
    .D(_00259_),
    .Q(\reg_module.gprf[157] ));
 sky130_fd_sc_hd__dfxtp_1 _12644_ (.CLK(clknet_leaf_83_clk),
    .D(_00260_),
    .Q(\reg_module.gprf[158] ));
 sky130_fd_sc_hd__dfxtp_1 _12645_ (.CLK(clknet_leaf_62_clk),
    .D(_00261_),
    .Q(\reg_module.gprf[159] ));
 sky130_fd_sc_hd__dfxtp_1 _12646_ (.CLK(clknet_leaf_12_clk),
    .D(_00262_),
    .Q(\reg_module.gprf[160] ));
 sky130_fd_sc_hd__dfxtp_1 _12647_ (.CLK(clknet_leaf_35_clk),
    .D(_00263_),
    .Q(\reg_module.gprf[161] ));
 sky130_fd_sc_hd__dfxtp_1 _12648_ (.CLK(clknet_leaf_14_clk),
    .D(_00264_),
    .Q(\reg_module.gprf[162] ));
 sky130_fd_sc_hd__dfxtp_1 _12649_ (.CLK(clknet_leaf_2_clk),
    .D(_00265_),
    .Q(\reg_module.gprf[163] ));
 sky130_fd_sc_hd__dfxtp_1 _12650_ (.CLK(clknet_leaf_35_clk),
    .D(_00266_),
    .Q(\reg_module.gprf[164] ));
 sky130_fd_sc_hd__dfxtp_1 _12651_ (.CLK(clknet_leaf_8_clk),
    .D(_00267_),
    .Q(\reg_module.gprf[165] ));
 sky130_fd_sc_hd__dfxtp_1 _12652_ (.CLK(clknet_leaf_0_clk),
    .D(_00268_),
    .Q(\reg_module.gprf[166] ));
 sky130_fd_sc_hd__dfxtp_1 _12653_ (.CLK(clknet_leaf_5_clk),
    .D(_00269_),
    .Q(\reg_module.gprf[167] ));
 sky130_fd_sc_hd__dfxtp_1 _12654_ (.CLK(clknet_leaf_29_clk),
    .D(_00270_),
    .Q(\reg_module.gprf[168] ));
 sky130_fd_sc_hd__dfxtp_1 _12655_ (.CLK(clknet_leaf_125_clk),
    .D(_00271_),
    .Q(\reg_module.gprf[169] ));
 sky130_fd_sc_hd__dfxtp_1 _12656_ (.CLK(clknet_leaf_0_clk),
    .D(_00272_),
    .Q(\reg_module.gprf[170] ));
 sky130_fd_sc_hd__dfxtp_1 _12657_ (.CLK(clknet_leaf_120_clk),
    .D(_00273_),
    .Q(\reg_module.gprf[171] ));
 sky130_fd_sc_hd__dfxtp_1 _12658_ (.CLK(clknet_leaf_118_clk),
    .D(_00274_),
    .Q(\reg_module.gprf[172] ));
 sky130_fd_sc_hd__dfxtp_1 _12659_ (.CLK(clknet_leaf_126_clk),
    .D(_00275_),
    .Q(\reg_module.gprf[173] ));
 sky130_fd_sc_hd__dfxtp_1 _12660_ (.CLK(clknet_leaf_17_clk),
    .D(_00276_),
    .Q(\reg_module.gprf[174] ));
 sky130_fd_sc_hd__dfxtp_1 _12661_ (.CLK(clknet_leaf_110_clk),
    .D(_00277_),
    .Q(\reg_module.gprf[175] ));
 sky130_fd_sc_hd__dfxtp_1 _12662_ (.CLK(clknet_leaf_54_clk),
    .D(_00278_),
    .Q(\reg_module.gprf[176] ));
 sky130_fd_sc_hd__dfxtp_1 _12663_ (.CLK(clknet_leaf_104_clk),
    .D(_00279_),
    .Q(\reg_module.gprf[177] ));
 sky130_fd_sc_hd__dfxtp_1 _12664_ (.CLK(clknet_leaf_120_clk),
    .D(_00280_),
    .Q(\reg_module.gprf[178] ));
 sky130_fd_sc_hd__dfxtp_1 _12665_ (.CLK(clknet_leaf_106_clk),
    .D(_00281_),
    .Q(\reg_module.gprf[179] ));
 sky130_fd_sc_hd__dfxtp_1 _12666_ (.CLK(clknet_leaf_116_clk),
    .D(_00282_),
    .Q(\reg_module.gprf[180] ));
 sky130_fd_sc_hd__dfxtp_1 _12667_ (.CLK(clknet_leaf_60_clk),
    .D(_00283_),
    .Q(\reg_module.gprf[181] ));
 sky130_fd_sc_hd__dfxtp_1 _12668_ (.CLK(clknet_leaf_68_clk),
    .D(_00284_),
    .Q(\reg_module.gprf[182] ));
 sky130_fd_sc_hd__dfxtp_1 _12669_ (.CLK(clknet_leaf_97_clk),
    .D(_00285_),
    .Q(\reg_module.gprf[183] ));
 sky130_fd_sc_hd__dfxtp_1 _12670_ (.CLK(clknet_leaf_87_clk),
    .D(_00286_),
    .Q(\reg_module.gprf[184] ));
 sky130_fd_sc_hd__dfxtp_1 _12671_ (.CLK(clknet_leaf_87_clk),
    .D(_00287_),
    .Q(\reg_module.gprf[185] ));
 sky130_fd_sc_hd__dfxtp_1 _12672_ (.CLK(clknet_leaf_79_clk),
    .D(_00288_),
    .Q(\reg_module.gprf[186] ));
 sky130_fd_sc_hd__dfxtp_1 _12673_ (.CLK(clknet_leaf_99_clk),
    .D(_00289_),
    .Q(\reg_module.gprf[187] ));
 sky130_fd_sc_hd__dfxtp_1 _12674_ (.CLK(clknet_leaf_94_clk),
    .D(_00290_),
    .Q(\reg_module.gprf[188] ));
 sky130_fd_sc_hd__dfxtp_1 _12675_ (.CLK(clknet_leaf_98_clk),
    .D(_00291_),
    .Q(\reg_module.gprf[189] ));
 sky130_fd_sc_hd__dfxtp_1 _12676_ (.CLK(clknet_leaf_83_clk),
    .D(_00292_),
    .Q(\reg_module.gprf[190] ));
 sky130_fd_sc_hd__dfxtp_1 _12677_ (.CLK(clknet_leaf_62_clk),
    .D(_00293_),
    .Q(\reg_module.gprf[191] ));
 sky130_fd_sc_hd__dfxtp_1 _12678_ (.CLK(clknet_leaf_12_clk),
    .D(_00294_),
    .Q(\reg_module.gprf[192] ));
 sky130_fd_sc_hd__dfxtp_1 _12679_ (.CLK(clknet_leaf_34_clk),
    .D(_00295_),
    .Q(\reg_module.gprf[193] ));
 sky130_fd_sc_hd__dfxtp_1 _12680_ (.CLK(clknet_leaf_116_clk),
    .D(_00296_),
    .Q(\reg_module.gprf[194] ));
 sky130_fd_sc_hd__dfxtp_1 _12681_ (.CLK(clknet_leaf_3_clk),
    .D(_00297_),
    .Q(\reg_module.gprf[195] ));
 sky130_fd_sc_hd__dfxtp_1 _12682_ (.CLK(clknet_leaf_31_clk),
    .D(_00298_),
    .Q(\reg_module.gprf[196] ));
 sky130_fd_sc_hd__dfxtp_1 _12683_ (.CLK(clknet_leaf_9_clk),
    .D(_00299_),
    .Q(\reg_module.gprf[197] ));
 sky130_fd_sc_hd__dfxtp_1 _12684_ (.CLK(clknet_leaf_2_clk),
    .D(_00300_),
    .Q(\reg_module.gprf[198] ));
 sky130_fd_sc_hd__dfxtp_1 _12685_ (.CLK(clknet_leaf_4_clk),
    .D(_00301_),
    .Q(\reg_module.gprf[199] ));
 sky130_fd_sc_hd__dfxtp_1 _12686_ (.CLK(clknet_leaf_29_clk),
    .D(_00302_),
    .Q(\reg_module.gprf[200] ));
 sky130_fd_sc_hd__dfxtp_1 _12687_ (.CLK(clknet_leaf_125_clk),
    .D(_00303_),
    .Q(\reg_module.gprf[201] ));
 sky130_fd_sc_hd__dfxtp_1 _12688_ (.CLK(clknet_leaf_0_clk),
    .D(_00304_),
    .Q(\reg_module.gprf[202] ));
 sky130_fd_sc_hd__dfxtp_1 _12689_ (.CLK(clknet_leaf_120_clk),
    .D(_00305_),
    .Q(\reg_module.gprf[203] ));
 sky130_fd_sc_hd__dfxtp_1 _12690_ (.CLK(clknet_leaf_118_clk),
    .D(_00306_),
    .Q(\reg_module.gprf[204] ));
 sky130_fd_sc_hd__dfxtp_1 _12691_ (.CLK(clknet_leaf_118_clk),
    .D(_00307_),
    .Q(\reg_module.gprf[205] ));
 sky130_fd_sc_hd__dfxtp_1 _12692_ (.CLK(clknet_leaf_18_clk),
    .D(_00308_),
    .Q(\reg_module.gprf[206] ));
 sky130_fd_sc_hd__dfxtp_1 _12693_ (.CLK(clknet_leaf_110_clk),
    .D(_00309_),
    .Q(\reg_module.gprf[207] ));
 sky130_fd_sc_hd__dfxtp_1 _12694_ (.CLK(clknet_leaf_61_clk),
    .D(_00310_),
    .Q(\reg_module.gprf[208] ));
 sky130_fd_sc_hd__dfxtp_1 _12695_ (.CLK(clknet_leaf_103_clk),
    .D(_00311_),
    .Q(\reg_module.gprf[209] ));
 sky130_fd_sc_hd__dfxtp_1 _12696_ (.CLK(clknet_leaf_103_clk),
    .D(_00312_),
    .Q(\reg_module.gprf[210] ));
 sky130_fd_sc_hd__dfxtp_1 _12697_ (.CLK(clknet_leaf_107_clk),
    .D(_00313_),
    .Q(\reg_module.gprf[211] ));
 sky130_fd_sc_hd__dfxtp_1 _12698_ (.CLK(clknet_leaf_115_clk),
    .D(_00314_),
    .Q(\reg_module.gprf[212] ));
 sky130_fd_sc_hd__dfxtp_1 _12699_ (.CLK(clknet_leaf_60_clk),
    .D(_00315_),
    .Q(\reg_module.gprf[213] ));
 sky130_fd_sc_hd__dfxtp_1 _12700_ (.CLK(clknet_leaf_68_clk),
    .D(_00316_),
    .Q(\reg_module.gprf[214] ));
 sky130_fd_sc_hd__dfxtp_1 _12701_ (.CLK(clknet_leaf_97_clk),
    .D(_00317_),
    .Q(\reg_module.gprf[215] ));
 sky130_fd_sc_hd__dfxtp_1 _12702_ (.CLK(clknet_leaf_87_clk),
    .D(_00318_),
    .Q(\reg_module.gprf[216] ));
 sky130_fd_sc_hd__dfxtp_1 _12703_ (.CLK(clknet_leaf_91_clk),
    .D(_00319_),
    .Q(\reg_module.gprf[217] ));
 sky130_fd_sc_hd__dfxtp_1 _12704_ (.CLK(clknet_leaf_78_clk),
    .D(_00320_),
    .Q(\reg_module.gprf[218] ));
 sky130_fd_sc_hd__dfxtp_1 _12705_ (.CLK(clknet_leaf_99_clk),
    .D(_00321_),
    .Q(\reg_module.gprf[219] ));
 sky130_fd_sc_hd__dfxtp_1 _12706_ (.CLK(clknet_leaf_92_clk),
    .D(_00322_),
    .Q(\reg_module.gprf[220] ));
 sky130_fd_sc_hd__dfxtp_1 _12707_ (.CLK(clknet_leaf_89_clk),
    .D(_00323_),
    .Q(\reg_module.gprf[221] ));
 sky130_fd_sc_hd__dfxtp_1 _12708_ (.CLK(clknet_leaf_83_clk),
    .D(_00324_),
    .Q(\reg_module.gprf[222] ));
 sky130_fd_sc_hd__dfxtp_1 _12709_ (.CLK(clknet_leaf_62_clk),
    .D(_00325_),
    .Q(\reg_module.gprf[223] ));
 sky130_fd_sc_hd__dfxtp_1 _12710_ (.CLK(clknet_leaf_12_clk),
    .D(_00326_),
    .Q(\reg_module.gprf[224] ));
 sky130_fd_sc_hd__dfxtp_1 _12711_ (.CLK(clknet_leaf_34_clk),
    .D(_00327_),
    .Q(\reg_module.gprf[225] ));
 sky130_fd_sc_hd__dfxtp_1 _12712_ (.CLK(clknet_leaf_117_clk),
    .D(_00328_),
    .Q(\reg_module.gprf[226] ));
 sky130_fd_sc_hd__dfxtp_1 _12713_ (.CLK(clknet_leaf_127_clk),
    .D(_00329_),
    .Q(\reg_module.gprf[227] ));
 sky130_fd_sc_hd__dfxtp_1 _12714_ (.CLK(clknet_leaf_35_clk),
    .D(_00330_),
    .Q(\reg_module.gprf[228] ));
 sky130_fd_sc_hd__dfxtp_1 _12715_ (.CLK(clknet_leaf_9_clk),
    .D(_00331_),
    .Q(\reg_module.gprf[229] ));
 sky130_fd_sc_hd__dfxtp_1 _12716_ (.CLK(clknet_leaf_0_clk),
    .D(_00332_),
    .Q(\reg_module.gprf[230] ));
 sky130_fd_sc_hd__dfxtp_1 _12717_ (.CLK(clknet_leaf_4_clk),
    .D(_00333_),
    .Q(\reg_module.gprf[231] ));
 sky130_fd_sc_hd__dfxtp_1 _12718_ (.CLK(clknet_leaf_29_clk),
    .D(_00334_),
    .Q(\reg_module.gprf[232] ));
 sky130_fd_sc_hd__dfxtp_1 _12719_ (.CLK(clknet_leaf_125_clk),
    .D(_00335_),
    .Q(\reg_module.gprf[233] ));
 sky130_fd_sc_hd__dfxtp_1 _12720_ (.CLK(clknet_leaf_128_clk),
    .D(_00336_),
    .Q(\reg_module.gprf[234] ));
 sky130_fd_sc_hd__dfxtp_1 _12721_ (.CLK(clknet_leaf_120_clk),
    .D(_00337_),
    .Q(\reg_module.gprf[235] ));
 sky130_fd_sc_hd__dfxtp_1 _12722_ (.CLK(clknet_leaf_120_clk),
    .D(_00338_),
    .Q(\reg_module.gprf[236] ));
 sky130_fd_sc_hd__dfxtp_1 _12723_ (.CLK(clknet_leaf_118_clk),
    .D(_00339_),
    .Q(\reg_module.gprf[237] ));
 sky130_fd_sc_hd__dfxtp_1 _12724_ (.CLK(clknet_leaf_17_clk),
    .D(_00340_),
    .Q(\reg_module.gprf[238] ));
 sky130_fd_sc_hd__dfxtp_1 _12725_ (.CLK(clknet_leaf_110_clk),
    .D(_00341_),
    .Q(\reg_module.gprf[239] ));
 sky130_fd_sc_hd__dfxtp_1 _12726_ (.CLK(clknet_leaf_61_clk),
    .D(_00342_),
    .Q(\reg_module.gprf[240] ));
 sky130_fd_sc_hd__dfxtp_1 _12727_ (.CLK(clknet_leaf_104_clk),
    .D(_00343_),
    .Q(\reg_module.gprf[241] ));
 sky130_fd_sc_hd__dfxtp_1 _12728_ (.CLK(clknet_leaf_103_clk),
    .D(_00344_),
    .Q(\reg_module.gprf[242] ));
 sky130_fd_sc_hd__dfxtp_1 _12729_ (.CLK(clknet_leaf_107_clk),
    .D(_00345_),
    .Q(\reg_module.gprf[243] ));
 sky130_fd_sc_hd__dfxtp_1 _12730_ (.CLK(clknet_leaf_115_clk),
    .D(_00346_),
    .Q(\reg_module.gprf[244] ));
 sky130_fd_sc_hd__dfxtp_1 _12731_ (.CLK(clknet_leaf_59_clk),
    .D(_00347_),
    .Q(\reg_module.gprf[245] ));
 sky130_fd_sc_hd__dfxtp_1 _12732_ (.CLK(clknet_leaf_65_clk),
    .D(_00348_),
    .Q(\reg_module.gprf[246] ));
 sky130_fd_sc_hd__dfxtp_1 _12733_ (.CLK(clknet_leaf_97_clk),
    .D(_00349_),
    .Q(\reg_module.gprf[247] ));
 sky130_fd_sc_hd__dfxtp_1 _12734_ (.CLK(clknet_leaf_87_clk),
    .D(_00350_),
    .Q(\reg_module.gprf[248] ));
 sky130_fd_sc_hd__dfxtp_1 _12735_ (.CLK(clknet_leaf_87_clk),
    .D(_00351_),
    .Q(\reg_module.gprf[249] ));
 sky130_fd_sc_hd__dfxtp_1 _12736_ (.CLK(clknet_leaf_79_clk),
    .D(_00352_),
    .Q(\reg_module.gprf[250] ));
 sky130_fd_sc_hd__dfxtp_1 _12737_ (.CLK(clknet_leaf_99_clk),
    .D(_00353_),
    .Q(\reg_module.gprf[251] ));
 sky130_fd_sc_hd__dfxtp_1 _12738_ (.CLK(clknet_leaf_93_clk),
    .D(_00354_),
    .Q(\reg_module.gprf[252] ));
 sky130_fd_sc_hd__dfxtp_1 _12739_ (.CLK(clknet_leaf_98_clk),
    .D(_00355_),
    .Q(\reg_module.gprf[253] ));
 sky130_fd_sc_hd__dfxtp_1 _12740_ (.CLK(clknet_leaf_83_clk),
    .D(_00356_),
    .Q(\reg_module.gprf[254] ));
 sky130_fd_sc_hd__dfxtp_1 _12741_ (.CLK(clknet_leaf_64_clk),
    .D(_00357_),
    .Q(\reg_module.gprf[255] ));
 sky130_fd_sc_hd__dfxtp_1 _12742_ (.CLK(clknet_leaf_25_clk),
    .D(_00358_),
    .Q(\reg_module.gprf[256] ));
 sky130_fd_sc_hd__dfxtp_1 _12743_ (.CLK(clknet_leaf_36_clk),
    .D(_00359_),
    .Q(\reg_module.gprf[257] ));
 sky130_fd_sc_hd__dfxtp_1 _12744_ (.CLK(clknet_leaf_116_clk),
    .D(_00360_),
    .Q(\reg_module.gprf[258] ));
 sky130_fd_sc_hd__dfxtp_1 _12745_ (.CLK(clknet_leaf_3_clk),
    .D(_00361_),
    .Q(\reg_module.gprf[259] ));
 sky130_fd_sc_hd__dfxtp_1 _12746_ (.CLK(clknet_leaf_35_clk),
    .D(_00362_),
    .Q(\reg_module.gprf[260] ));
 sky130_fd_sc_hd__dfxtp_1 _12747_ (.CLK(clknet_leaf_28_clk),
    .D(_00363_),
    .Q(\reg_module.gprf[261] ));
 sky130_fd_sc_hd__dfxtp_1 _12748_ (.CLK(clknet_leaf_1_clk),
    .D(_00364_),
    .Q(\reg_module.gprf[262] ));
 sky130_fd_sc_hd__dfxtp_1 _12749_ (.CLK(clknet_leaf_6_clk),
    .D(_00365_),
    .Q(\reg_module.gprf[263] ));
 sky130_fd_sc_hd__dfxtp_1 _12750_ (.CLK(clknet_leaf_30_clk),
    .D(_00366_),
    .Q(\reg_module.gprf[264] ));
 sky130_fd_sc_hd__dfxtp_1 _12751_ (.CLK(clknet_leaf_124_clk),
    .D(_00367_),
    .Q(\reg_module.gprf[265] ));
 sky130_fd_sc_hd__dfxtp_1 _12752_ (.CLK(clknet_leaf_129_clk),
    .D(_00368_),
    .Q(\reg_module.gprf[266] ));
 sky130_fd_sc_hd__dfxtp_1 _12753_ (.CLK(clknet_leaf_121_clk),
    .D(_00369_),
    .Q(\reg_module.gprf[267] ));
 sky130_fd_sc_hd__dfxtp_1 _12754_ (.CLK(clknet_leaf_119_clk),
    .D(_00370_),
    .Q(\reg_module.gprf[268] ));
 sky130_fd_sc_hd__dfxtp_1 _12755_ (.CLK(clknet_leaf_117_clk),
    .D(_00371_),
    .Q(\reg_module.gprf[269] ));
 sky130_fd_sc_hd__dfxtp_1 _12756_ (.CLK(clknet_leaf_111_clk),
    .D(_00372_),
    .Q(\reg_module.gprf[270] ));
 sky130_fd_sc_hd__dfxtp_1 _12757_ (.CLK(clknet_leaf_108_clk),
    .D(_00373_),
    .Q(\reg_module.gprf[271] ));
 sky130_fd_sc_hd__dfxtp_1 _12758_ (.CLK(clknet_leaf_55_clk),
    .D(_00374_),
    .Q(\reg_module.gprf[272] ));
 sky130_fd_sc_hd__dfxtp_1 _12759_ (.CLK(clknet_leaf_102_clk),
    .D(_00375_),
    .Q(\reg_module.gprf[273] ));
 sky130_fd_sc_hd__dfxtp_1 _12760_ (.CLK(clknet_leaf_102_clk),
    .D(_00376_),
    .Q(\reg_module.gprf[274] ));
 sky130_fd_sc_hd__dfxtp_1 _12761_ (.CLK(clknet_leaf_107_clk),
    .D(_00377_),
    .Q(\reg_module.gprf[275] ));
 sky130_fd_sc_hd__dfxtp_1 _12762_ (.CLK(clknet_leaf_114_clk),
    .D(_00378_),
    .Q(\reg_module.gprf[276] ));
 sky130_fd_sc_hd__dfxtp_1 _12763_ (.CLK(clknet_leaf_58_clk),
    .D(_00379_),
    .Q(\reg_module.gprf[277] ));
 sky130_fd_sc_hd__dfxtp_1 _12764_ (.CLK(clknet_leaf_66_clk),
    .D(_00380_),
    .Q(\reg_module.gprf[278] ));
 sky130_fd_sc_hd__dfxtp_1 _12765_ (.CLK(clknet_leaf_94_clk),
    .D(_00381_),
    .Q(\reg_module.gprf[279] ));
 sky130_fd_sc_hd__dfxtp_1 _12766_ (.CLK(clknet_leaf_86_clk),
    .D(_00382_),
    .Q(\reg_module.gprf[280] ));
 sky130_fd_sc_hd__dfxtp_1 _12767_ (.CLK(clknet_leaf_91_clk),
    .D(_00383_),
    .Q(\reg_module.gprf[281] ));
 sky130_fd_sc_hd__dfxtp_1 _12768_ (.CLK(clknet_leaf_79_clk),
    .D(_00384_),
    .Q(\reg_module.gprf[282] ));
 sky130_fd_sc_hd__dfxtp_1 _12769_ (.CLK(clknet_leaf_96_clk),
    .D(_00385_),
    .Q(\reg_module.gprf[283] ));
 sky130_fd_sc_hd__dfxtp_1 _12770_ (.CLK(clknet_leaf_93_clk),
    .D(_00386_),
    .Q(\reg_module.gprf[284] ));
 sky130_fd_sc_hd__dfxtp_1 _12771_ (.CLK(clknet_leaf_81_clk),
    .D(_00387_),
    .Q(\reg_module.gprf[285] ));
 sky130_fd_sc_hd__dfxtp_1 _12772_ (.CLK(clknet_leaf_67_clk),
    .D(_00388_),
    .Q(\reg_module.gprf[286] ));
 sky130_fd_sc_hd__dfxtp_1 _12773_ (.CLK(clknet_leaf_63_clk),
    .D(_00389_),
    .Q(\reg_module.gprf[287] ));
 sky130_fd_sc_hd__dfxtp_1 _12774_ (.CLK(clknet_leaf_26_clk),
    .D(_00390_),
    .Q(\reg_module.gprf[288] ));
 sky130_fd_sc_hd__dfxtp_1 _12775_ (.CLK(clknet_leaf_36_clk),
    .D(_00391_),
    .Q(\reg_module.gprf[289] ));
 sky130_fd_sc_hd__dfxtp_1 _12776_ (.CLK(clknet_leaf_15_clk),
    .D(_00392_),
    .Q(\reg_module.gprf[290] ));
 sky130_fd_sc_hd__dfxtp_1 _12777_ (.CLK(clknet_leaf_3_clk),
    .D(_00393_),
    .Q(\reg_module.gprf[291] ));
 sky130_fd_sc_hd__dfxtp_1 _12778_ (.CLK(clknet_leaf_35_clk),
    .D(_00394_),
    .Q(\reg_module.gprf[292] ));
 sky130_fd_sc_hd__dfxtp_1 _12779_ (.CLK(clknet_leaf_28_clk),
    .D(_00395_),
    .Q(\reg_module.gprf[293] ));
 sky130_fd_sc_hd__dfxtp_1 _12780_ (.CLK(clknet_leaf_1_clk),
    .D(_00396_),
    .Q(\reg_module.gprf[294] ));
 sky130_fd_sc_hd__dfxtp_1 _12781_ (.CLK(clknet_leaf_7_clk),
    .D(_00397_),
    .Q(\reg_module.gprf[295] ));
 sky130_fd_sc_hd__dfxtp_1 _12782_ (.CLK(clknet_leaf_30_clk),
    .D(_00398_),
    .Q(\reg_module.gprf[296] ));
 sky130_fd_sc_hd__dfxtp_1 _12783_ (.CLK(clknet_leaf_124_clk),
    .D(_00399_),
    .Q(\reg_module.gprf[297] ));
 sky130_fd_sc_hd__dfxtp_1 _12784_ (.CLK(clknet_leaf_130_clk),
    .D(_00400_),
    .Q(\reg_module.gprf[298] ));
 sky130_fd_sc_hd__dfxtp_1 _12785_ (.CLK(clknet_leaf_122_clk),
    .D(_00401_),
    .Q(\reg_module.gprf[299] ));
 sky130_fd_sc_hd__dfxtp_1 _12786_ (.CLK(clknet_leaf_119_clk),
    .D(_00402_),
    .Q(\reg_module.gprf[300] ));
 sky130_fd_sc_hd__dfxtp_1 _12787_ (.CLK(clknet_leaf_3_clk),
    .D(_00403_),
    .Q(\reg_module.gprf[301] ));
 sky130_fd_sc_hd__dfxtp_1 _12788_ (.CLK(clknet_leaf_112_clk),
    .D(_00404_),
    .Q(\reg_module.gprf[302] ));
 sky130_fd_sc_hd__dfxtp_1 _12789_ (.CLK(clknet_leaf_108_clk),
    .D(_00405_),
    .Q(\reg_module.gprf[303] ));
 sky130_fd_sc_hd__dfxtp_1 _12790_ (.CLK(clknet_leaf_55_clk),
    .D(_00406_),
    .Q(\reg_module.gprf[304] ));
 sky130_fd_sc_hd__dfxtp_1 _12791_ (.CLK(clknet_leaf_102_clk),
    .D(_00407_),
    .Q(\reg_module.gprf[305] ));
 sky130_fd_sc_hd__dfxtp_1 _12792_ (.CLK(clknet_leaf_102_clk),
    .D(_00408_),
    .Q(\reg_module.gprf[306] ));
 sky130_fd_sc_hd__dfxtp_1 _12793_ (.CLK(clknet_leaf_107_clk),
    .D(_00409_),
    .Q(\reg_module.gprf[307] ));
 sky130_fd_sc_hd__dfxtp_1 _12794_ (.CLK(clknet_leaf_114_clk),
    .D(_00410_),
    .Q(\reg_module.gprf[308] ));
 sky130_fd_sc_hd__dfxtp_1 _12795_ (.CLK(clknet_leaf_58_clk),
    .D(_00411_),
    .Q(\reg_module.gprf[309] ));
 sky130_fd_sc_hd__dfxtp_1 _12796_ (.CLK(clknet_leaf_65_clk),
    .D(_00412_),
    .Q(\reg_module.gprf[310] ));
 sky130_fd_sc_hd__dfxtp_1 _12797_ (.CLK(clknet_leaf_95_clk),
    .D(_00413_),
    .Q(\reg_module.gprf[311] ));
 sky130_fd_sc_hd__dfxtp_1 _12798_ (.CLK(clknet_leaf_85_clk),
    .D(_00414_),
    .Q(\reg_module.gprf[312] ));
 sky130_fd_sc_hd__dfxtp_1 _12799_ (.CLK(clknet_leaf_91_clk),
    .D(_00415_),
    .Q(\reg_module.gprf[313] ));
 sky130_fd_sc_hd__dfxtp_1 _12800_ (.CLK(clknet_leaf_79_clk),
    .D(_00416_),
    .Q(\reg_module.gprf[314] ));
 sky130_fd_sc_hd__dfxtp_1 _12801_ (.CLK(clknet_leaf_100_clk),
    .D(_00417_),
    .Q(\reg_module.gprf[315] ));
 sky130_fd_sc_hd__dfxtp_1 _12802_ (.CLK(clknet_leaf_93_clk),
    .D(_00418_),
    .Q(\reg_module.gprf[316] ));
 sky130_fd_sc_hd__dfxtp_1 _12803_ (.CLK(clknet_leaf_82_clk),
    .D(_00419_),
    .Q(\reg_module.gprf[317] ));
 sky130_fd_sc_hd__dfxtp_1 _12804_ (.CLK(clknet_leaf_84_clk),
    .D(_00420_),
    .Q(\reg_module.gprf[318] ));
 sky130_fd_sc_hd__dfxtp_1 _12805_ (.CLK(clknet_leaf_63_clk),
    .D(_00421_),
    .Q(\reg_module.gprf[319] ));
 sky130_fd_sc_hd__dfxtp_1 _12806_ (.CLK(clknet_leaf_26_clk),
    .D(_00422_),
    .Q(\reg_module.gprf[320] ));
 sky130_fd_sc_hd__dfxtp_1 _12807_ (.CLK(clknet_leaf_37_clk),
    .D(_00423_),
    .Q(\reg_module.gprf[321] ));
 sky130_fd_sc_hd__dfxtp_1 _12808_ (.CLK(clknet_leaf_15_clk),
    .D(_00424_),
    .Q(\reg_module.gprf[322] ));
 sky130_fd_sc_hd__dfxtp_1 _12809_ (.CLK(clknet_leaf_13_clk),
    .D(_00425_),
    .Q(\reg_module.gprf[323] ));
 sky130_fd_sc_hd__dfxtp_1 _12810_ (.CLK(clknet_leaf_35_clk),
    .D(_00426_),
    .Q(\reg_module.gprf[324] ));
 sky130_fd_sc_hd__dfxtp_1 _12811_ (.CLK(clknet_leaf_28_clk),
    .D(_00427_),
    .Q(\reg_module.gprf[325] ));
 sky130_fd_sc_hd__dfxtp_1 _12812_ (.CLK(clknet_leaf_1_clk),
    .D(_00428_),
    .Q(\reg_module.gprf[326] ));
 sky130_fd_sc_hd__dfxtp_1 _12813_ (.CLK(clknet_leaf_7_clk),
    .D(_00429_),
    .Q(\reg_module.gprf[327] ));
 sky130_fd_sc_hd__dfxtp_1 _12814_ (.CLK(clknet_leaf_30_clk),
    .D(_00430_),
    .Q(\reg_module.gprf[328] ));
 sky130_fd_sc_hd__dfxtp_1 _12815_ (.CLK(clknet_leaf_124_clk),
    .D(_00431_),
    .Q(\reg_module.gprf[329] ));
 sky130_fd_sc_hd__dfxtp_1 _12816_ (.CLK(clknet_leaf_129_clk),
    .D(_00432_),
    .Q(\reg_module.gprf[330] ));
 sky130_fd_sc_hd__dfxtp_1 _12817_ (.CLK(clknet_leaf_122_clk),
    .D(_00433_),
    .Q(\reg_module.gprf[331] ));
 sky130_fd_sc_hd__dfxtp_1 _12818_ (.CLK(clknet_leaf_104_clk),
    .D(_00434_),
    .Q(\reg_module.gprf[332] ));
 sky130_fd_sc_hd__dfxtp_1 _12819_ (.CLK(clknet_leaf_14_clk),
    .D(_00435_),
    .Q(\reg_module.gprf[333] ));
 sky130_fd_sc_hd__dfxtp_1 _12820_ (.CLK(clknet_leaf_110_clk),
    .D(_00436_),
    .Q(\reg_module.gprf[334] ));
 sky130_fd_sc_hd__dfxtp_1 _12821_ (.CLK(clknet_leaf_108_clk),
    .D(_00437_),
    .Q(\reg_module.gprf[335] ));
 sky130_fd_sc_hd__dfxtp_1 _12822_ (.CLK(clknet_leaf_55_clk),
    .D(_00438_),
    .Q(\reg_module.gprf[336] ));
 sky130_fd_sc_hd__dfxtp_1 _12823_ (.CLK(clknet_leaf_102_clk),
    .D(_00439_),
    .Q(\reg_module.gprf[337] ));
 sky130_fd_sc_hd__dfxtp_1 _12824_ (.CLK(clknet_leaf_102_clk),
    .D(_00440_),
    .Q(\reg_module.gprf[338] ));
 sky130_fd_sc_hd__dfxtp_1 _12825_ (.CLK(clknet_leaf_80_clk),
    .D(_00441_),
    .Q(\reg_module.gprf[339] ));
 sky130_fd_sc_hd__dfxtp_1 _12826_ (.CLK(clknet_leaf_114_clk),
    .D(_00442_),
    .Q(\reg_module.gprf[340] ));
 sky130_fd_sc_hd__dfxtp_1 _12827_ (.CLK(clknet_leaf_58_clk),
    .D(_00443_),
    .Q(\reg_module.gprf[341] ));
 sky130_fd_sc_hd__dfxtp_1 _12828_ (.CLK(clknet_leaf_66_clk),
    .D(_00444_),
    .Q(\reg_module.gprf[342] ));
 sky130_fd_sc_hd__dfxtp_1 _12829_ (.CLK(clknet_leaf_95_clk),
    .D(_00445_),
    .Q(\reg_module.gprf[343] ));
 sky130_fd_sc_hd__dfxtp_1 _12830_ (.CLK(clknet_leaf_86_clk),
    .D(_00446_),
    .Q(\reg_module.gprf[344] ));
 sky130_fd_sc_hd__dfxtp_1 _12831_ (.CLK(clknet_leaf_91_clk),
    .D(_00447_),
    .Q(\reg_module.gprf[345] ));
 sky130_fd_sc_hd__dfxtp_1 _12832_ (.CLK(clknet_leaf_79_clk),
    .D(_00448_),
    .Q(\reg_module.gprf[346] ));
 sky130_fd_sc_hd__dfxtp_1 _12833_ (.CLK(clknet_leaf_100_clk),
    .D(_00449_),
    .Q(\reg_module.gprf[347] ));
 sky130_fd_sc_hd__dfxtp_1 _12834_ (.CLK(clknet_leaf_93_clk),
    .D(_00450_),
    .Q(\reg_module.gprf[348] ));
 sky130_fd_sc_hd__dfxtp_1 _12835_ (.CLK(clknet_leaf_81_clk),
    .D(_00451_),
    .Q(\reg_module.gprf[349] ));
 sky130_fd_sc_hd__dfxtp_1 _12836_ (.CLK(clknet_leaf_67_clk),
    .D(_00452_),
    .Q(\reg_module.gprf[350] ));
 sky130_fd_sc_hd__dfxtp_1 _12837_ (.CLK(clknet_leaf_63_clk),
    .D(_00453_),
    .Q(\reg_module.gprf[351] ));
 sky130_fd_sc_hd__dfxtp_1 _12838_ (.CLK(clknet_leaf_26_clk),
    .D(_00454_),
    .Q(\reg_module.gprf[352] ));
 sky130_fd_sc_hd__dfxtp_1 _12839_ (.CLK(clknet_leaf_37_clk),
    .D(_00455_),
    .Q(\reg_module.gprf[353] ));
 sky130_fd_sc_hd__dfxtp_1 _12840_ (.CLK(clknet_leaf_116_clk),
    .D(_00456_),
    .Q(\reg_module.gprf[354] ));
 sky130_fd_sc_hd__dfxtp_1 _12841_ (.CLK(clknet_leaf_14_clk),
    .D(_00457_),
    .Q(\reg_module.gprf[355] ));
 sky130_fd_sc_hd__dfxtp_1 _12842_ (.CLK(clknet_leaf_35_clk),
    .D(_00458_),
    .Q(\reg_module.gprf[356] ));
 sky130_fd_sc_hd__dfxtp_1 _12843_ (.CLK(clknet_leaf_28_clk),
    .D(_00459_),
    .Q(\reg_module.gprf[357] ));
 sky130_fd_sc_hd__dfxtp_1 _12844_ (.CLK(clknet_leaf_1_clk),
    .D(_00460_),
    .Q(\reg_module.gprf[358] ));
 sky130_fd_sc_hd__dfxtp_1 _12845_ (.CLK(clknet_leaf_7_clk),
    .D(_00461_),
    .Q(\reg_module.gprf[359] ));
 sky130_fd_sc_hd__dfxtp_1 _12846_ (.CLK(clknet_leaf_30_clk),
    .D(_00462_),
    .Q(\reg_module.gprf[360] ));
 sky130_fd_sc_hd__dfxtp_1 _12847_ (.CLK(clknet_leaf_124_clk),
    .D(_00463_),
    .Q(\reg_module.gprf[361] ));
 sky130_fd_sc_hd__dfxtp_1 _12848_ (.CLK(clknet_leaf_129_clk),
    .D(_00464_),
    .Q(\reg_module.gprf[362] ));
 sky130_fd_sc_hd__dfxtp_1 _12849_ (.CLK(clknet_leaf_121_clk),
    .D(_00465_),
    .Q(\reg_module.gprf[363] ));
 sky130_fd_sc_hd__dfxtp_1 _12850_ (.CLK(clknet_leaf_105_clk),
    .D(_00466_),
    .Q(\reg_module.gprf[364] ));
 sky130_fd_sc_hd__dfxtp_1 _12851_ (.CLK(clknet_leaf_117_clk),
    .D(_00467_),
    .Q(\reg_module.gprf[365] ));
 sky130_fd_sc_hd__dfxtp_1 _12852_ (.CLK(clknet_leaf_111_clk),
    .D(_00468_),
    .Q(\reg_module.gprf[366] ));
 sky130_fd_sc_hd__dfxtp_1 _12853_ (.CLK(clknet_leaf_108_clk),
    .D(_00469_),
    .Q(\reg_module.gprf[367] ));
 sky130_fd_sc_hd__dfxtp_1 _12854_ (.CLK(clknet_leaf_55_clk),
    .D(_00470_),
    .Q(\reg_module.gprf[368] ));
 sky130_fd_sc_hd__dfxtp_1 _12855_ (.CLK(clknet_leaf_100_clk),
    .D(_00471_),
    .Q(\reg_module.gprf[369] ));
 sky130_fd_sc_hd__dfxtp_1 _12856_ (.CLK(clknet_leaf_102_clk),
    .D(_00472_),
    .Q(\reg_module.gprf[370] ));
 sky130_fd_sc_hd__dfxtp_1 _12857_ (.CLK(clknet_leaf_80_clk),
    .D(_00473_),
    .Q(\reg_module.gprf[371] ));
 sky130_fd_sc_hd__dfxtp_1 _12858_ (.CLK(clknet_leaf_114_clk),
    .D(_00474_),
    .Q(\reg_module.gprf[372] ));
 sky130_fd_sc_hd__dfxtp_1 _12859_ (.CLK(clknet_leaf_58_clk),
    .D(_00475_),
    .Q(\reg_module.gprf[373] ));
 sky130_fd_sc_hd__dfxtp_1 _12860_ (.CLK(clknet_leaf_66_clk),
    .D(_00476_),
    .Q(\reg_module.gprf[374] ));
 sky130_fd_sc_hd__dfxtp_1 _12861_ (.CLK(clknet_leaf_94_clk),
    .D(_00477_),
    .Q(\reg_module.gprf[375] ));
 sky130_fd_sc_hd__dfxtp_1 _12862_ (.CLK(clknet_leaf_86_clk),
    .D(_00478_),
    .Q(\reg_module.gprf[376] ));
 sky130_fd_sc_hd__dfxtp_1 _12863_ (.CLK(clknet_leaf_91_clk),
    .D(_00479_),
    .Q(\reg_module.gprf[377] ));
 sky130_fd_sc_hd__dfxtp_1 _12864_ (.CLK(clknet_leaf_80_clk),
    .D(_00480_),
    .Q(\reg_module.gprf[378] ));
 sky130_fd_sc_hd__dfxtp_1 _12865_ (.CLK(clknet_leaf_95_clk),
    .D(_00481_),
    .Q(\reg_module.gprf[379] ));
 sky130_fd_sc_hd__dfxtp_1 _12866_ (.CLK(clknet_leaf_93_clk),
    .D(_00482_),
    .Q(\reg_module.gprf[380] ));
 sky130_fd_sc_hd__dfxtp_1 _12867_ (.CLK(clknet_leaf_81_clk),
    .D(_00483_),
    .Q(\reg_module.gprf[381] ));
 sky130_fd_sc_hd__dfxtp_1 _12868_ (.CLK(clknet_leaf_84_clk),
    .D(_00484_),
    .Q(\reg_module.gprf[382] ));
 sky130_fd_sc_hd__dfxtp_1 _12869_ (.CLK(clknet_leaf_63_clk),
    .D(_00485_),
    .Q(\reg_module.gprf[383] ));
 sky130_fd_sc_hd__dfxtp_1 _12870_ (.CLK(clknet_leaf_11_clk),
    .D(_00486_),
    .Q(\reg_module.gprf[384] ));
 sky130_fd_sc_hd__dfxtp_1 _12871_ (.CLK(clknet_leaf_40_clk),
    .D(_00487_),
    .Q(\reg_module.gprf[385] ));
 sky130_fd_sc_hd__dfxtp_1 _12872_ (.CLK(clknet_leaf_15_clk),
    .D(_00488_),
    .Q(\reg_module.gprf[386] ));
 sky130_fd_sc_hd__dfxtp_1 _12873_ (.CLK(clknet_leaf_13_clk),
    .D(_00489_),
    .Q(\reg_module.gprf[387] ));
 sky130_fd_sc_hd__dfxtp_1 _12874_ (.CLK(clknet_leaf_37_clk),
    .D(_00490_),
    .Q(\reg_module.gprf[388] ));
 sky130_fd_sc_hd__dfxtp_1 _12875_ (.CLK(clknet_leaf_28_clk),
    .D(_00491_),
    .Q(\reg_module.gprf[389] ));
 sky130_fd_sc_hd__dfxtp_1 _12876_ (.CLK(clknet_leaf_5_clk),
    .D(_00492_),
    .Q(\reg_module.gprf[390] ));
 sky130_fd_sc_hd__dfxtp_1 _12877_ (.CLK(clknet_leaf_7_clk),
    .D(_00493_),
    .Q(\reg_module.gprf[391] ));
 sky130_fd_sc_hd__dfxtp_1 _12878_ (.CLK(clknet_leaf_29_clk),
    .D(_00494_),
    .Q(\reg_module.gprf[392] ));
 sky130_fd_sc_hd__dfxtp_1 _12879_ (.CLK(clknet_leaf_129_clk),
    .D(_00495_),
    .Q(\reg_module.gprf[393] ));
 sky130_fd_sc_hd__dfxtp_1 _12880_ (.CLK(clknet_leaf_131_clk),
    .D(_00496_),
    .Q(\reg_module.gprf[394] ));
 sky130_fd_sc_hd__dfxtp_1 _12881_ (.CLK(clknet_leaf_123_clk),
    .D(_00497_),
    .Q(\reg_module.gprf[395] ));
 sky130_fd_sc_hd__dfxtp_1 _12882_ (.CLK(clknet_leaf_114_clk),
    .D(_00498_),
    .Q(\reg_module.gprf[396] ));
 sky130_fd_sc_hd__dfxtp_1 _12883_ (.CLK(clknet_leaf_127_clk),
    .D(_00499_),
    .Q(\reg_module.gprf[397] ));
 sky130_fd_sc_hd__dfxtp_1 _12884_ (.CLK(clknet_leaf_112_clk),
    .D(_00500_),
    .Q(\reg_module.gprf[398] ));
 sky130_fd_sc_hd__dfxtp_1 _12885_ (.CLK(clknet_leaf_77_clk),
    .D(_00501_),
    .Q(\reg_module.gprf[399] ));
 sky130_fd_sc_hd__dfxtp_1 _12886_ (.CLK(clknet_leaf_53_clk),
    .D(_00502_),
    .Q(\reg_module.gprf[400] ));
 sky130_fd_sc_hd__dfxtp_1 _12887_ (.CLK(clknet_leaf_101_clk),
    .D(_00503_),
    .Q(\reg_module.gprf[401] ));
 sky130_fd_sc_hd__dfxtp_1 _12888_ (.CLK(clknet_leaf_121_clk),
    .D(_00504_),
    .Q(\reg_module.gprf[402] ));
 sky130_fd_sc_hd__dfxtp_1 _12889_ (.CLK(clknet_leaf_106_clk),
    .D(_00505_),
    .Q(\reg_module.gprf[403] ));
 sky130_fd_sc_hd__dfxtp_1 _12890_ (.CLK(clknet_leaf_109_clk),
    .D(_00506_),
    .Q(\reg_module.gprf[404] ));
 sky130_fd_sc_hd__dfxtp_1 _12891_ (.CLK(clknet_leaf_55_clk),
    .D(_00507_),
    .Q(\reg_module.gprf[405] ));
 sky130_fd_sc_hd__dfxtp_1 _12892_ (.CLK(clknet_leaf_64_clk),
    .D(_00508_),
    .Q(\reg_module.gprf[406] ));
 sky130_fd_sc_hd__dfxtp_1 _12893_ (.CLK(clknet_leaf_96_clk),
    .D(_00509_),
    .Q(\reg_module.gprf[407] ));
 sky130_fd_sc_hd__dfxtp_1 _12894_ (.CLK(clknet_leaf_85_clk),
    .D(_00510_),
    .Q(\reg_module.gprf[408] ));
 sky130_fd_sc_hd__dfxtp_1 _12895_ (.CLK(clknet_leaf_87_clk),
    .D(_00511_),
    .Q(\reg_module.gprf[409] ));
 sky130_fd_sc_hd__dfxtp_1 _12896_ (.CLK(clknet_leaf_78_clk),
    .D(_00512_),
    .Q(\reg_module.gprf[410] ));
 sky130_fd_sc_hd__dfxtp_1 _12897_ (.CLK(clknet_leaf_99_clk),
    .D(_00513_),
    .Q(\reg_module.gprf[411] ));
 sky130_fd_sc_hd__dfxtp_1 _12898_ (.CLK(clknet_leaf_92_clk),
    .D(_00514_),
    .Q(\reg_module.gprf[412] ));
 sky130_fd_sc_hd__dfxtp_1 _12899_ (.CLK(clknet_leaf_80_clk),
    .D(_00515_),
    .Q(\reg_module.gprf[413] ));
 sky130_fd_sc_hd__dfxtp_1 _12900_ (.CLK(clknet_leaf_66_clk),
    .D(_00516_),
    .Q(\reg_module.gprf[414] ));
 sky130_fd_sc_hd__dfxtp_1 _12901_ (.CLK(clknet_leaf_59_clk),
    .D(_00517_),
    .Q(\reg_module.gprf[415] ));
 sky130_fd_sc_hd__dfxtp_1 _12902_ (.CLK(clknet_leaf_10_clk),
    .D(_00518_),
    .Q(\reg_module.gprf[416] ));
 sky130_fd_sc_hd__dfxtp_1 _12903_ (.CLK(clknet_leaf_37_clk),
    .D(_00519_),
    .Q(\reg_module.gprf[417] ));
 sky130_fd_sc_hd__dfxtp_1 _12904_ (.CLK(clknet_leaf_15_clk),
    .D(_00520_),
    .Q(\reg_module.gprf[418] ));
 sky130_fd_sc_hd__dfxtp_1 _12905_ (.CLK(clknet_leaf_13_clk),
    .D(_00521_),
    .Q(\reg_module.gprf[419] ));
 sky130_fd_sc_hd__dfxtp_1 _12906_ (.CLK(clknet_leaf_37_clk),
    .D(_00522_),
    .Q(\reg_module.gprf[420] ));
 sky130_fd_sc_hd__dfxtp_1 _12907_ (.CLK(clknet_leaf_28_clk),
    .D(_00523_),
    .Q(\reg_module.gprf[421] ));
 sky130_fd_sc_hd__dfxtp_1 _12908_ (.CLK(clknet_leaf_1_clk),
    .D(_00524_),
    .Q(\reg_module.gprf[422] ));
 sky130_fd_sc_hd__dfxtp_1 _12909_ (.CLK(clknet_leaf_7_clk),
    .D(_00525_),
    .Q(\reg_module.gprf[423] ));
 sky130_fd_sc_hd__dfxtp_1 _12910_ (.CLK(clknet_leaf_29_clk),
    .D(_00526_),
    .Q(\reg_module.gprf[424] ));
 sky130_fd_sc_hd__dfxtp_1 _12911_ (.CLK(clknet_leaf_129_clk),
    .D(_00527_),
    .Q(\reg_module.gprf[425] ));
 sky130_fd_sc_hd__dfxtp_1 _12912_ (.CLK(clknet_leaf_130_clk),
    .D(_00528_),
    .Q(\reg_module.gprf[426] ));
 sky130_fd_sc_hd__dfxtp_1 _12913_ (.CLK(clknet_leaf_123_clk),
    .D(_00529_),
    .Q(\reg_module.gprf[427] ));
 sky130_fd_sc_hd__dfxtp_1 _12914_ (.CLK(clknet_leaf_119_clk),
    .D(_00530_),
    .Q(\reg_module.gprf[428] ));
 sky130_fd_sc_hd__dfxtp_1 _12915_ (.CLK(clknet_leaf_127_clk),
    .D(_00531_),
    .Q(\reg_module.gprf[429] ));
 sky130_fd_sc_hd__dfxtp_1 _12916_ (.CLK(clknet_leaf_112_clk),
    .D(_00532_),
    .Q(\reg_module.gprf[430] ));
 sky130_fd_sc_hd__dfxtp_1 _12917_ (.CLK(clknet_leaf_77_clk),
    .D(_00533_),
    .Q(\reg_module.gprf[431] ));
 sky130_fd_sc_hd__dfxtp_1 _12918_ (.CLK(clknet_leaf_53_clk),
    .D(_00534_),
    .Q(\reg_module.gprf[432] ));
 sky130_fd_sc_hd__dfxtp_1 _12919_ (.CLK(clknet_leaf_101_clk),
    .D(_00535_),
    .Q(\reg_module.gprf[433] ));
 sky130_fd_sc_hd__dfxtp_1 _12920_ (.CLK(clknet_leaf_121_clk),
    .D(_00536_),
    .Q(\reg_module.gprf[434] ));
 sky130_fd_sc_hd__dfxtp_1 _12921_ (.CLK(clknet_leaf_109_clk),
    .D(_00537_),
    .Q(\reg_module.gprf[435] ));
 sky130_fd_sc_hd__dfxtp_1 _12922_ (.CLK(clknet_leaf_114_clk),
    .D(_00538_),
    .Q(\reg_module.gprf[436] ));
 sky130_fd_sc_hd__dfxtp_1 _12923_ (.CLK(clknet_leaf_55_clk),
    .D(_00539_),
    .Q(\reg_module.gprf[437] ));
 sky130_fd_sc_hd__dfxtp_1 _12924_ (.CLK(clknet_leaf_64_clk),
    .D(_00540_),
    .Q(\reg_module.gprf[438] ));
 sky130_fd_sc_hd__dfxtp_1 _12925_ (.CLK(clknet_leaf_94_clk),
    .D(_00541_),
    .Q(\reg_module.gprf[439] ));
 sky130_fd_sc_hd__dfxtp_1 _12926_ (.CLK(clknet_leaf_85_clk),
    .D(_00542_),
    .Q(\reg_module.gprf[440] ));
 sky130_fd_sc_hd__dfxtp_1 _12927_ (.CLK(clknet_leaf_87_clk),
    .D(_00543_),
    .Q(\reg_module.gprf[441] ));
 sky130_fd_sc_hd__dfxtp_1 _12928_ (.CLK(clknet_leaf_78_clk),
    .D(_00544_),
    .Q(\reg_module.gprf[442] ));
 sky130_fd_sc_hd__dfxtp_1 _12929_ (.CLK(clknet_leaf_99_clk),
    .D(_00545_),
    .Q(\reg_module.gprf[443] ));
 sky130_fd_sc_hd__dfxtp_1 _12930_ (.CLK(clknet_leaf_92_clk),
    .D(_00546_),
    .Q(\reg_module.gprf[444] ));
 sky130_fd_sc_hd__dfxtp_1 _12931_ (.CLK(clknet_leaf_80_clk),
    .D(_00547_),
    .Q(\reg_module.gprf[445] ));
 sky130_fd_sc_hd__dfxtp_1 _12932_ (.CLK(clknet_leaf_68_clk),
    .D(_00548_),
    .Q(\reg_module.gprf[446] ));
 sky130_fd_sc_hd__dfxtp_1 _12933_ (.CLK(clknet_leaf_59_clk),
    .D(_00549_),
    .Q(\reg_module.gprf[447] ));
 sky130_fd_sc_hd__dfxtp_1 _12934_ (.CLK(clknet_leaf_11_clk),
    .D(_00550_),
    .Q(\reg_module.gprf[448] ));
 sky130_fd_sc_hd__dfxtp_1 _12935_ (.CLK(clknet_leaf_40_clk),
    .D(_00551_),
    .Q(\reg_module.gprf[449] ));
 sky130_fd_sc_hd__dfxtp_1 _12936_ (.CLK(clknet_leaf_15_clk),
    .D(_00552_),
    .Q(\reg_module.gprf[450] ));
 sky130_fd_sc_hd__dfxtp_1 _12937_ (.CLK(clknet_leaf_13_clk),
    .D(_00553_),
    .Q(\reg_module.gprf[451] ));
 sky130_fd_sc_hd__dfxtp_1 _12938_ (.CLK(clknet_leaf_37_clk),
    .D(_00554_),
    .Q(\reg_module.gprf[452] ));
 sky130_fd_sc_hd__dfxtp_1 _12939_ (.CLK(clknet_leaf_27_clk),
    .D(_00555_),
    .Q(\reg_module.gprf[453] ));
 sky130_fd_sc_hd__dfxtp_1 _12940_ (.CLK(clknet_leaf_5_clk),
    .D(_00556_),
    .Q(\reg_module.gprf[454] ));
 sky130_fd_sc_hd__dfxtp_1 _12941_ (.CLK(clknet_leaf_10_clk),
    .D(_00557_),
    .Q(\reg_module.gprf[455] ));
 sky130_fd_sc_hd__dfxtp_1 _12942_ (.CLK(clknet_leaf_32_clk),
    .D(_00558_),
    .Q(\reg_module.gprf[456] ));
 sky130_fd_sc_hd__dfxtp_1 _12943_ (.CLK(clknet_leaf_124_clk),
    .D(_00559_),
    .Q(\reg_module.gprf[457] ));
 sky130_fd_sc_hd__dfxtp_1 _12944_ (.CLK(clknet_leaf_130_clk),
    .D(_00560_),
    .Q(\reg_module.gprf[458] ));
 sky130_fd_sc_hd__dfxtp_1 _12945_ (.CLK(clknet_leaf_122_clk),
    .D(_00561_),
    .Q(\reg_module.gprf[459] ));
 sky130_fd_sc_hd__dfxtp_1 _12946_ (.CLK(clknet_leaf_109_clk),
    .D(_00562_),
    .Q(\reg_module.gprf[460] ));
 sky130_fd_sc_hd__dfxtp_1 _12947_ (.CLK(clknet_leaf_126_clk),
    .D(_00563_),
    .Q(\reg_module.gprf[461] ));
 sky130_fd_sc_hd__dfxtp_1 _12948_ (.CLK(clknet_leaf_111_clk),
    .D(_00564_),
    .Q(\reg_module.gprf[462] ));
 sky130_fd_sc_hd__dfxtp_1 _12949_ (.CLK(clknet_leaf_77_clk),
    .D(_00565_),
    .Q(\reg_module.gprf[463] ));
 sky130_fd_sc_hd__dfxtp_1 _12950_ (.CLK(clknet_leaf_53_clk),
    .D(_00566_),
    .Q(\reg_module.gprf[464] ));
 sky130_fd_sc_hd__dfxtp_1 _12951_ (.CLK(clknet_leaf_101_clk),
    .D(_00567_),
    .Q(\reg_module.gprf[465] ));
 sky130_fd_sc_hd__dfxtp_1 _12952_ (.CLK(clknet_leaf_121_clk),
    .D(_00568_),
    .Q(\reg_module.gprf[466] ));
 sky130_fd_sc_hd__dfxtp_1 _12953_ (.CLK(clknet_leaf_106_clk),
    .D(_00569_),
    .Q(\reg_module.gprf[467] ));
 sky130_fd_sc_hd__dfxtp_1 _12954_ (.CLK(clknet_leaf_110_clk),
    .D(_00570_),
    .Q(\reg_module.gprf[468] ));
 sky130_fd_sc_hd__dfxtp_1 _12955_ (.CLK(clknet_leaf_58_clk),
    .D(_00571_),
    .Q(\reg_module.gprf[469] ));
 sky130_fd_sc_hd__dfxtp_1 _12956_ (.CLK(clknet_leaf_64_clk),
    .D(_00572_),
    .Q(\reg_module.gprf[470] ));
 sky130_fd_sc_hd__dfxtp_1 _12957_ (.CLK(clknet_leaf_94_clk),
    .D(_00573_),
    .Q(\reg_module.gprf[471] ));
 sky130_fd_sc_hd__dfxtp_1 _12958_ (.CLK(clknet_leaf_84_clk),
    .D(_00574_),
    .Q(\reg_module.gprf[472] ));
 sky130_fd_sc_hd__dfxtp_1 _12959_ (.CLK(clknet_leaf_86_clk),
    .D(_00575_),
    .Q(\reg_module.gprf[473] ));
 sky130_fd_sc_hd__dfxtp_1 _12960_ (.CLK(clknet_leaf_78_clk),
    .D(_00576_),
    .Q(\reg_module.gprf[474] ));
 sky130_fd_sc_hd__dfxtp_1 _12961_ (.CLK(clknet_leaf_100_clk),
    .D(_00577_),
    .Q(\reg_module.gprf[475] ));
 sky130_fd_sc_hd__dfxtp_1 _12962_ (.CLK(clknet_leaf_92_clk),
    .D(_00578_),
    .Q(\reg_module.gprf[476] ));
 sky130_fd_sc_hd__dfxtp_1 _12963_ (.CLK(clknet_leaf_80_clk),
    .D(_00579_),
    .Q(\reg_module.gprf[477] ));
 sky130_fd_sc_hd__dfxtp_1 _12964_ (.CLK(clknet_leaf_66_clk),
    .D(_00580_),
    .Q(\reg_module.gprf[478] ));
 sky130_fd_sc_hd__dfxtp_1 _12965_ (.CLK(clknet_leaf_59_clk),
    .D(_00581_),
    .Q(\reg_module.gprf[479] ));
 sky130_fd_sc_hd__dfxtp_1 _12966_ (.CLK(clknet_leaf_11_clk),
    .D(_00582_),
    .Q(\reg_module.gprf[480] ));
 sky130_fd_sc_hd__dfxtp_1 _12967_ (.CLK(clknet_leaf_40_clk),
    .D(_00583_),
    .Q(\reg_module.gprf[481] ));
 sky130_fd_sc_hd__dfxtp_1 _12968_ (.CLK(clknet_leaf_15_clk),
    .D(_00584_),
    .Q(\reg_module.gprf[482] ));
 sky130_fd_sc_hd__dfxtp_1 _12969_ (.CLK(clknet_leaf_13_clk),
    .D(_00585_),
    .Q(\reg_module.gprf[483] ));
 sky130_fd_sc_hd__dfxtp_1 _12970_ (.CLK(clknet_leaf_34_clk),
    .D(_00586_),
    .Q(\reg_module.gprf[484] ));
 sky130_fd_sc_hd__dfxtp_1 _12971_ (.CLK(clknet_leaf_27_clk),
    .D(_00587_),
    .Q(\reg_module.gprf[485] ));
 sky130_fd_sc_hd__dfxtp_1 _12972_ (.CLK(clknet_leaf_2_clk),
    .D(_00588_),
    .Q(\reg_module.gprf[486] ));
 sky130_fd_sc_hd__dfxtp_1 _12973_ (.CLK(clknet_leaf_12_clk),
    .D(_00589_),
    .Q(\reg_module.gprf[487] ));
 sky130_fd_sc_hd__dfxtp_1 _12974_ (.CLK(clknet_leaf_32_clk),
    .D(_00590_),
    .Q(\reg_module.gprf[488] ));
 sky130_fd_sc_hd__dfxtp_1 _12975_ (.CLK(clknet_leaf_125_clk),
    .D(_00591_),
    .Q(\reg_module.gprf[489] ));
 sky130_fd_sc_hd__dfxtp_1 _12976_ (.CLK(clknet_leaf_128_clk),
    .D(_00592_),
    .Q(\reg_module.gprf[490] ));
 sky130_fd_sc_hd__dfxtp_1 _12977_ (.CLK(clknet_leaf_122_clk),
    .D(_00593_),
    .Q(\reg_module.gprf[491] ));
 sky130_fd_sc_hd__dfxtp_1 _12978_ (.CLK(clknet_leaf_114_clk),
    .D(_00594_),
    .Q(\reg_module.gprf[492] ));
 sky130_fd_sc_hd__dfxtp_1 _12979_ (.CLK(clknet_leaf_117_clk),
    .D(_00595_),
    .Q(\reg_module.gprf[493] ));
 sky130_fd_sc_hd__dfxtp_1 _12980_ (.CLK(clknet_leaf_76_clk),
    .D(_00596_),
    .Q(\reg_module.gprf[494] ));
 sky130_fd_sc_hd__dfxtp_1 _12981_ (.CLK(clknet_leaf_76_clk),
    .D(_00597_),
    .Q(\reg_module.gprf[495] ));
 sky130_fd_sc_hd__dfxtp_1 _12982_ (.CLK(clknet_leaf_53_clk),
    .D(_00598_),
    .Q(\reg_module.gprf[496] ));
 sky130_fd_sc_hd__dfxtp_1 _12983_ (.CLK(clknet_leaf_101_clk),
    .D(_00599_),
    .Q(\reg_module.gprf[497] ));
 sky130_fd_sc_hd__dfxtp_1 _12984_ (.CLK(clknet_leaf_103_clk),
    .D(_00600_),
    .Q(\reg_module.gprf[498] ));
 sky130_fd_sc_hd__dfxtp_1 _12985_ (.CLK(clknet_leaf_105_clk),
    .D(_00601_),
    .Q(\reg_module.gprf[499] ));
 sky130_fd_sc_hd__dfxtp_1 _12986_ (.CLK(clknet_leaf_110_clk),
    .D(_00602_),
    .Q(\reg_module.gprf[500] ));
 sky130_fd_sc_hd__dfxtp_1 _12987_ (.CLK(clknet_leaf_55_clk),
    .D(_00603_),
    .Q(\reg_module.gprf[501] ));
 sky130_fd_sc_hd__dfxtp_1 _12988_ (.CLK(clknet_leaf_62_clk),
    .D(_00604_),
    .Q(\reg_module.gprf[502] ));
 sky130_fd_sc_hd__dfxtp_1 _12989_ (.CLK(clknet_leaf_94_clk),
    .D(_00605_),
    .Q(\reg_module.gprf[503] ));
 sky130_fd_sc_hd__dfxtp_1 _12990_ (.CLK(clknet_leaf_83_clk),
    .D(_00606_),
    .Q(\reg_module.gprf[504] ));
 sky130_fd_sc_hd__dfxtp_1 _12991_ (.CLK(clknet_leaf_87_clk),
    .D(_00607_),
    .Q(\reg_module.gprf[505] ));
 sky130_fd_sc_hd__dfxtp_1 _12992_ (.CLK(clknet_leaf_78_clk),
    .D(_00608_),
    .Q(\reg_module.gprf[506] ));
 sky130_fd_sc_hd__dfxtp_1 _12993_ (.CLK(clknet_leaf_99_clk),
    .D(_00609_),
    .Q(\reg_module.gprf[507] ));
 sky130_fd_sc_hd__dfxtp_1 _12994_ (.CLK(clknet_leaf_90_clk),
    .D(_00610_),
    .Q(\reg_module.gprf[508] ));
 sky130_fd_sc_hd__dfxtp_1 _12995_ (.CLK(clknet_leaf_81_clk),
    .D(_00611_),
    .Q(\reg_module.gprf[509] ));
 sky130_fd_sc_hd__dfxtp_1 _12996_ (.CLK(clknet_leaf_68_clk),
    .D(_00612_),
    .Q(\reg_module.gprf[510] ));
 sky130_fd_sc_hd__dfxtp_1 _12997_ (.CLK(clknet_leaf_59_clk),
    .D(_00613_),
    .Q(\reg_module.gprf[511] ));
 sky130_fd_sc_hd__dfxtp_1 _12998_ (.CLK(clknet_leaf_16_clk),
    .D(_00614_),
    .Q(\reg_module.gprf[512] ));
 sky130_fd_sc_hd__dfxtp_1 _12999_ (.CLK(clknet_leaf_40_clk),
    .D(_00615_),
    .Q(\reg_module.gprf[513] ));
 sky130_fd_sc_hd__dfxtp_1 _13000_ (.CLK(clknet_leaf_12_clk),
    .D(_00616_),
    .Q(\reg_module.gprf[514] ));
 sky130_fd_sc_hd__dfxtp_1 _13001_ (.CLK(clknet_leaf_4_clk),
    .D(_00617_),
    .Q(\reg_module.gprf[515] ));
 sky130_fd_sc_hd__dfxtp_1 _13002_ (.CLK(clknet_leaf_31_clk),
    .D(_00618_),
    .Q(\reg_module.gprf[516] ));
 sky130_fd_sc_hd__dfxtp_1 _13003_ (.CLK(clknet_leaf_27_clk),
    .D(_00619_),
    .Q(\reg_module.gprf[517] ));
 sky130_fd_sc_hd__dfxtp_1 _13004_ (.CLK(clknet_leaf_2_clk),
    .D(_00620_),
    .Q(\reg_module.gprf[518] ));
 sky130_fd_sc_hd__dfxtp_1 _13005_ (.CLK(clknet_leaf_10_clk),
    .D(_00621_),
    .Q(\reg_module.gprf[519] ));
 sky130_fd_sc_hd__dfxtp_1 _13006_ (.CLK(clknet_leaf_25_clk),
    .D(_00622_),
    .Q(\reg_module.gprf[520] ));
 sky130_fd_sc_hd__dfxtp_1 _13007_ (.CLK(clknet_leaf_126_clk),
    .D(_00623_),
    .Q(\reg_module.gprf[521] ));
 sky130_fd_sc_hd__dfxtp_1 _13008_ (.CLK(clknet_leaf_2_clk),
    .D(_00624_),
    .Q(\reg_module.gprf[522] ));
 sky130_fd_sc_hd__dfxtp_1 _13009_ (.CLK(clknet_leaf_120_clk),
    .D(_00625_),
    .Q(\reg_module.gprf[523] ));
 sky130_fd_sc_hd__dfxtp_1 _13010_ (.CLK(clknet_leaf_114_clk),
    .D(_00626_),
    .Q(\reg_module.gprf[524] ));
 sky130_fd_sc_hd__dfxtp_1 _13011_ (.CLK(clknet_leaf_117_clk),
    .D(_00627_),
    .Q(\reg_module.gprf[525] ));
 sky130_fd_sc_hd__dfxtp_1 _13012_ (.CLK(clknet_leaf_18_clk),
    .D(_00628_),
    .Q(\reg_module.gprf[526] ));
 sky130_fd_sc_hd__dfxtp_1 _13013_ (.CLK(clknet_leaf_76_clk),
    .D(_00629_),
    .Q(\reg_module.gprf[527] ));
 sky130_fd_sc_hd__dfxtp_1 _13014_ (.CLK(clknet_leaf_53_clk),
    .D(_00630_),
    .Q(\reg_module.gprf[528] ));
 sky130_fd_sc_hd__dfxtp_1 _13015_ (.CLK(clknet_leaf_106_clk),
    .D(_00631_),
    .Q(\reg_module.gprf[529] ));
 sky130_fd_sc_hd__dfxtp_1 _13016_ (.CLK(clknet_leaf_104_clk),
    .D(_00632_),
    .Q(\reg_module.gprf[530] ));
 sky130_fd_sc_hd__dfxtp_1 _13017_ (.CLK(clknet_leaf_105_clk),
    .D(_00633_),
    .Q(\reg_module.gprf[531] ));
 sky130_fd_sc_hd__dfxtp_1 _13018_ (.CLK(clknet_leaf_113_clk),
    .D(_00634_),
    .Q(\reg_module.gprf[532] ));
 sky130_fd_sc_hd__dfxtp_1 _13019_ (.CLK(clknet_leaf_55_clk),
    .D(_00635_),
    .Q(\reg_module.gprf[533] ));
 sky130_fd_sc_hd__dfxtp_1 _13020_ (.CLK(clknet_leaf_71_clk),
    .D(_00636_),
    .Q(\reg_module.gprf[534] ));
 sky130_fd_sc_hd__dfxtp_1 _13021_ (.CLK(clknet_leaf_98_clk),
    .D(_00637_),
    .Q(\reg_module.gprf[535] ));
 sky130_fd_sc_hd__dfxtp_1 _13022_ (.CLK(clknet_leaf_81_clk),
    .D(_00638_),
    .Q(\reg_module.gprf[536] ));
 sky130_fd_sc_hd__dfxtp_1 _13023_ (.CLK(clknet_leaf_88_clk),
    .D(_00639_),
    .Q(\reg_module.gprf[537] ));
 sky130_fd_sc_hd__dfxtp_1 _13024_ (.CLK(clknet_leaf_78_clk),
    .D(_00640_),
    .Q(\reg_module.gprf[538] ));
 sky130_fd_sc_hd__dfxtp_1 _13025_ (.CLK(clknet_leaf_98_clk),
    .D(_00641_),
    .Q(\reg_module.gprf[539] ));
 sky130_fd_sc_hd__dfxtp_1 _13026_ (.CLK(clknet_leaf_90_clk),
    .D(_00642_),
    .Q(\reg_module.gprf[540] ));
 sky130_fd_sc_hd__dfxtp_1 _13027_ (.CLK(clknet_leaf_80_clk),
    .D(_00643_),
    .Q(\reg_module.gprf[541] ));
 sky130_fd_sc_hd__dfxtp_1 _13028_ (.CLK(clknet_leaf_69_clk),
    .D(_00644_),
    .Q(\reg_module.gprf[542] ));
 sky130_fd_sc_hd__dfxtp_1 _13029_ (.CLK(clknet_leaf_61_clk),
    .D(_00645_),
    .Q(\reg_module.gprf[543] ));
 sky130_fd_sc_hd__dfxtp_1 _13030_ (.CLK(clknet_leaf_11_clk),
    .D(_00646_),
    .Q(\reg_module.gprf[544] ));
 sky130_fd_sc_hd__dfxtp_1 _13031_ (.CLK(clknet_leaf_34_clk),
    .D(_00647_),
    .Q(\reg_module.gprf[545] ));
 sky130_fd_sc_hd__dfxtp_1 _13032_ (.CLK(clknet_leaf_13_clk),
    .D(_00648_),
    .Q(\reg_module.gprf[546] ));
 sky130_fd_sc_hd__dfxtp_1 _13033_ (.CLK(clknet_leaf_4_clk),
    .D(_00649_),
    .Q(\reg_module.gprf[547] ));
 sky130_fd_sc_hd__dfxtp_1 _13034_ (.CLK(clknet_leaf_32_clk),
    .D(_00650_),
    .Q(\reg_module.gprf[548] ));
 sky130_fd_sc_hd__dfxtp_1 _13035_ (.CLK(clknet_leaf_9_clk),
    .D(_00651_),
    .Q(\reg_module.gprf[549] ));
 sky130_fd_sc_hd__dfxtp_1 _13036_ (.CLK(clknet_leaf_2_clk),
    .D(_00652_),
    .Q(\reg_module.gprf[550] ));
 sky130_fd_sc_hd__dfxtp_1 _13037_ (.CLK(clknet_leaf_4_clk),
    .D(_00653_),
    .Q(\reg_module.gprf[551] ));
 sky130_fd_sc_hd__dfxtp_1 _13038_ (.CLK(clknet_leaf_27_clk),
    .D(_00654_),
    .Q(\reg_module.gprf[552] ));
 sky130_fd_sc_hd__dfxtp_1 _13039_ (.CLK(clknet_leaf_128_clk),
    .D(_00655_),
    .Q(\reg_module.gprf[553] ));
 sky130_fd_sc_hd__dfxtp_1 _13040_ (.CLK(clknet_leaf_2_clk),
    .D(_00656_),
    .Q(\reg_module.gprf[554] ));
 sky130_fd_sc_hd__dfxtp_1 _13041_ (.CLK(clknet_leaf_126_clk),
    .D(_00657_),
    .Q(\reg_module.gprf[555] ));
 sky130_fd_sc_hd__dfxtp_1 _13042_ (.CLK(clknet_leaf_115_clk),
    .D(_00658_),
    .Q(\reg_module.gprf[556] ));
 sky130_fd_sc_hd__dfxtp_1 _13043_ (.CLK(clknet_leaf_117_clk),
    .D(_00659_),
    .Q(\reg_module.gprf[557] ));
 sky130_fd_sc_hd__dfxtp_1 _13044_ (.CLK(clknet_leaf_18_clk),
    .D(_00660_),
    .Q(\reg_module.gprf[558] ));
 sky130_fd_sc_hd__dfxtp_1 _13045_ (.CLK(clknet_leaf_111_clk),
    .D(_00661_),
    .Q(\reg_module.gprf[559] ));
 sky130_fd_sc_hd__dfxtp_1 _13046_ (.CLK(clknet_leaf_53_clk),
    .D(_00662_),
    .Q(\reg_module.gprf[560] ));
 sky130_fd_sc_hd__dfxtp_1 _13047_ (.CLK(clknet_leaf_106_clk),
    .D(_00663_),
    .Q(\reg_module.gprf[561] ));
 sky130_fd_sc_hd__dfxtp_1 _13048_ (.CLK(clknet_leaf_104_clk),
    .D(_00664_),
    .Q(\reg_module.gprf[562] ));
 sky130_fd_sc_hd__dfxtp_1 _13049_ (.CLK(clknet_leaf_105_clk),
    .D(_00665_),
    .Q(\reg_module.gprf[563] ));
 sky130_fd_sc_hd__dfxtp_1 _13050_ (.CLK(clknet_leaf_115_clk),
    .D(_00666_),
    .Q(\reg_module.gprf[564] ));
 sky130_fd_sc_hd__dfxtp_1 _13051_ (.CLK(clknet_leaf_60_clk),
    .D(_00667_),
    .Q(\reg_module.gprf[565] ));
 sky130_fd_sc_hd__dfxtp_1 _13052_ (.CLK(clknet_leaf_70_clk),
    .D(_00668_),
    .Q(\reg_module.gprf[566] ));
 sky130_fd_sc_hd__dfxtp_1 _13053_ (.CLK(clknet_leaf_98_clk),
    .D(_00669_),
    .Q(\reg_module.gprf[567] ));
 sky130_fd_sc_hd__dfxtp_1 _13054_ (.CLK(clknet_leaf_81_clk),
    .D(_00670_),
    .Q(\reg_module.gprf[568] ));
 sky130_fd_sc_hd__dfxtp_1 _13055_ (.CLK(clknet_leaf_89_clk),
    .D(_00671_),
    .Q(\reg_module.gprf[569] ));
 sky130_fd_sc_hd__dfxtp_1 _13056_ (.CLK(clknet_leaf_77_clk),
    .D(_00672_),
    .Q(\reg_module.gprf[570] ));
 sky130_fd_sc_hd__dfxtp_1 _13057_ (.CLK(clknet_leaf_98_clk),
    .D(_00673_),
    .Q(\reg_module.gprf[571] ));
 sky130_fd_sc_hd__dfxtp_1 _13058_ (.CLK(clknet_leaf_90_clk),
    .D(_00674_),
    .Q(\reg_module.gprf[572] ));
 sky130_fd_sc_hd__dfxtp_1 _13059_ (.CLK(clknet_leaf_89_clk),
    .D(_00675_),
    .Q(\reg_module.gprf[573] ));
 sky130_fd_sc_hd__dfxtp_1 _13060_ (.CLK(clknet_leaf_69_clk),
    .D(_00676_),
    .Q(\reg_module.gprf[574] ));
 sky130_fd_sc_hd__dfxtp_1 _13061_ (.CLK(clknet_leaf_61_clk),
    .D(_00677_),
    .Q(\reg_module.gprf[575] ));
 sky130_fd_sc_hd__dfxtp_1 _13062_ (.CLK(clknet_leaf_16_clk),
    .D(_00678_),
    .Q(\reg_module.gprf[576] ));
 sky130_fd_sc_hd__dfxtp_1 _13063_ (.CLK(clknet_leaf_34_clk),
    .D(_00679_),
    .Q(\reg_module.gprf[577] ));
 sky130_fd_sc_hd__dfxtp_1 _13064_ (.CLK(clknet_leaf_13_clk),
    .D(_00680_),
    .Q(\reg_module.gprf[578] ));
 sky130_fd_sc_hd__dfxtp_1 _13065_ (.CLK(clknet_leaf_4_clk),
    .D(_00681_),
    .Q(\reg_module.gprf[579] ));
 sky130_fd_sc_hd__dfxtp_1 _13066_ (.CLK(clknet_leaf_32_clk),
    .D(_00682_),
    .Q(\reg_module.gprf[580] ));
 sky130_fd_sc_hd__dfxtp_1 _13067_ (.CLK(clknet_leaf_9_clk),
    .D(_00683_),
    .Q(\reg_module.gprf[581] ));
 sky130_fd_sc_hd__dfxtp_1 _13068_ (.CLK(clknet_leaf_2_clk),
    .D(_00684_),
    .Q(\reg_module.gprf[582] ));
 sky130_fd_sc_hd__dfxtp_1 _13069_ (.CLK(clknet_leaf_4_clk),
    .D(_00685_),
    .Q(\reg_module.gprf[583] ));
 sky130_fd_sc_hd__dfxtp_1 _13070_ (.CLK(clknet_leaf_25_clk),
    .D(_00686_),
    .Q(\reg_module.gprf[584] ));
 sky130_fd_sc_hd__dfxtp_1 _13071_ (.CLK(clknet_leaf_127_clk),
    .D(_00687_),
    .Q(\reg_module.gprf[585] ));
 sky130_fd_sc_hd__dfxtp_1 _13072_ (.CLK(clknet_leaf_128_clk),
    .D(_00688_),
    .Q(\reg_module.gprf[586] ));
 sky130_fd_sc_hd__dfxtp_1 _13073_ (.CLK(clknet_leaf_118_clk),
    .D(_00689_),
    .Q(\reg_module.gprf[587] ));
 sky130_fd_sc_hd__dfxtp_1 _13074_ (.CLK(clknet_leaf_118_clk),
    .D(_00690_),
    .Q(\reg_module.gprf[588] ));
 sky130_fd_sc_hd__dfxtp_1 _13075_ (.CLK(clknet_leaf_116_clk),
    .D(_00691_),
    .Q(\reg_module.gprf[589] ));
 sky130_fd_sc_hd__dfxtp_1 _13076_ (.CLK(clknet_leaf_18_clk),
    .D(_00692_),
    .Q(\reg_module.gprf[590] ));
 sky130_fd_sc_hd__dfxtp_1 _13077_ (.CLK(clknet_leaf_76_clk),
    .D(_00693_),
    .Q(\reg_module.gprf[591] ));
 sky130_fd_sc_hd__dfxtp_1 _13078_ (.CLK(clknet_leaf_53_clk),
    .D(_00694_),
    .Q(\reg_module.gprf[592] ));
 sky130_fd_sc_hd__dfxtp_1 _13079_ (.CLK(clknet_leaf_106_clk),
    .D(_00695_),
    .Q(\reg_module.gprf[593] ));
 sky130_fd_sc_hd__dfxtp_1 _13080_ (.CLK(clknet_leaf_104_clk),
    .D(_00696_),
    .Q(\reg_module.gprf[594] ));
 sky130_fd_sc_hd__dfxtp_1 _13081_ (.CLK(clknet_leaf_105_clk),
    .D(_00697_),
    .Q(\reg_module.gprf[595] ));
 sky130_fd_sc_hd__dfxtp_1 _13082_ (.CLK(clknet_leaf_113_clk),
    .D(_00698_),
    .Q(\reg_module.gprf[596] ));
 sky130_fd_sc_hd__dfxtp_1 _13083_ (.CLK(clknet_leaf_55_clk),
    .D(_00699_),
    .Q(\reg_module.gprf[597] ));
 sky130_fd_sc_hd__dfxtp_1 _13084_ (.CLK(clknet_leaf_70_clk),
    .D(_00700_),
    .Q(\reg_module.gprf[598] ));
 sky130_fd_sc_hd__dfxtp_1 _13085_ (.CLK(clknet_leaf_98_clk),
    .D(_00701_),
    .Q(\reg_module.gprf[599] ));
 sky130_fd_sc_hd__dfxtp_1 _13086_ (.CLK(clknet_leaf_81_clk),
    .D(_00702_),
    .Q(\reg_module.gprf[600] ));
 sky130_fd_sc_hd__dfxtp_1 _13087_ (.CLK(clknet_leaf_89_clk),
    .D(_00703_),
    .Q(\reg_module.gprf[601] ));
 sky130_fd_sc_hd__dfxtp_1 _13088_ (.CLK(clknet_leaf_77_clk),
    .D(_00704_),
    .Q(\reg_module.gprf[602] ));
 sky130_fd_sc_hd__dfxtp_1 _13089_ (.CLK(clknet_leaf_98_clk),
    .D(_00705_),
    .Q(\reg_module.gprf[603] ));
 sky130_fd_sc_hd__dfxtp_1 _13090_ (.CLK(clknet_leaf_90_clk),
    .D(_00706_),
    .Q(\reg_module.gprf[604] ));
 sky130_fd_sc_hd__dfxtp_1 _13091_ (.CLK(clknet_leaf_89_clk),
    .D(_00707_),
    .Q(\reg_module.gprf[605] ));
 sky130_fd_sc_hd__dfxtp_1 _13092_ (.CLK(clknet_leaf_68_clk),
    .D(_00708_),
    .Q(\reg_module.gprf[606] ));
 sky130_fd_sc_hd__dfxtp_1 _13093_ (.CLK(clknet_leaf_62_clk),
    .D(_00709_),
    .Q(\reg_module.gprf[607] ));
 sky130_fd_sc_hd__dfxtp_1 _13094_ (.CLK(clknet_leaf_16_clk),
    .D(_00710_),
    .Q(\reg_module.gprf[608] ));
 sky130_fd_sc_hd__dfxtp_1 _13095_ (.CLK(clknet_leaf_34_clk),
    .D(_00711_),
    .Q(\reg_module.gprf[609] ));
 sky130_fd_sc_hd__dfxtp_1 _13096_ (.CLK(clknet_leaf_13_clk),
    .D(_00712_),
    .Q(\reg_module.gprf[610] ));
 sky130_fd_sc_hd__dfxtp_1 _13097_ (.CLK(clknet_leaf_4_clk),
    .D(_00713_),
    .Q(\reg_module.gprf[611] ));
 sky130_fd_sc_hd__dfxtp_1 _13098_ (.CLK(clknet_leaf_32_clk),
    .D(_00714_),
    .Q(\reg_module.gprf[612] ));
 sky130_fd_sc_hd__dfxtp_1 _13099_ (.CLK(clknet_leaf_10_clk),
    .D(_00715_),
    .Q(\reg_module.gprf[613] ));
 sky130_fd_sc_hd__dfxtp_1 _13100_ (.CLK(clknet_leaf_2_clk),
    .D(_00716_),
    .Q(\reg_module.gprf[614] ));
 sky130_fd_sc_hd__dfxtp_1 _13101_ (.CLK(clknet_leaf_12_clk),
    .D(_00717_),
    .Q(\reg_module.gprf[615] ));
 sky130_fd_sc_hd__dfxtp_1 _13102_ (.CLK(clknet_leaf_26_clk),
    .D(_00718_),
    .Q(\reg_module.gprf[616] ));
 sky130_fd_sc_hd__dfxtp_1 _13103_ (.CLK(clknet_leaf_126_clk),
    .D(_00719_),
    .Q(\reg_module.gprf[617] ));
 sky130_fd_sc_hd__dfxtp_1 _13104_ (.CLK(clknet_leaf_128_clk),
    .D(_00720_),
    .Q(\reg_module.gprf[618] ));
 sky130_fd_sc_hd__dfxtp_1 _13105_ (.CLK(clknet_leaf_118_clk),
    .D(_00721_),
    .Q(\reg_module.gprf[619] ));
 sky130_fd_sc_hd__dfxtp_1 _13106_ (.CLK(clknet_leaf_118_clk),
    .D(_00722_),
    .Q(\reg_module.gprf[620] ));
 sky130_fd_sc_hd__dfxtp_1 _13107_ (.CLK(clknet_leaf_117_clk),
    .D(_00723_),
    .Q(\reg_module.gprf[621] ));
 sky130_fd_sc_hd__dfxtp_1 _13108_ (.CLK(clknet_leaf_112_clk),
    .D(_00724_),
    .Q(\reg_module.gprf[622] ));
 sky130_fd_sc_hd__dfxtp_1 _13109_ (.CLK(clknet_leaf_76_clk),
    .D(_00725_),
    .Q(\reg_module.gprf[623] ));
 sky130_fd_sc_hd__dfxtp_1 _13110_ (.CLK(clknet_leaf_54_clk),
    .D(_00726_),
    .Q(\reg_module.gprf[624] ));
 sky130_fd_sc_hd__dfxtp_1 _13111_ (.CLK(clknet_leaf_106_clk),
    .D(_00727_),
    .Q(\reg_module.gprf[625] ));
 sky130_fd_sc_hd__dfxtp_1 _13112_ (.CLK(clknet_leaf_104_clk),
    .D(_00728_),
    .Q(\reg_module.gprf[626] ));
 sky130_fd_sc_hd__dfxtp_1 _13113_ (.CLK(clknet_leaf_105_clk),
    .D(_00729_),
    .Q(\reg_module.gprf[627] ));
 sky130_fd_sc_hd__dfxtp_1 _13114_ (.CLK(clknet_leaf_115_clk),
    .D(_00730_),
    .Q(\reg_module.gprf[628] ));
 sky130_fd_sc_hd__dfxtp_1 _13115_ (.CLK(clknet_leaf_60_clk),
    .D(_00731_),
    .Q(\reg_module.gprf[629] ));
 sky130_fd_sc_hd__dfxtp_1 _13116_ (.CLK(clknet_leaf_65_clk),
    .D(_00732_),
    .Q(\reg_module.gprf[630] ));
 sky130_fd_sc_hd__dfxtp_1 _13117_ (.CLK(clknet_leaf_89_clk),
    .D(_00733_),
    .Q(\reg_module.gprf[631] ));
 sky130_fd_sc_hd__dfxtp_1 _13118_ (.CLK(clknet_leaf_88_clk),
    .D(_00734_),
    .Q(\reg_module.gprf[632] ));
 sky130_fd_sc_hd__dfxtp_1 _13119_ (.CLK(clknet_leaf_88_clk),
    .D(_00735_),
    .Q(\reg_module.gprf[633] ));
 sky130_fd_sc_hd__dfxtp_1 _13120_ (.CLK(clknet_leaf_78_clk),
    .D(_00736_),
    .Q(\reg_module.gprf[634] ));
 sky130_fd_sc_hd__dfxtp_1 _13121_ (.CLK(clknet_leaf_97_clk),
    .D(_00737_),
    .Q(\reg_module.gprf[635] ));
 sky130_fd_sc_hd__dfxtp_1 _13122_ (.CLK(clknet_leaf_90_clk),
    .D(_00738_),
    .Q(\reg_module.gprf[636] ));
 sky130_fd_sc_hd__dfxtp_1 _13123_ (.CLK(clknet_leaf_89_clk),
    .D(_00739_),
    .Q(\reg_module.gprf[637] ));
 sky130_fd_sc_hd__dfxtp_1 _13124_ (.CLK(clknet_leaf_83_clk),
    .D(_00740_),
    .Q(\reg_module.gprf[638] ));
 sky130_fd_sc_hd__dfxtp_1 _13125_ (.CLK(clknet_leaf_61_clk),
    .D(_00741_),
    .Q(\reg_module.gprf[639] ));
 sky130_fd_sc_hd__dfxtp_1 _13126_ (.CLK(clknet_leaf_11_clk),
    .D(_00742_),
    .Q(\reg_module.gprf[640] ));
 sky130_fd_sc_hd__dfxtp_1 _13127_ (.CLK(clknet_leaf_34_clk),
    .D(_00743_),
    .Q(\reg_module.gprf[641] ));
 sky130_fd_sc_hd__dfxtp_1 _13128_ (.CLK(clknet_leaf_13_clk),
    .D(_00744_),
    .Q(\reg_module.gprf[642] ));
 sky130_fd_sc_hd__dfxtp_1 _13129_ (.CLK(clknet_leaf_4_clk),
    .D(_00745_),
    .Q(\reg_module.gprf[643] ));
 sky130_fd_sc_hd__dfxtp_1 _13130_ (.CLK(clknet_leaf_31_clk),
    .D(_00746_),
    .Q(\reg_module.gprf[644] ));
 sky130_fd_sc_hd__dfxtp_1 _13131_ (.CLK(clknet_leaf_8_clk),
    .D(_00747_),
    .Q(\reg_module.gprf[645] ));
 sky130_fd_sc_hd__dfxtp_1 _13132_ (.CLK(clknet_leaf_1_clk),
    .D(_00748_),
    .Q(\reg_module.gprf[646] ));
 sky130_fd_sc_hd__dfxtp_1 _13133_ (.CLK(clknet_leaf_6_clk),
    .D(_00749_),
    .Q(\reg_module.gprf[647] ));
 sky130_fd_sc_hd__dfxtp_1 _13134_ (.CLK(clknet_leaf_27_clk),
    .D(_00750_),
    .Q(\reg_module.gprf[648] ));
 sky130_fd_sc_hd__dfxtp_1 _13135_ (.CLK(clknet_leaf_128_clk),
    .D(_00751_),
    .Q(\reg_module.gprf[649] ));
 sky130_fd_sc_hd__dfxtp_1 _13136_ (.CLK(clknet_leaf_2_clk),
    .D(_00752_),
    .Q(\reg_module.gprf[650] ));
 sky130_fd_sc_hd__dfxtp_1 _13137_ (.CLK(clknet_leaf_125_clk),
    .D(_00753_),
    .Q(\reg_module.gprf[651] ));
 sky130_fd_sc_hd__dfxtp_1 _13138_ (.CLK(clknet_leaf_118_clk),
    .D(_00754_),
    .Q(\reg_module.gprf[652] ));
 sky130_fd_sc_hd__dfxtp_1 _13139_ (.CLK(clknet_leaf_118_clk),
    .D(_00755_),
    .Q(\reg_module.gprf[653] ));
 sky130_fd_sc_hd__dfxtp_1 _13140_ (.CLK(clknet_leaf_17_clk),
    .D(_00756_),
    .Q(\reg_module.gprf[654] ));
 sky130_fd_sc_hd__dfxtp_1 _13141_ (.CLK(clknet_leaf_111_clk),
    .D(_00757_),
    .Q(\reg_module.gprf[655] ));
 sky130_fd_sc_hd__dfxtp_1 _13142_ (.CLK(clknet_leaf_61_clk),
    .D(_00758_),
    .Q(\reg_module.gprf[656] ));
 sky130_fd_sc_hd__dfxtp_1 _13143_ (.CLK(clknet_leaf_99_clk),
    .D(_00759_),
    .Q(\reg_module.gprf[657] ));
 sky130_fd_sc_hd__dfxtp_1 _13144_ (.CLK(clknet_leaf_119_clk),
    .D(_00760_),
    .Q(\reg_module.gprf[658] ));
 sky130_fd_sc_hd__dfxtp_1 _13145_ (.CLK(clknet_leaf_106_clk),
    .D(_00761_),
    .Q(\reg_module.gprf[659] ));
 sky130_fd_sc_hd__dfxtp_1 _13146_ (.CLK(clknet_leaf_15_clk),
    .D(_00762_),
    .Q(\reg_module.gprf[660] ));
 sky130_fd_sc_hd__dfxtp_1 _13147_ (.CLK(clknet_leaf_60_clk),
    .D(_00763_),
    .Q(\reg_module.gprf[661] ));
 sky130_fd_sc_hd__dfxtp_1 _13148_ (.CLK(clknet_leaf_68_clk),
    .D(_00764_),
    .Q(\reg_module.gprf[662] ));
 sky130_fd_sc_hd__dfxtp_1 _13149_ (.CLK(clknet_leaf_97_clk),
    .D(_00765_),
    .Q(\reg_module.gprf[663] ));
 sky130_fd_sc_hd__dfxtp_1 _13150_ (.CLK(clknet_leaf_88_clk),
    .D(_00766_),
    .Q(\reg_module.gprf[664] ));
 sky130_fd_sc_hd__dfxtp_1 _13151_ (.CLK(clknet_leaf_89_clk),
    .D(_00767_),
    .Q(\reg_module.gprf[665] ));
 sky130_fd_sc_hd__dfxtp_1 _13152_ (.CLK(clknet_leaf_77_clk),
    .D(_00768_),
    .Q(\reg_module.gprf[666] ));
 sky130_fd_sc_hd__dfxtp_1 _13153_ (.CLK(clknet_leaf_99_clk),
    .D(_00769_),
    .Q(\reg_module.gprf[667] ));
 sky130_fd_sc_hd__dfxtp_1 _13154_ (.CLK(clknet_leaf_97_clk),
    .D(_00770_),
    .Q(\reg_module.gprf[668] ));
 sky130_fd_sc_hd__dfxtp_1 _13155_ (.CLK(clknet_leaf_89_clk),
    .D(_00771_),
    .Q(\reg_module.gprf[669] ));
 sky130_fd_sc_hd__dfxtp_1 _13156_ (.CLK(clknet_leaf_83_clk),
    .D(_00772_),
    .Q(\reg_module.gprf[670] ));
 sky130_fd_sc_hd__dfxtp_1 _13157_ (.CLK(clknet_leaf_62_clk),
    .D(_00773_),
    .Q(\reg_module.gprf[671] ));
 sky130_fd_sc_hd__dfxtp_1 _13158_ (.CLK(clknet_leaf_11_clk),
    .D(_00774_),
    .Q(\reg_module.gprf[672] ));
 sky130_fd_sc_hd__dfxtp_1 _13159_ (.CLK(clknet_leaf_34_clk),
    .D(_00775_),
    .Q(\reg_module.gprf[673] ));
 sky130_fd_sc_hd__dfxtp_1 _13160_ (.CLK(clknet_leaf_13_clk),
    .D(_00776_),
    .Q(\reg_module.gprf[674] ));
 sky130_fd_sc_hd__dfxtp_1 _13161_ (.CLK(clknet_leaf_4_clk),
    .D(_00777_),
    .Q(\reg_module.gprf[675] ));
 sky130_fd_sc_hd__dfxtp_1 _13162_ (.CLK(clknet_leaf_31_clk),
    .D(_00778_),
    .Q(\reg_module.gprf[676] ));
 sky130_fd_sc_hd__dfxtp_1 _13163_ (.CLK(clknet_leaf_8_clk),
    .D(_00779_),
    .Q(\reg_module.gprf[677] ));
 sky130_fd_sc_hd__dfxtp_1 _13164_ (.CLK(clknet_leaf_1_clk),
    .D(_00780_),
    .Q(\reg_module.gprf[678] ));
 sky130_fd_sc_hd__dfxtp_1 _13165_ (.CLK(clknet_leaf_6_clk),
    .D(_00781_),
    .Q(\reg_module.gprf[679] ));
 sky130_fd_sc_hd__dfxtp_1 _13166_ (.CLK(clknet_leaf_27_clk),
    .D(_00782_),
    .Q(\reg_module.gprf[680] ));
 sky130_fd_sc_hd__dfxtp_1 _13167_ (.CLK(clknet_leaf_128_clk),
    .D(_00783_),
    .Q(\reg_module.gprf[681] ));
 sky130_fd_sc_hd__dfxtp_1 _13168_ (.CLK(clknet_leaf_2_clk),
    .D(_00784_),
    .Q(\reg_module.gprf[682] ));
 sky130_fd_sc_hd__dfxtp_1 _13169_ (.CLK(clknet_leaf_125_clk),
    .D(_00785_),
    .Q(\reg_module.gprf[683] ));
 sky130_fd_sc_hd__dfxtp_1 _13170_ (.CLK(clknet_leaf_118_clk),
    .D(_00786_),
    .Q(\reg_module.gprf[684] ));
 sky130_fd_sc_hd__dfxtp_1 _13171_ (.CLK(clknet_leaf_117_clk),
    .D(_00787_),
    .Q(\reg_module.gprf[685] ));
 sky130_fd_sc_hd__dfxtp_1 _13172_ (.CLK(clknet_leaf_17_clk),
    .D(_00788_),
    .Q(\reg_module.gprf[686] ));
 sky130_fd_sc_hd__dfxtp_1 _13173_ (.CLK(clknet_leaf_111_clk),
    .D(_00789_),
    .Q(\reg_module.gprf[687] ));
 sky130_fd_sc_hd__dfxtp_1 _13174_ (.CLK(clknet_leaf_54_clk),
    .D(_00790_),
    .Q(\reg_module.gprf[688] ));
 sky130_fd_sc_hd__dfxtp_1 _13175_ (.CLK(clknet_leaf_101_clk),
    .D(_00791_),
    .Q(\reg_module.gprf[689] ));
 sky130_fd_sc_hd__dfxtp_1 _13176_ (.CLK(clknet_leaf_119_clk),
    .D(_00792_),
    .Q(\reg_module.gprf[690] ));
 sky130_fd_sc_hd__dfxtp_1 _13177_ (.CLK(clknet_leaf_106_clk),
    .D(_00793_),
    .Q(\reg_module.gprf[691] ));
 sky130_fd_sc_hd__dfxtp_1 _13178_ (.CLK(clknet_leaf_116_clk),
    .D(_00794_),
    .Q(\reg_module.gprf[692] ));
 sky130_fd_sc_hd__dfxtp_1 _13179_ (.CLK(clknet_leaf_61_clk),
    .D(_00795_),
    .Q(\reg_module.gprf[693] ));
 sky130_fd_sc_hd__dfxtp_1 _13180_ (.CLK(clknet_leaf_70_clk),
    .D(_00796_),
    .Q(\reg_module.gprf[694] ));
 sky130_fd_sc_hd__dfxtp_1 _13181_ (.CLK(clknet_leaf_97_clk),
    .D(_00797_),
    .Q(\reg_module.gprf[695] ));
 sky130_fd_sc_hd__dfxtp_1 _13182_ (.CLK(clknet_leaf_88_clk),
    .D(_00798_),
    .Q(\reg_module.gprf[696] ));
 sky130_fd_sc_hd__dfxtp_1 _13183_ (.CLK(clknet_leaf_89_clk),
    .D(_00799_),
    .Q(\reg_module.gprf[697] ));
 sky130_fd_sc_hd__dfxtp_1 _13184_ (.CLK(clknet_leaf_77_clk),
    .D(_00800_),
    .Q(\reg_module.gprf[698] ));
 sky130_fd_sc_hd__dfxtp_1 _13185_ (.CLK(clknet_leaf_99_clk),
    .D(_00801_),
    .Q(\reg_module.gprf[699] ));
 sky130_fd_sc_hd__dfxtp_1 _13186_ (.CLK(clknet_leaf_97_clk),
    .D(_00802_),
    .Q(\reg_module.gprf[700] ));
 sky130_fd_sc_hd__dfxtp_1 _13187_ (.CLK(clknet_leaf_98_clk),
    .D(_00803_),
    .Q(\reg_module.gprf[701] ));
 sky130_fd_sc_hd__dfxtp_1 _13188_ (.CLK(clknet_leaf_83_clk),
    .D(_00804_),
    .Q(\reg_module.gprf[702] ));
 sky130_fd_sc_hd__dfxtp_1 _13189_ (.CLK(clknet_leaf_62_clk),
    .D(_00805_),
    .Q(\reg_module.gprf[703] ));
 sky130_fd_sc_hd__dfxtp_1 _13190_ (.CLK(clknet_leaf_12_clk),
    .D(_00806_),
    .Q(\reg_module.gprf[704] ));
 sky130_fd_sc_hd__dfxtp_1 _13191_ (.CLK(clknet_leaf_34_clk),
    .D(_00807_),
    .Q(\reg_module.gprf[705] ));
 sky130_fd_sc_hd__dfxtp_1 _13192_ (.CLK(clknet_leaf_14_clk),
    .D(_00808_),
    .Q(\reg_module.gprf[706] ));
 sky130_fd_sc_hd__dfxtp_1 _13193_ (.CLK(clknet_leaf_3_clk),
    .D(_00809_),
    .Q(\reg_module.gprf[707] ));
 sky130_fd_sc_hd__dfxtp_1 _13194_ (.CLK(clknet_leaf_31_clk),
    .D(_00810_),
    .Q(\reg_module.gprf[708] ));
 sky130_fd_sc_hd__dfxtp_1 _13195_ (.CLK(clknet_leaf_9_clk),
    .D(_00811_),
    .Q(\reg_module.gprf[709] ));
 sky130_fd_sc_hd__dfxtp_1 _13196_ (.CLK(clknet_leaf_2_clk),
    .D(_00812_),
    .Q(\reg_module.gprf[710] ));
 sky130_fd_sc_hd__dfxtp_1 _13197_ (.CLK(clknet_leaf_6_clk),
    .D(_00813_),
    .Q(\reg_module.gprf[711] ));
 sky130_fd_sc_hd__dfxtp_1 _13198_ (.CLK(clknet_leaf_27_clk),
    .D(_00814_),
    .Q(\reg_module.gprf[712] ));
 sky130_fd_sc_hd__dfxtp_1 _13199_ (.CLK(clknet_leaf_128_clk),
    .D(_00815_),
    .Q(\reg_module.gprf[713] ));
 sky130_fd_sc_hd__dfxtp_1 _13200_ (.CLK(clknet_leaf_2_clk),
    .D(_00816_),
    .Q(\reg_module.gprf[714] ));
 sky130_fd_sc_hd__dfxtp_1 _13201_ (.CLK(clknet_leaf_123_clk),
    .D(_00817_),
    .Q(\reg_module.gprf[715] ));
 sky130_fd_sc_hd__dfxtp_1 _13202_ (.CLK(clknet_leaf_118_clk),
    .D(_00818_),
    .Q(\reg_module.gprf[716] ));
 sky130_fd_sc_hd__dfxtp_1 _13203_ (.CLK(clknet_leaf_118_clk),
    .D(_00819_),
    .Q(\reg_module.gprf[717] ));
 sky130_fd_sc_hd__dfxtp_1 _13204_ (.CLK(clknet_leaf_18_clk),
    .D(_00820_),
    .Q(\reg_module.gprf[718] ));
 sky130_fd_sc_hd__dfxtp_1 _13205_ (.CLK(clknet_leaf_111_clk),
    .D(_00821_),
    .Q(\reg_module.gprf[719] ));
 sky130_fd_sc_hd__dfxtp_1 _13206_ (.CLK(clknet_leaf_61_clk),
    .D(_00822_),
    .Q(\reg_module.gprf[720] ));
 sky130_fd_sc_hd__dfxtp_1 _13207_ (.CLK(clknet_leaf_103_clk),
    .D(_00823_),
    .Q(\reg_module.gprf[721] ));
 sky130_fd_sc_hd__dfxtp_1 _13208_ (.CLK(clknet_leaf_119_clk),
    .D(_00824_),
    .Q(\reg_module.gprf[722] ));
 sky130_fd_sc_hd__dfxtp_1 _13209_ (.CLK(clknet_leaf_106_clk),
    .D(_00825_),
    .Q(\reg_module.gprf[723] ));
 sky130_fd_sc_hd__dfxtp_1 _13210_ (.CLK(clknet_leaf_116_clk),
    .D(_00826_),
    .Q(\reg_module.gprf[724] ));
 sky130_fd_sc_hd__dfxtp_1 _13211_ (.CLK(clknet_leaf_60_clk),
    .D(_00827_),
    .Q(\reg_module.gprf[725] ));
 sky130_fd_sc_hd__dfxtp_1 _13212_ (.CLK(clknet_leaf_68_clk),
    .D(_00828_),
    .Q(\reg_module.gprf[726] ));
 sky130_fd_sc_hd__dfxtp_1 _13213_ (.CLK(clknet_leaf_90_clk),
    .D(_00829_),
    .Q(\reg_module.gprf[727] ));
 sky130_fd_sc_hd__dfxtp_1 _13214_ (.CLK(clknet_leaf_88_clk),
    .D(_00830_),
    .Q(\reg_module.gprf[728] ));
 sky130_fd_sc_hd__dfxtp_1 _13215_ (.CLK(clknet_leaf_90_clk),
    .D(_00831_),
    .Q(\reg_module.gprf[729] ));
 sky130_fd_sc_hd__dfxtp_1 _13216_ (.CLK(clknet_leaf_77_clk),
    .D(_00832_),
    .Q(\reg_module.gprf[730] ));
 sky130_fd_sc_hd__dfxtp_1 _13217_ (.CLK(clknet_leaf_99_clk),
    .D(_00833_),
    .Q(\reg_module.gprf[731] ));
 sky130_fd_sc_hd__dfxtp_1 _13218_ (.CLK(clknet_leaf_90_clk),
    .D(_00834_),
    .Q(\reg_module.gprf[732] ));
 sky130_fd_sc_hd__dfxtp_1 _13219_ (.CLK(clknet_leaf_89_clk),
    .D(_00835_),
    .Q(\reg_module.gprf[733] ));
 sky130_fd_sc_hd__dfxtp_1 _13220_ (.CLK(clknet_leaf_83_clk),
    .D(_00836_),
    .Q(\reg_module.gprf[734] ));
 sky130_fd_sc_hd__dfxtp_1 _13221_ (.CLK(clknet_leaf_62_clk),
    .D(_00837_),
    .Q(\reg_module.gprf[735] ));
 sky130_fd_sc_hd__dfxtp_1 _13222_ (.CLK(clknet_leaf_16_clk),
    .D(_00838_),
    .Q(\reg_module.gprf[736] ));
 sky130_fd_sc_hd__dfxtp_1 _13223_ (.CLK(clknet_leaf_34_clk),
    .D(_00839_),
    .Q(\reg_module.gprf[737] ));
 sky130_fd_sc_hd__dfxtp_1 _13224_ (.CLK(clknet_leaf_14_clk),
    .D(_00840_),
    .Q(\reg_module.gprf[738] ));
 sky130_fd_sc_hd__dfxtp_1 _13225_ (.CLK(clknet_leaf_3_clk),
    .D(_00841_),
    .Q(\reg_module.gprf[739] ));
 sky130_fd_sc_hd__dfxtp_1 _13226_ (.CLK(clknet_leaf_32_clk),
    .D(_00842_),
    .Q(\reg_module.gprf[740] ));
 sky130_fd_sc_hd__dfxtp_1 _13227_ (.CLK(clknet_leaf_9_clk),
    .D(_00843_),
    .Q(\reg_module.gprf[741] ));
 sky130_fd_sc_hd__dfxtp_1 _13228_ (.CLK(clknet_leaf_2_clk),
    .D(_00844_),
    .Q(\reg_module.gprf[742] ));
 sky130_fd_sc_hd__dfxtp_1 _13229_ (.CLK(clknet_leaf_7_clk),
    .D(_00845_),
    .Q(\reg_module.gprf[743] ));
 sky130_fd_sc_hd__dfxtp_1 _13230_ (.CLK(clknet_leaf_26_clk),
    .D(_00846_),
    .Q(\reg_module.gprf[744] ));
 sky130_fd_sc_hd__dfxtp_1 _13231_ (.CLK(clknet_leaf_128_clk),
    .D(_00847_),
    .Q(\reg_module.gprf[745] ));
 sky130_fd_sc_hd__dfxtp_1 _13232_ (.CLK(clknet_leaf_2_clk),
    .D(_00848_),
    .Q(\reg_module.gprf[746] ));
 sky130_fd_sc_hd__dfxtp_1 _13233_ (.CLK(clknet_leaf_123_clk),
    .D(_00849_),
    .Q(\reg_module.gprf[747] ));
 sky130_fd_sc_hd__dfxtp_1 _13234_ (.CLK(clknet_leaf_118_clk),
    .D(_00850_),
    .Q(\reg_module.gprf[748] ));
 sky130_fd_sc_hd__dfxtp_1 _13235_ (.CLK(clknet_leaf_118_clk),
    .D(_00851_),
    .Q(\reg_module.gprf[749] ));
 sky130_fd_sc_hd__dfxtp_1 _13236_ (.CLK(clknet_leaf_18_clk),
    .D(_00852_),
    .Q(\reg_module.gprf[750] ));
 sky130_fd_sc_hd__dfxtp_1 _13237_ (.CLK(clknet_leaf_77_clk),
    .D(_00853_),
    .Q(\reg_module.gprf[751] ));
 sky130_fd_sc_hd__dfxtp_1 _13238_ (.CLK(clknet_leaf_61_clk),
    .D(_00854_),
    .Q(\reg_module.gprf[752] ));
 sky130_fd_sc_hd__dfxtp_1 _13239_ (.CLK(clknet_leaf_101_clk),
    .D(_00855_),
    .Q(\reg_module.gprf[753] ));
 sky130_fd_sc_hd__dfxtp_1 _13240_ (.CLK(clknet_leaf_104_clk),
    .D(_00856_),
    .Q(\reg_module.gprf[754] ));
 sky130_fd_sc_hd__dfxtp_1 _13241_ (.CLK(clknet_leaf_106_clk),
    .D(_00857_),
    .Q(\reg_module.gprf[755] ));
 sky130_fd_sc_hd__dfxtp_1 _13242_ (.CLK(clknet_leaf_113_clk),
    .D(_00858_),
    .Q(\reg_module.gprf[756] ));
 sky130_fd_sc_hd__dfxtp_1 _13243_ (.CLK(clknet_leaf_60_clk),
    .D(_00859_),
    .Q(\reg_module.gprf[757] ));
 sky130_fd_sc_hd__dfxtp_1 _13244_ (.CLK(clknet_leaf_68_clk),
    .D(_00860_),
    .Q(\reg_module.gprf[758] ));
 sky130_fd_sc_hd__dfxtp_1 _13245_ (.CLK(clknet_leaf_90_clk),
    .D(_00861_),
    .Q(\reg_module.gprf[759] ));
 sky130_fd_sc_hd__dfxtp_1 _13246_ (.CLK(clknet_leaf_88_clk),
    .D(_00862_),
    .Q(\reg_module.gprf[760] ));
 sky130_fd_sc_hd__dfxtp_1 _13247_ (.CLK(clknet_leaf_90_clk),
    .D(_00863_),
    .Q(\reg_module.gprf[761] ));
 sky130_fd_sc_hd__dfxtp_1 _13248_ (.CLK(clknet_leaf_78_clk),
    .D(_00864_),
    .Q(\reg_module.gprf[762] ));
 sky130_fd_sc_hd__dfxtp_1 _13249_ (.CLK(clknet_leaf_99_clk),
    .D(_00865_),
    .Q(\reg_module.gprf[763] ));
 sky130_fd_sc_hd__dfxtp_1 _13250_ (.CLK(clknet_leaf_94_clk),
    .D(_00866_),
    .Q(\reg_module.gprf[764] ));
 sky130_fd_sc_hd__dfxtp_1 _13251_ (.CLK(clknet_leaf_89_clk),
    .D(_00867_),
    .Q(\reg_module.gprf[765] ));
 sky130_fd_sc_hd__dfxtp_1 _13252_ (.CLK(clknet_leaf_83_clk),
    .D(_00868_),
    .Q(\reg_module.gprf[766] ));
 sky130_fd_sc_hd__dfxtp_1 _13253_ (.CLK(clknet_leaf_62_clk),
    .D(_00869_),
    .Q(\reg_module.gprf[767] ));
 sky130_fd_sc_hd__dfxtp_1 _13254_ (.CLK(clknet_leaf_25_clk),
    .D(_00870_),
    .Q(\reg_module.gprf[768] ));
 sky130_fd_sc_hd__dfxtp_1 _13255_ (.CLK(clknet_leaf_37_clk),
    .D(_00871_),
    .Q(\reg_module.gprf[769] ));
 sky130_fd_sc_hd__dfxtp_1 _13256_ (.CLK(clknet_leaf_14_clk),
    .D(_00872_),
    .Q(\reg_module.gprf[770] ));
 sky130_fd_sc_hd__dfxtp_1 _13257_ (.CLK(clknet_leaf_4_clk),
    .D(_00873_),
    .Q(\reg_module.gprf[771] ));
 sky130_fd_sc_hd__dfxtp_1 _13258_ (.CLK(clknet_leaf_36_clk),
    .D(_00874_),
    .Q(\reg_module.gprf[772] ));
 sky130_fd_sc_hd__dfxtp_1 _13259_ (.CLK(clknet_leaf_28_clk),
    .D(_00875_),
    .Q(\reg_module.gprf[773] ));
 sky130_fd_sc_hd__dfxtp_1 _13260_ (.CLK(clknet_leaf_5_clk),
    .D(_00876_),
    .Q(\reg_module.gprf[774] ));
 sky130_fd_sc_hd__dfxtp_1 _13261_ (.CLK(clknet_leaf_8_clk),
    .D(_00877_),
    .Q(\reg_module.gprf[775] ));
 sky130_fd_sc_hd__dfxtp_1 _13262_ (.CLK(clknet_leaf_30_clk),
    .D(_00878_),
    .Q(\reg_module.gprf[776] ));
 sky130_fd_sc_hd__dfxtp_1 _13263_ (.CLK(clknet_leaf_129_clk),
    .D(_00879_),
    .Q(\reg_module.gprf[777] ));
 sky130_fd_sc_hd__dfxtp_1 _13264_ (.CLK(clknet_leaf_131_clk),
    .D(_00880_),
    .Q(\reg_module.gprf[778] ));
 sky130_fd_sc_hd__dfxtp_1 _13265_ (.CLK(clknet_leaf_124_clk),
    .D(_00881_),
    .Q(\reg_module.gprf[779] ));
 sky130_fd_sc_hd__dfxtp_1 _13266_ (.CLK(clknet_leaf_105_clk),
    .D(_00882_),
    .Q(\reg_module.gprf[780] ));
 sky130_fd_sc_hd__dfxtp_1 _13267_ (.CLK(clknet_leaf_3_clk),
    .D(_00883_),
    .Q(\reg_module.gprf[781] ));
 sky130_fd_sc_hd__dfxtp_1 _13268_ (.CLK(clknet_leaf_112_clk),
    .D(_00884_),
    .Q(\reg_module.gprf[782] ));
 sky130_fd_sc_hd__dfxtp_1 _13269_ (.CLK(clknet_leaf_109_clk),
    .D(_00885_),
    .Q(\reg_module.gprf[783] ));
 sky130_fd_sc_hd__dfxtp_1 _13270_ (.CLK(clknet_leaf_56_clk),
    .D(_00886_),
    .Q(\reg_module.gprf[784] ));
 sky130_fd_sc_hd__dfxtp_1 _13271_ (.CLK(clknet_leaf_101_clk),
    .D(_00887_),
    .Q(\reg_module.gprf[785] ));
 sky130_fd_sc_hd__dfxtp_1 _13272_ (.CLK(clknet_leaf_121_clk),
    .D(_00888_),
    .Q(\reg_module.gprf[786] ));
 sky130_fd_sc_hd__dfxtp_1 _13273_ (.CLK(clknet_leaf_108_clk),
    .D(_00889_),
    .Q(\reg_module.gprf[787] ));
 sky130_fd_sc_hd__dfxtp_1 _13274_ (.CLK(clknet_leaf_113_clk),
    .D(_00890_),
    .Q(\reg_module.gprf[788] ));
 sky130_fd_sc_hd__dfxtp_1 _13275_ (.CLK(clknet_leaf_57_clk),
    .D(_00891_),
    .Q(\reg_module.gprf[789] ));
 sky130_fd_sc_hd__dfxtp_1 _13276_ (.CLK(clknet_leaf_64_clk),
    .D(_00892_),
    .Q(\reg_module.gprf[790] ));
 sky130_fd_sc_hd__dfxtp_1 _13277_ (.CLK(clknet_leaf_95_clk),
    .D(_00893_),
    .Q(\reg_module.gprf[791] ));
 sky130_fd_sc_hd__dfxtp_1 _13278_ (.CLK(clknet_leaf_85_clk),
    .D(_00894_),
    .Q(\reg_module.gprf[792] ));
 sky130_fd_sc_hd__dfxtp_1 _13279_ (.CLK(clknet_leaf_91_clk),
    .D(_00895_),
    .Q(\reg_module.gprf[793] ));
 sky130_fd_sc_hd__dfxtp_1 _13280_ (.CLK(clknet_leaf_78_clk),
    .D(_00896_),
    .Q(\reg_module.gprf[794] ));
 sky130_fd_sc_hd__dfxtp_1 _13281_ (.CLK(clknet_leaf_100_clk),
    .D(_00897_),
    .Q(\reg_module.gprf[795] ));
 sky130_fd_sc_hd__dfxtp_1 _13282_ (.CLK(clknet_leaf_93_clk),
    .D(_00898_),
    .Q(\reg_module.gprf[796] ));
 sky130_fd_sc_hd__dfxtp_1 _13283_ (.CLK(clknet_leaf_81_clk),
    .D(_00899_),
    .Q(\reg_module.gprf[797] ));
 sky130_fd_sc_hd__dfxtp_1 _13284_ (.CLK(clknet_leaf_83_clk),
    .D(_00900_),
    .Q(\reg_module.gprf[798] ));
 sky130_fd_sc_hd__dfxtp_1 _13285_ (.CLK(clknet_leaf_63_clk),
    .D(_00901_),
    .Q(\reg_module.gprf[799] ));
 sky130_fd_sc_hd__dfxtp_1 _13286_ (.CLK(clknet_leaf_26_clk),
    .D(_00902_),
    .Q(\reg_module.gprf[800] ));
 sky130_fd_sc_hd__dfxtp_1 _13287_ (.CLK(clknet_leaf_37_clk),
    .D(_00903_),
    .Q(\reg_module.gprf[801] ));
 sky130_fd_sc_hd__dfxtp_1 _13288_ (.CLK(clknet_leaf_14_clk),
    .D(_00904_),
    .Q(\reg_module.gprf[802] ));
 sky130_fd_sc_hd__dfxtp_1 _13289_ (.CLK(clknet_leaf_3_clk),
    .D(_00905_),
    .Q(\reg_module.gprf[803] ));
 sky130_fd_sc_hd__dfxtp_1 _13290_ (.CLK(clknet_leaf_36_clk),
    .D(_00906_),
    .Q(\reg_module.gprf[804] ));
 sky130_fd_sc_hd__dfxtp_1 _13291_ (.CLK(clknet_leaf_28_clk),
    .D(_00907_),
    .Q(\reg_module.gprf[805] ));
 sky130_fd_sc_hd__dfxtp_1 _13292_ (.CLK(clknet_leaf_1_clk),
    .D(_00908_),
    .Q(\reg_module.gprf[806] ));
 sky130_fd_sc_hd__dfxtp_1 _13293_ (.CLK(clknet_leaf_8_clk),
    .D(_00909_),
    .Q(\reg_module.gprf[807] ));
 sky130_fd_sc_hd__dfxtp_1 _13294_ (.CLK(clknet_leaf_30_clk),
    .D(_00910_),
    .Q(\reg_module.gprf[808] ));
 sky130_fd_sc_hd__dfxtp_1 _13295_ (.CLK(clknet_leaf_129_clk),
    .D(_00911_),
    .Q(\reg_module.gprf[809] ));
 sky130_fd_sc_hd__dfxtp_1 _13296_ (.CLK(clknet_leaf_130_clk),
    .D(_00912_),
    .Q(\reg_module.gprf[810] ));
 sky130_fd_sc_hd__dfxtp_1 _13297_ (.CLK(clknet_leaf_124_clk),
    .D(_00913_),
    .Q(\reg_module.gprf[811] ));
 sky130_fd_sc_hd__dfxtp_1 _13298_ (.CLK(clknet_leaf_105_clk),
    .D(_00914_),
    .Q(\reg_module.gprf[812] ));
 sky130_fd_sc_hd__dfxtp_1 _13299_ (.CLK(clknet_leaf_127_clk),
    .D(_00915_),
    .Q(\reg_module.gprf[813] ));
 sky130_fd_sc_hd__dfxtp_1 _13300_ (.CLK(clknet_leaf_112_clk),
    .D(_00916_),
    .Q(\reg_module.gprf[814] ));
 sky130_fd_sc_hd__dfxtp_1 _13301_ (.CLK(clknet_leaf_109_clk),
    .D(_00917_),
    .Q(\reg_module.gprf[815] ));
 sky130_fd_sc_hd__dfxtp_1 _13302_ (.CLK(clknet_leaf_55_clk),
    .D(_00918_),
    .Q(\reg_module.gprf[816] ));
 sky130_fd_sc_hd__dfxtp_1 _13303_ (.CLK(clknet_leaf_102_clk),
    .D(_00919_),
    .Q(\reg_module.gprf[817] ));
 sky130_fd_sc_hd__dfxtp_1 _13304_ (.CLK(clknet_leaf_121_clk),
    .D(_00920_),
    .Q(\reg_module.gprf[818] ));
 sky130_fd_sc_hd__dfxtp_1 _13305_ (.CLK(clknet_leaf_108_clk),
    .D(_00921_),
    .Q(\reg_module.gprf[819] ));
 sky130_fd_sc_hd__dfxtp_1 _13306_ (.CLK(clknet_leaf_115_clk),
    .D(_00922_),
    .Q(\reg_module.gprf[820] ));
 sky130_fd_sc_hd__dfxtp_1 _13307_ (.CLK(clknet_leaf_57_clk),
    .D(_00923_),
    .Q(\reg_module.gprf[821] ));
 sky130_fd_sc_hd__dfxtp_1 _13308_ (.CLK(clknet_leaf_65_clk),
    .D(_00924_),
    .Q(\reg_module.gprf[822] ));
 sky130_fd_sc_hd__dfxtp_1 _13309_ (.CLK(clknet_leaf_95_clk),
    .D(_00925_),
    .Q(\reg_module.gprf[823] ));
 sky130_fd_sc_hd__dfxtp_1 _13310_ (.CLK(clknet_leaf_85_clk),
    .D(_00926_),
    .Q(\reg_module.gprf[824] ));
 sky130_fd_sc_hd__dfxtp_1 _13311_ (.CLK(clknet_leaf_91_clk),
    .D(_00927_),
    .Q(\reg_module.gprf[825] ));
 sky130_fd_sc_hd__dfxtp_1 _13312_ (.CLK(clknet_leaf_78_clk),
    .D(_00928_),
    .Q(\reg_module.gprf[826] ));
 sky130_fd_sc_hd__dfxtp_1 _13313_ (.CLK(clknet_leaf_100_clk),
    .D(_00929_),
    .Q(\reg_module.gprf[827] ));
 sky130_fd_sc_hd__dfxtp_1 _13314_ (.CLK(clknet_leaf_94_clk),
    .D(_00930_),
    .Q(\reg_module.gprf[828] ));
 sky130_fd_sc_hd__dfxtp_1 _13315_ (.CLK(clknet_leaf_82_clk),
    .D(_00931_),
    .Q(\reg_module.gprf[829] ));
 sky130_fd_sc_hd__dfxtp_1 _13316_ (.CLK(clknet_leaf_84_clk),
    .D(_00932_),
    .Q(\reg_module.gprf[830] ));
 sky130_fd_sc_hd__dfxtp_1 _13317_ (.CLK(clknet_leaf_62_clk),
    .D(_00933_),
    .Q(\reg_module.gprf[831] ));
 sky130_fd_sc_hd__dfxtp_1 _13318_ (.CLK(clknet_leaf_25_clk),
    .D(_00934_),
    .Q(\reg_module.gprf[832] ));
 sky130_fd_sc_hd__dfxtp_1 _13319_ (.CLK(clknet_leaf_37_clk),
    .D(_00935_),
    .Q(\reg_module.gprf[833] ));
 sky130_fd_sc_hd__dfxtp_1 _13320_ (.CLK(clknet_leaf_15_clk),
    .D(_00936_),
    .Q(\reg_module.gprf[834] ));
 sky130_fd_sc_hd__dfxtp_1 _13321_ (.CLK(clknet_leaf_3_clk),
    .D(_00937_),
    .Q(\reg_module.gprf[835] ));
 sky130_fd_sc_hd__dfxtp_1 _13322_ (.CLK(clknet_leaf_36_clk),
    .D(_00938_),
    .Q(\reg_module.gprf[836] ));
 sky130_fd_sc_hd__dfxtp_1 _13323_ (.CLK(clknet_leaf_28_clk),
    .D(_00939_),
    .Q(\reg_module.gprf[837] ));
 sky130_fd_sc_hd__dfxtp_1 _13324_ (.CLK(clknet_leaf_5_clk),
    .D(_00940_),
    .Q(\reg_module.gprf[838] ));
 sky130_fd_sc_hd__dfxtp_1 _13325_ (.CLK(clknet_leaf_8_clk),
    .D(_00941_),
    .Q(\reg_module.gprf[839] ));
 sky130_fd_sc_hd__dfxtp_1 _13326_ (.CLK(clknet_leaf_30_clk),
    .D(_00942_),
    .Q(\reg_module.gprf[840] ));
 sky130_fd_sc_hd__dfxtp_1 _13327_ (.CLK(clknet_leaf_124_clk),
    .D(_00943_),
    .Q(\reg_module.gprf[841] ));
 sky130_fd_sc_hd__dfxtp_1 _13328_ (.CLK(clknet_leaf_130_clk),
    .D(_00944_),
    .Q(\reg_module.gprf[842] ));
 sky130_fd_sc_hd__dfxtp_1 _13329_ (.CLK(clknet_leaf_122_clk),
    .D(_00945_),
    .Q(\reg_module.gprf[843] ));
 sky130_fd_sc_hd__dfxtp_1 _13330_ (.CLK(clknet_leaf_104_clk),
    .D(_00946_),
    .Q(\reg_module.gprf[844] ));
 sky130_fd_sc_hd__dfxtp_1 _13331_ (.CLK(clknet_leaf_14_clk),
    .D(_00947_),
    .Q(\reg_module.gprf[845] ));
 sky130_fd_sc_hd__dfxtp_1 _13332_ (.CLK(clknet_leaf_113_clk),
    .D(_00948_),
    .Q(\reg_module.gprf[846] ));
 sky130_fd_sc_hd__dfxtp_1 _13333_ (.CLK(clknet_leaf_108_clk),
    .D(_00949_),
    .Q(\reg_module.gprf[847] ));
 sky130_fd_sc_hd__dfxtp_1 _13334_ (.CLK(clknet_leaf_55_clk),
    .D(_00950_),
    .Q(\reg_module.gprf[848] ));
 sky130_fd_sc_hd__dfxtp_1 _13335_ (.CLK(clknet_leaf_101_clk),
    .D(_00951_),
    .Q(\reg_module.gprf[849] ));
 sky130_fd_sc_hd__dfxtp_1 _13336_ (.CLK(clknet_leaf_102_clk),
    .D(_00952_),
    .Q(\reg_module.gprf[850] ));
 sky130_fd_sc_hd__dfxtp_1 _13337_ (.CLK(clknet_leaf_80_clk),
    .D(_00953_),
    .Q(\reg_module.gprf[851] ));
 sky130_fd_sc_hd__dfxtp_1 _13338_ (.CLK(clknet_leaf_113_clk),
    .D(_00954_),
    .Q(\reg_module.gprf[852] ));
 sky130_fd_sc_hd__dfxtp_1 _13339_ (.CLK(clknet_leaf_58_clk),
    .D(_00955_),
    .Q(\reg_module.gprf[853] ));
 sky130_fd_sc_hd__dfxtp_1 _13340_ (.CLK(clknet_leaf_65_clk),
    .D(_00956_),
    .Q(\reg_module.gprf[854] ));
 sky130_fd_sc_hd__dfxtp_1 _13341_ (.CLK(clknet_leaf_95_clk),
    .D(_00957_),
    .Q(\reg_module.gprf[855] ));
 sky130_fd_sc_hd__dfxtp_1 _13342_ (.CLK(clknet_leaf_86_clk),
    .D(_00958_),
    .Q(\reg_module.gprf[856] ));
 sky130_fd_sc_hd__dfxtp_1 _13343_ (.CLK(clknet_leaf_91_clk),
    .D(_00959_),
    .Q(\reg_module.gprf[857] ));
 sky130_fd_sc_hd__dfxtp_1 _13344_ (.CLK(clknet_leaf_79_clk),
    .D(_00960_),
    .Q(\reg_module.gprf[858] ));
 sky130_fd_sc_hd__dfxtp_1 _13345_ (.CLK(clknet_leaf_100_clk),
    .D(_00961_),
    .Q(\reg_module.gprf[859] ));
 sky130_fd_sc_hd__dfxtp_1 _13346_ (.CLK(clknet_leaf_93_clk),
    .D(_00962_),
    .Q(\reg_module.gprf[860] ));
 sky130_fd_sc_hd__dfxtp_1 _13347_ (.CLK(clknet_leaf_81_clk),
    .D(_00963_),
    .Q(\reg_module.gprf[861] ));
 sky130_fd_sc_hd__dfxtp_1 _13348_ (.CLK(clknet_leaf_84_clk),
    .D(_00964_),
    .Q(\reg_module.gprf[862] ));
 sky130_fd_sc_hd__dfxtp_1 _13349_ (.CLK(clknet_leaf_63_clk),
    .D(_00965_),
    .Q(\reg_module.gprf[863] ));
 sky130_fd_sc_hd__dfxtp_1 _13350_ (.CLK(clknet_leaf_25_clk),
    .D(_00966_),
    .Q(\reg_module.gprf[864] ));
 sky130_fd_sc_hd__dfxtp_1 _13351_ (.CLK(clknet_leaf_37_clk),
    .D(_00967_),
    .Q(\reg_module.gprf[865] ));
 sky130_fd_sc_hd__dfxtp_1 _13352_ (.CLK(clknet_leaf_15_clk),
    .D(_00968_),
    .Q(\reg_module.gprf[866] ));
 sky130_fd_sc_hd__dfxtp_1 _13353_ (.CLK(clknet_leaf_13_clk),
    .D(_00969_),
    .Q(\reg_module.gprf[867] ));
 sky130_fd_sc_hd__dfxtp_1 _13354_ (.CLK(clknet_leaf_35_clk),
    .D(_00970_),
    .Q(\reg_module.gprf[868] ));
 sky130_fd_sc_hd__dfxtp_1 _13355_ (.CLK(clknet_leaf_28_clk),
    .D(_00971_),
    .Q(\reg_module.gprf[869] ));
 sky130_fd_sc_hd__dfxtp_1 _13356_ (.CLK(clknet_leaf_5_clk),
    .D(_00972_),
    .Q(\reg_module.gprf[870] ));
 sky130_fd_sc_hd__dfxtp_1 _13357_ (.CLK(clknet_leaf_8_clk),
    .D(_00973_),
    .Q(\reg_module.gprf[871] ));
 sky130_fd_sc_hd__dfxtp_1 _13358_ (.CLK(clknet_leaf_31_clk),
    .D(_00974_),
    .Q(\reg_module.gprf[872] ));
 sky130_fd_sc_hd__dfxtp_1 _13359_ (.CLK(clknet_leaf_124_clk),
    .D(_00975_),
    .Q(\reg_module.gprf[873] ));
 sky130_fd_sc_hd__dfxtp_1 _13360_ (.CLK(clknet_leaf_129_clk),
    .D(_00976_),
    .Q(\reg_module.gprf[874] ));
 sky130_fd_sc_hd__dfxtp_1 _13361_ (.CLK(clknet_leaf_122_clk),
    .D(_00977_),
    .Q(\reg_module.gprf[875] ));
 sky130_fd_sc_hd__dfxtp_1 _13362_ (.CLK(clknet_leaf_105_clk),
    .D(_00978_),
    .Q(\reg_module.gprf[876] ));
 sky130_fd_sc_hd__dfxtp_1 _13363_ (.CLK(clknet_leaf_127_clk),
    .D(_00979_),
    .Q(\reg_module.gprf[877] ));
 sky130_fd_sc_hd__dfxtp_1 _13364_ (.CLK(clknet_leaf_112_clk),
    .D(_00980_),
    .Q(\reg_module.gprf[878] ));
 sky130_fd_sc_hd__dfxtp_1 _13365_ (.CLK(clknet_leaf_108_clk),
    .D(_00981_),
    .Q(\reg_module.gprf[879] ));
 sky130_fd_sc_hd__dfxtp_1 _13366_ (.CLK(clknet_leaf_55_clk),
    .D(_00982_),
    .Q(\reg_module.gprf[880] ));
 sky130_fd_sc_hd__dfxtp_1 _13367_ (.CLK(clknet_leaf_100_clk),
    .D(_00983_),
    .Q(\reg_module.gprf[881] ));
 sky130_fd_sc_hd__dfxtp_1 _13368_ (.CLK(clknet_leaf_102_clk),
    .D(_00984_),
    .Q(\reg_module.gprf[882] ));
 sky130_fd_sc_hd__dfxtp_1 _13369_ (.CLK(clknet_leaf_80_clk),
    .D(_00985_),
    .Q(\reg_module.gprf[883] ));
 sky130_fd_sc_hd__dfxtp_1 _13370_ (.CLK(clknet_leaf_114_clk),
    .D(_00986_),
    .Q(\reg_module.gprf[884] ));
 sky130_fd_sc_hd__dfxtp_1 _13371_ (.CLK(clknet_leaf_58_clk),
    .D(_00987_),
    .Q(\reg_module.gprf[885] ));
 sky130_fd_sc_hd__dfxtp_1 _13372_ (.CLK(clknet_leaf_66_clk),
    .D(_00988_),
    .Q(\reg_module.gprf[886] ));
 sky130_fd_sc_hd__dfxtp_1 _13373_ (.CLK(clknet_leaf_94_clk),
    .D(_00989_),
    .Q(\reg_module.gprf[887] ));
 sky130_fd_sc_hd__dfxtp_1 _13374_ (.CLK(clknet_leaf_86_clk),
    .D(_00990_),
    .Q(\reg_module.gprf[888] ));
 sky130_fd_sc_hd__dfxtp_1 _13375_ (.CLK(clknet_leaf_91_clk),
    .D(_00991_),
    .Q(\reg_module.gprf[889] ));
 sky130_fd_sc_hd__dfxtp_1 _13376_ (.CLK(clknet_leaf_81_clk),
    .D(_00992_),
    .Q(\reg_module.gprf[890] ));
 sky130_fd_sc_hd__dfxtp_1 _13377_ (.CLK(clknet_leaf_95_clk),
    .D(_00993_),
    .Q(\reg_module.gprf[891] ));
 sky130_fd_sc_hd__dfxtp_1 _13378_ (.CLK(clknet_leaf_93_clk),
    .D(_00994_),
    .Q(\reg_module.gprf[892] ));
 sky130_fd_sc_hd__dfxtp_1 _13379_ (.CLK(clknet_leaf_81_clk),
    .D(_00995_),
    .Q(\reg_module.gprf[893] ));
 sky130_fd_sc_hd__dfxtp_1 _13380_ (.CLK(clknet_leaf_84_clk),
    .D(_00996_),
    .Q(\reg_module.gprf[894] ));
 sky130_fd_sc_hd__dfxtp_1 _13381_ (.CLK(clknet_leaf_63_clk),
    .D(_00997_),
    .Q(\reg_module.gprf[895] ));
 sky130_fd_sc_hd__dfxtp_1 _13382_ (.CLK(clknet_leaf_26_clk),
    .D(_00998_),
    .Q(\reg_module.gprf[896] ));
 sky130_fd_sc_hd__dfxtp_1 _13383_ (.CLK(clknet_leaf_38_clk),
    .D(_00999_),
    .Q(\reg_module.gprf[897] ));
 sky130_fd_sc_hd__dfxtp_1 _13384_ (.CLK(clknet_leaf_16_clk),
    .D(_01000_),
    .Q(\reg_module.gprf[898] ));
 sky130_fd_sc_hd__dfxtp_1 _13385_ (.CLK(clknet_leaf_12_clk),
    .D(_01001_),
    .Q(\reg_module.gprf[899] ));
 sky130_fd_sc_hd__dfxtp_1 _13386_ (.CLK(clknet_leaf_37_clk),
    .D(_01002_),
    .Q(\reg_module.gprf[900] ));
 sky130_fd_sc_hd__dfxtp_1 _13387_ (.CLK(clknet_leaf_28_clk),
    .D(_01003_),
    .Q(\reg_module.gprf[901] ));
 sky130_fd_sc_hd__dfxtp_1 _13388_ (.CLK(clknet_leaf_5_clk),
    .D(_01004_),
    .Q(\reg_module.gprf[902] ));
 sky130_fd_sc_hd__dfxtp_1 _13389_ (.CLK(clknet_leaf_7_clk),
    .D(_01005_),
    .Q(\reg_module.gprf[903] ));
 sky130_fd_sc_hd__dfxtp_1 _13390_ (.CLK(clknet_leaf_32_clk),
    .D(_01006_),
    .Q(\reg_module.gprf[904] ));
 sky130_fd_sc_hd__dfxtp_1 _13391_ (.CLK(clknet_leaf_129_clk),
    .D(_01007_),
    .Q(\reg_module.gprf[905] ));
 sky130_fd_sc_hd__dfxtp_1 _13392_ (.CLK(clknet_leaf_131_clk),
    .D(_01008_),
    .Q(\reg_module.gprf[906] ));
 sky130_fd_sc_hd__dfxtp_1 _13393_ (.CLK(clknet_leaf_123_clk),
    .D(_01009_),
    .Q(\reg_module.gprf[907] ));
 sky130_fd_sc_hd__dfxtp_1 _13394_ (.CLK(clknet_leaf_109_clk),
    .D(_01010_),
    .Q(\reg_module.gprf[908] ));
 sky130_fd_sc_hd__dfxtp_1 _13395_ (.CLK(clknet_leaf_127_clk),
    .D(_01011_),
    .Q(\reg_module.gprf[909] ));
 sky130_fd_sc_hd__dfxtp_1 _13396_ (.CLK(clknet_leaf_19_clk),
    .D(_01012_),
    .Q(\reg_module.gprf[910] ));
 sky130_fd_sc_hd__dfxtp_1 _13397_ (.CLK(clknet_leaf_77_clk),
    .D(_01013_),
    .Q(\reg_module.gprf[911] ));
 sky130_fd_sc_hd__dfxtp_1 _13398_ (.CLK(clknet_leaf_53_clk),
    .D(_01014_),
    .Q(\reg_module.gprf[912] ));
 sky130_fd_sc_hd__dfxtp_1 _13399_ (.CLK(clknet_leaf_101_clk),
    .D(_01015_),
    .Q(\reg_module.gprf[913] ));
 sky130_fd_sc_hd__dfxtp_1 _13400_ (.CLK(clknet_leaf_121_clk),
    .D(_01016_),
    .Q(\reg_module.gprf[914] ));
 sky130_fd_sc_hd__dfxtp_1 _13401_ (.CLK(clknet_leaf_107_clk),
    .D(_01017_),
    .Q(\reg_module.gprf[915] ));
 sky130_fd_sc_hd__dfxtp_1 _13402_ (.CLK(clknet_leaf_114_clk),
    .D(_01018_),
    .Q(\reg_module.gprf[916] ));
 sky130_fd_sc_hd__dfxtp_1 _13403_ (.CLK(clknet_leaf_56_clk),
    .D(_01019_),
    .Q(\reg_module.gprf[917] ));
 sky130_fd_sc_hd__dfxtp_1 _13404_ (.CLK(clknet_leaf_63_clk),
    .D(_01020_),
    .Q(\reg_module.gprf[918] ));
 sky130_fd_sc_hd__dfxtp_1 _13405_ (.CLK(clknet_leaf_96_clk),
    .D(_01021_),
    .Q(\reg_module.gprf[919] ));
 sky130_fd_sc_hd__dfxtp_1 _13406_ (.CLK(clknet_leaf_85_clk),
    .D(_01022_),
    .Q(\reg_module.gprf[920] ));
 sky130_fd_sc_hd__dfxtp_1 _13407_ (.CLK(clknet_leaf_86_clk),
    .D(_01023_),
    .Q(\reg_module.gprf[921] ));
 sky130_fd_sc_hd__dfxtp_1 _13408_ (.CLK(clknet_leaf_78_clk),
    .D(_01024_),
    .Q(\reg_module.gprf[922] ));
 sky130_fd_sc_hd__dfxtp_1 _13409_ (.CLK(clknet_leaf_100_clk),
    .D(_01025_),
    .Q(\reg_module.gprf[923] ));
 sky130_fd_sc_hd__dfxtp_1 _13410_ (.CLK(clknet_leaf_91_clk),
    .D(_01026_),
    .Q(\reg_module.gprf[924] ));
 sky130_fd_sc_hd__dfxtp_1 _13411_ (.CLK(clknet_leaf_80_clk),
    .D(_01027_),
    .Q(\reg_module.gprf[925] ));
 sky130_fd_sc_hd__dfxtp_1 _13412_ (.CLK(clknet_leaf_66_clk),
    .D(_01028_),
    .Q(\reg_module.gprf[926] ));
 sky130_fd_sc_hd__dfxtp_1 _13413_ (.CLK(clknet_leaf_59_clk),
    .D(_01029_),
    .Q(\reg_module.gprf[927] ));
 sky130_fd_sc_hd__dfxtp_1 _13414_ (.CLK(clknet_leaf_26_clk),
    .D(_01030_),
    .Q(\reg_module.gprf[928] ));
 sky130_fd_sc_hd__dfxtp_1 _13415_ (.CLK(clknet_leaf_38_clk),
    .D(_01031_),
    .Q(\reg_module.gprf[929] ));
 sky130_fd_sc_hd__dfxtp_1 _13416_ (.CLK(clknet_leaf_15_clk),
    .D(_01032_),
    .Q(\reg_module.gprf[930] ));
 sky130_fd_sc_hd__dfxtp_1 _13417_ (.CLK(clknet_leaf_12_clk),
    .D(_01033_),
    .Q(\reg_module.gprf[931] ));
 sky130_fd_sc_hd__dfxtp_1 _13418_ (.CLK(clknet_leaf_37_clk),
    .D(_01034_),
    .Q(\reg_module.gprf[932] ));
 sky130_fd_sc_hd__dfxtp_1 _13419_ (.CLK(clknet_leaf_29_clk),
    .D(_01035_),
    .Q(\reg_module.gprf[933] ));
 sky130_fd_sc_hd__dfxtp_1 _13420_ (.CLK(clknet_leaf_5_clk),
    .D(_01036_),
    .Q(\reg_module.gprf[934] ));
 sky130_fd_sc_hd__dfxtp_1 _13421_ (.CLK(clknet_leaf_7_clk),
    .D(_01037_),
    .Q(\reg_module.gprf[935] ));
 sky130_fd_sc_hd__dfxtp_1 _13422_ (.CLK(clknet_leaf_30_clk),
    .D(_01038_),
    .Q(\reg_module.gprf[936] ));
 sky130_fd_sc_hd__dfxtp_1 _13423_ (.CLK(clknet_leaf_129_clk),
    .D(_01039_),
    .Q(\reg_module.gprf[937] ));
 sky130_fd_sc_hd__dfxtp_1 _13424_ (.CLK(clknet_leaf_131_clk),
    .D(_01040_),
    .Q(\reg_module.gprf[938] ));
 sky130_fd_sc_hd__dfxtp_1 _13425_ (.CLK(clknet_leaf_124_clk),
    .D(_01041_),
    .Q(\reg_module.gprf[939] ));
 sky130_fd_sc_hd__dfxtp_1 _13426_ (.CLK(clknet_leaf_105_clk),
    .D(_01042_),
    .Q(\reg_module.gprf[940] ));
 sky130_fd_sc_hd__dfxtp_1 _13427_ (.CLK(clknet_leaf_127_clk),
    .D(_01043_),
    .Q(\reg_module.gprf[941] ));
 sky130_fd_sc_hd__dfxtp_1 _13428_ (.CLK(clknet_leaf_112_clk),
    .D(_01044_),
    .Q(\reg_module.gprf[942] ));
 sky130_fd_sc_hd__dfxtp_1 _13429_ (.CLK(clknet_leaf_110_clk),
    .D(_01045_),
    .Q(\reg_module.gprf[943] ));
 sky130_fd_sc_hd__dfxtp_1 _13430_ (.CLK(clknet_leaf_53_clk),
    .D(_01046_),
    .Q(\reg_module.gprf[944] ));
 sky130_fd_sc_hd__dfxtp_1 _13431_ (.CLK(clknet_leaf_101_clk),
    .D(_01047_),
    .Q(\reg_module.gprf[945] ));
 sky130_fd_sc_hd__dfxtp_1 _13432_ (.CLK(clknet_leaf_121_clk),
    .D(_01048_),
    .Q(\reg_module.gprf[946] ));
 sky130_fd_sc_hd__dfxtp_1 _13433_ (.CLK(clknet_leaf_108_clk),
    .D(_01049_),
    .Q(\reg_module.gprf[947] ));
 sky130_fd_sc_hd__dfxtp_1 _13434_ (.CLK(clknet_leaf_114_clk),
    .D(_01050_),
    .Q(\reg_module.gprf[948] ));
 sky130_fd_sc_hd__dfxtp_1 _13435_ (.CLK(clknet_leaf_55_clk),
    .D(_01051_),
    .Q(\reg_module.gprf[949] ));
 sky130_fd_sc_hd__dfxtp_1 _13436_ (.CLK(clknet_leaf_64_clk),
    .D(_01052_),
    .Q(\reg_module.gprf[950] ));
 sky130_fd_sc_hd__dfxtp_1 _13437_ (.CLK(clknet_leaf_96_clk),
    .D(_01053_),
    .Q(\reg_module.gprf[951] ));
 sky130_fd_sc_hd__dfxtp_1 _13438_ (.CLK(clknet_leaf_85_clk),
    .D(_01054_),
    .Q(\reg_module.gprf[952] ));
 sky130_fd_sc_hd__dfxtp_1 _13439_ (.CLK(clknet_leaf_87_clk),
    .D(_01055_),
    .Q(\reg_module.gprf[953] ));
 sky130_fd_sc_hd__dfxtp_1 _13440_ (.CLK(clknet_leaf_78_clk),
    .D(_01056_),
    .Q(\reg_module.gprf[954] ));
 sky130_fd_sc_hd__dfxtp_1 _13441_ (.CLK(clknet_leaf_100_clk),
    .D(_01057_),
    .Q(\reg_module.gprf[955] ));
 sky130_fd_sc_hd__dfxtp_1 _13442_ (.CLK(clknet_leaf_92_clk),
    .D(_01058_),
    .Q(\reg_module.gprf[956] ));
 sky130_fd_sc_hd__dfxtp_1 _13443_ (.CLK(clknet_leaf_80_clk),
    .D(_01059_),
    .Q(\reg_module.gprf[957] ));
 sky130_fd_sc_hd__dfxtp_1 _13444_ (.CLK(clknet_leaf_67_clk),
    .D(_01060_),
    .Q(\reg_module.gprf[958] ));
 sky130_fd_sc_hd__dfxtp_1 _13445_ (.CLK(clknet_leaf_59_clk),
    .D(_01061_),
    .Q(\reg_module.gprf[959] ));
 sky130_fd_sc_hd__dfxtp_1 _13446_ (.CLK(clknet_leaf_26_clk),
    .D(_01062_),
    .Q(\reg_module.gprf[960] ));
 sky130_fd_sc_hd__dfxtp_1 _13447_ (.CLK(clknet_leaf_40_clk),
    .D(_01063_),
    .Q(\reg_module.gprf[961] ));
 sky130_fd_sc_hd__dfxtp_1 _13448_ (.CLK(clknet_leaf_16_clk),
    .D(_01064_),
    .Q(\reg_module.gprf[962] ));
 sky130_fd_sc_hd__dfxtp_1 _13449_ (.CLK(clknet_leaf_13_clk),
    .D(_01065_),
    .Q(\reg_module.gprf[963] ));
 sky130_fd_sc_hd__dfxtp_1 _13450_ (.CLK(clknet_leaf_38_clk),
    .D(_01066_),
    .Q(\reg_module.gprf[964] ));
 sky130_fd_sc_hd__dfxtp_1 _13451_ (.CLK(clknet_leaf_27_clk),
    .D(_01067_),
    .Q(\reg_module.gprf[965] ));
 sky130_fd_sc_hd__dfxtp_1 _13452_ (.CLK(clknet_leaf_4_clk),
    .D(_01068_),
    .Q(\reg_module.gprf[966] ));
 sky130_fd_sc_hd__dfxtp_1 _13453_ (.CLK(clknet_leaf_9_clk),
    .D(_01069_),
    .Q(\reg_module.gprf[967] ));
 sky130_fd_sc_hd__dfxtp_1 _13454_ (.CLK(clknet_leaf_32_clk),
    .D(_01070_),
    .Q(\reg_module.gprf[968] ));
 sky130_fd_sc_hd__dfxtp_1 _13455_ (.CLK(clknet_leaf_124_clk),
    .D(_01071_),
    .Q(\reg_module.gprf[969] ));
 sky130_fd_sc_hd__dfxtp_1 _13456_ (.CLK(clknet_leaf_130_clk),
    .D(_01072_),
    .Q(\reg_module.gprf[970] ));
 sky130_fd_sc_hd__dfxtp_1 _13457_ (.CLK(clknet_leaf_123_clk),
    .D(_01073_),
    .Q(\reg_module.gprf[971] ));
 sky130_fd_sc_hd__dfxtp_1 _13458_ (.CLK(clknet_leaf_109_clk),
    .D(_01074_),
    .Q(\reg_module.gprf[972] ));
 sky130_fd_sc_hd__dfxtp_1 _13459_ (.CLK(clknet_leaf_126_clk),
    .D(_01075_),
    .Q(\reg_module.gprf[973] ));
 sky130_fd_sc_hd__dfxtp_1 _13460_ (.CLK(clknet_leaf_111_clk),
    .D(_01076_),
    .Q(\reg_module.gprf[974] ));
 sky130_fd_sc_hd__dfxtp_1 _13461_ (.CLK(clknet_leaf_108_clk),
    .D(_01077_),
    .Q(\reg_module.gprf[975] ));
 sky130_fd_sc_hd__dfxtp_1 _13462_ (.CLK(clknet_leaf_53_clk),
    .D(_01078_),
    .Q(\reg_module.gprf[976] ));
 sky130_fd_sc_hd__dfxtp_1 _13463_ (.CLK(clknet_leaf_101_clk),
    .D(_01079_),
    .Q(\reg_module.gprf[977] ));
 sky130_fd_sc_hd__dfxtp_1 _13464_ (.CLK(clknet_leaf_102_clk),
    .D(_01080_),
    .Q(\reg_module.gprf[978] ));
 sky130_fd_sc_hd__dfxtp_1 _13465_ (.CLK(clknet_leaf_108_clk),
    .D(_01081_),
    .Q(\reg_module.gprf[979] ));
 sky130_fd_sc_hd__dfxtp_1 _13466_ (.CLK(clknet_leaf_110_clk),
    .D(_01082_),
    .Q(\reg_module.gprf[980] ));
 sky130_fd_sc_hd__dfxtp_1 _13467_ (.CLK(clknet_leaf_57_clk),
    .D(_01083_),
    .Q(\reg_module.gprf[981] ));
 sky130_fd_sc_hd__dfxtp_1 _13468_ (.CLK(clknet_leaf_64_clk),
    .D(_01084_),
    .Q(\reg_module.gprf[982] ));
 sky130_fd_sc_hd__dfxtp_1 _13469_ (.CLK(clknet_leaf_95_clk),
    .D(_01085_),
    .Q(\reg_module.gprf[983] ));
 sky130_fd_sc_hd__dfxtp_1 _13470_ (.CLK(clknet_leaf_85_clk),
    .D(_01086_),
    .Q(\reg_module.gprf[984] ));
 sky130_fd_sc_hd__dfxtp_1 _13471_ (.CLK(clknet_leaf_86_clk),
    .D(_01087_),
    .Q(\reg_module.gprf[985] ));
 sky130_fd_sc_hd__dfxtp_1 _13472_ (.CLK(clknet_leaf_82_clk),
    .D(_01088_),
    .Q(\reg_module.gprf[986] ));
 sky130_fd_sc_hd__dfxtp_1 _13473_ (.CLK(clknet_leaf_100_clk),
    .D(_01089_),
    .Q(\reg_module.gprf[987] ));
 sky130_fd_sc_hd__dfxtp_1 _13474_ (.CLK(clknet_leaf_92_clk),
    .D(_01090_),
    .Q(\reg_module.gprf[988] ));
 sky130_fd_sc_hd__dfxtp_1 _13475_ (.CLK(clknet_leaf_80_clk),
    .D(_01091_),
    .Q(\reg_module.gprf[989] ));
 sky130_fd_sc_hd__dfxtp_1 _13476_ (.CLK(clknet_leaf_66_clk),
    .D(_01092_),
    .Q(\reg_module.gprf[990] ));
 sky130_fd_sc_hd__dfxtp_1 _13477_ (.CLK(clknet_leaf_59_clk),
    .D(_01093_),
    .Q(\reg_module.gprf[991] ));
 sky130_fd_sc_hd__dfxtp_1 _13478_ (.CLK(clknet_leaf_26_clk),
    .D(_01094_),
    .Q(\reg_module.gprf[992] ));
 sky130_fd_sc_hd__dfxtp_1 _13479_ (.CLK(clknet_leaf_40_clk),
    .D(_01095_),
    .Q(\reg_module.gprf[993] ));
 sky130_fd_sc_hd__dfxtp_1 _13480_ (.CLK(clknet_leaf_15_clk),
    .D(_01096_),
    .Q(\reg_module.gprf[994] ));
 sky130_fd_sc_hd__dfxtp_1 _13481_ (.CLK(clknet_leaf_12_clk),
    .D(_01097_),
    .Q(\reg_module.gprf[995] ));
 sky130_fd_sc_hd__dfxtp_1 _13482_ (.CLK(clknet_leaf_38_clk),
    .D(_01098_),
    .Q(\reg_module.gprf[996] ));
 sky130_fd_sc_hd__dfxtp_1 _13483_ (.CLK(clknet_leaf_27_clk),
    .D(_01099_),
    .Q(\reg_module.gprf[997] ));
 sky130_fd_sc_hd__dfxtp_1 _13484_ (.CLK(clknet_leaf_4_clk),
    .D(_01100_),
    .Q(\reg_module.gprf[998] ));
 sky130_fd_sc_hd__dfxtp_1 _13485_ (.CLK(clknet_leaf_7_clk),
    .D(_01101_),
    .Q(\reg_module.gprf[999] ));
 sky130_fd_sc_hd__dfxtp_1 _13486_ (.CLK(clknet_leaf_32_clk),
    .D(_01102_),
    .Q(\reg_module.gprf[1000] ));
 sky130_fd_sc_hd__dfxtp_1 _13487_ (.CLK(clknet_leaf_129_clk),
    .D(_01103_),
    .Q(\reg_module.gprf[1001] ));
 sky130_fd_sc_hd__dfxtp_1 _13488_ (.CLK(clknet_leaf_131_clk),
    .D(_01104_),
    .Q(\reg_module.gprf[1002] ));
 sky130_fd_sc_hd__dfxtp_1 _13489_ (.CLK(clknet_leaf_123_clk),
    .D(_01105_),
    .Q(\reg_module.gprf[1003] ));
 sky130_fd_sc_hd__dfxtp_1 _13490_ (.CLK(clknet_leaf_109_clk),
    .D(_01106_),
    .Q(\reg_module.gprf[1004] ));
 sky130_fd_sc_hd__dfxtp_1 _13491_ (.CLK(clknet_leaf_126_clk),
    .D(_01107_),
    .Q(\reg_module.gprf[1005] ));
 sky130_fd_sc_hd__dfxtp_1 _13492_ (.CLK(clknet_leaf_112_clk),
    .D(_01108_),
    .Q(\reg_module.gprf[1006] ));
 sky130_fd_sc_hd__dfxtp_1 _13493_ (.CLK(clknet_leaf_108_clk),
    .D(_01109_),
    .Q(\reg_module.gprf[1007] ));
 sky130_fd_sc_hd__dfxtp_1 _13494_ (.CLK(clknet_leaf_56_clk),
    .D(_01110_),
    .Q(\reg_module.gprf[1008] ));
 sky130_fd_sc_hd__dfxtp_1 _13495_ (.CLK(clknet_leaf_100_clk),
    .D(_01111_),
    .Q(\reg_module.gprf[1009] ));
 sky130_fd_sc_hd__dfxtp_1 _13496_ (.CLK(clknet_leaf_121_clk),
    .D(_01112_),
    .Q(\reg_module.gprf[1010] ));
 sky130_fd_sc_hd__dfxtp_1 _13497_ (.CLK(clknet_leaf_108_clk),
    .D(_01113_),
    .Q(\reg_module.gprf[1011] ));
 sky130_fd_sc_hd__dfxtp_1 _13498_ (.CLK(clknet_leaf_110_clk),
    .D(_01114_),
    .Q(\reg_module.gprf[1012] ));
 sky130_fd_sc_hd__dfxtp_1 _13499_ (.CLK(clknet_leaf_57_clk),
    .D(_01115_),
    .Q(\reg_module.gprf[1013] ));
 sky130_fd_sc_hd__dfxtp_1 _13500_ (.CLK(clknet_leaf_64_clk),
    .D(_01116_),
    .Q(\reg_module.gprf[1014] ));
 sky130_fd_sc_hd__dfxtp_1 _13501_ (.CLK(clknet_leaf_95_clk),
    .D(_01117_),
    .Q(\reg_module.gprf[1015] ));
 sky130_fd_sc_hd__dfxtp_1 _13502_ (.CLK(clknet_leaf_85_clk),
    .D(_01118_),
    .Q(\reg_module.gprf[1016] ));
 sky130_fd_sc_hd__dfxtp_1 _13503_ (.CLK(clknet_leaf_86_clk),
    .D(_01119_),
    .Q(\reg_module.gprf[1017] ));
 sky130_fd_sc_hd__dfxtp_1 _13504_ (.CLK(clknet_leaf_82_clk),
    .D(_01120_),
    .Q(\reg_module.gprf[1018] ));
 sky130_fd_sc_hd__dfxtp_1 _13505_ (.CLK(clknet_leaf_100_clk),
    .D(_01121_),
    .Q(\reg_module.gprf[1019] ));
 sky130_fd_sc_hd__dfxtp_1 _13506_ (.CLK(clknet_leaf_92_clk),
    .D(_01122_),
    .Q(\reg_module.gprf[1020] ));
 sky130_fd_sc_hd__dfxtp_1 _13507_ (.CLK(clknet_leaf_89_clk),
    .D(_01123_),
    .Q(\reg_module.gprf[1021] ));
 sky130_fd_sc_hd__dfxtp_1 _13508_ (.CLK(clknet_leaf_66_clk),
    .D(_01124_),
    .Q(\reg_module.gprf[1022] ));
 sky130_fd_sc_hd__dfxtp_1 _13509_ (.CLK(clknet_leaf_59_clk),
    .D(_01125_),
    .Q(\reg_module.gprf[1023] ));
 sky130_fd_sc_hd__dfxtp_4 _13510_ (.CLK(clknet_leaf_46_clk),
    .D(_01126_),
    .Q(net157));
 sky130_fd_sc_hd__dfxtp_4 _13511_ (.CLK(clknet_leaf_46_clk),
    .D(_01127_),
    .Q(net160));
 sky130_fd_sc_hd__dfxtp_2 _13512_ (.CLK(clknet_leaf_46_clk),
    .D(_01128_),
    .Q(net161));
 sky130_fd_sc_hd__dfxtp_2 _13513_ (.CLK(clknet_leaf_23_clk),
    .D(_01129_),
    .Q(net162));
 sky130_fd_sc_hd__dfxtp_2 _13514_ (.CLK(clknet_leaf_21_clk),
    .D(_01130_),
    .Q(net163));
 sky130_fd_sc_hd__dfxtp_2 _13515_ (.CLK(clknet_leaf_21_clk),
    .D(_01131_),
    .Q(net164));
 sky130_fd_sc_hd__dfxtp_2 _13516_ (.CLK(clknet_leaf_21_clk),
    .D(_01132_),
    .Q(net165));
 sky130_fd_sc_hd__dfxtp_4 _13517_ (.CLK(clknet_leaf_21_clk),
    .D(_01133_),
    .Q(net166));
 sky130_fd_sc_hd__dfxtp_2 _13518_ (.CLK(clknet_leaf_20_clk),
    .D(_01134_),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_2 _13519_ (.CLK(clknet_leaf_19_clk),
    .D(_01135_),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_2 _13520_ (.CLK(clknet_leaf_19_clk),
    .D(_01136_),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_2 _13521_ (.CLK(clknet_leaf_49_clk),
    .D(_01137_),
    .Q(net139));
 sky130_fd_sc_hd__dfxtp_2 _13522_ (.CLK(clknet_leaf_49_clk),
    .D(_01138_),
    .Q(net140));
 sky130_fd_sc_hd__dfxtp_4 _13523_ (.CLK(clknet_leaf_50_clk),
    .D(_01139_),
    .Q(net141));
 sky130_fd_sc_hd__dfxtp_2 _13524_ (.CLK(clknet_leaf_50_clk),
    .D(_01140_),
    .Q(net142));
 sky130_fd_sc_hd__dfxtp_4 _13525_ (.CLK(clknet_leaf_51_clk),
    .D(_01141_),
    .Q(net143));
 sky130_fd_sc_hd__dfxtp_2 _13526_ (.CLK(clknet_leaf_50_clk),
    .D(_01142_),
    .Q(net144));
 sky130_fd_sc_hd__dfxtp_2 _13527_ (.CLK(clknet_leaf_75_clk),
    .D(_01143_),
    .Q(net145));
 sky130_fd_sc_hd__dfxtp_2 _13528_ (.CLK(clknet_leaf_75_clk),
    .D(_01144_),
    .Q(net147));
 sky130_fd_sc_hd__dfxtp_4 _13529_ (.CLK(clknet_leaf_75_clk),
    .D(_01145_),
    .Q(net148));
 sky130_fd_sc_hd__dfxtp_2 _13530_ (.CLK(clknet_leaf_74_clk),
    .D(_01146_),
    .Q(net149));
 sky130_fd_sc_hd__dfxtp_2 _13531_ (.CLK(clknet_leaf_74_clk),
    .D(_01147_),
    .Q(net150));
 sky130_fd_sc_hd__dfxtp_2 _13532_ (.CLK(clknet_leaf_69_clk),
    .D(_01148_),
    .Q(net151));
 sky130_fd_sc_hd__dfxtp_2 _13533_ (.CLK(clknet_leaf_69_clk),
    .D(_01149_),
    .Q(net152));
 sky130_fd_sc_hd__dfxtp_2 _13534_ (.CLK(clknet_leaf_70_clk),
    .D(_01150_),
    .Q(net153));
 sky130_fd_sc_hd__dfxtp_2 _13535_ (.CLK(clknet_leaf_70_clk),
    .D(_01151_),
    .Q(net154));
 sky130_fd_sc_hd__dfxtp_2 _13536_ (.CLK(clknet_leaf_71_clk),
    .D(_01152_),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_2 _13537_ (.CLK(clknet_leaf_71_clk),
    .D(_01153_),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_2 _13538_ (.CLK(clknet_leaf_61_clk),
    .D(_01154_),
    .Q(net158));
 sky130_fd_sc_hd__dfxtp_2 _13539_ (.CLK(clknet_leaf_61_clk),
    .D(_01155_),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_2 _13540_ (.CLK(clknet_leaf_42_clk),
    .D(_01156_),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_1 _13541_ (.CLK(clknet_leaf_42_clk),
    .D(_01157_),
    .Q(net146));
 sky130_fd_sc_hd__dfxtp_1 _13542_ (.CLK(clknet_leaf_42_clk),
    .D(_01158_),
    .Q(\brancher.rJumping ));
 sky130_fd_sc_hd__dfxtp_1 _13543_ (.CLK(clknet_leaf_42_clk),
    .D(_01159_),
    .Q(\brancher.imm13_b[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13544_ (.CLK(clknet_leaf_41_clk),
    .D(_01160_),
    .Q(\brancher.imm13_b[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13545_ (.CLK(clknet_leaf_40_clk),
    .D(_01161_),
    .Q(\brancher.imm13_b[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13546_ (.CLK(clknet_leaf_40_clk),
    .D(_01162_),
    .Q(\brancher.imm13_b[4] ));
 sky130_fd_sc_hd__dfxtp_2 _13547_ (.CLK(clknet_leaf_25_clk),
    .D(_01163_),
    .Q(\brancher.imm13_b[5] ));
 sky130_fd_sc_hd__dfxtp_2 _13548_ (.CLK(clknet_leaf_24_clk),
    .D(_01164_),
    .Q(\brancher.imm13_b[6] ));
 sky130_fd_sc_hd__dfxtp_2 _13549_ (.CLK(clknet_leaf_25_clk),
    .D(_01165_),
    .Q(\brancher.imm13_b[7] ));
 sky130_fd_sc_hd__dfxtp_2 _13550_ (.CLK(clknet_leaf_47_clk),
    .D(_01166_),
    .Q(\brancher.imm13_b[8] ));
 sky130_fd_sc_hd__dfxtp_2 _13551_ (.CLK(clknet_leaf_23_clk),
    .D(_01167_),
    .Q(\brancher.imm13_b[9] ));
 sky130_fd_sc_hd__dfxtp_2 _13552_ (.CLK(clknet_leaf_42_clk),
    .D(_01168_),
    .Q(\brancher.imm13_b[10] ));
 sky130_fd_sc_hd__dfxtp_2 _13553_ (.CLK(clknet_leaf_39_clk),
    .D(_01169_),
    .Q(\brancher.imm13_b[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13554_ (.CLK(clknet_leaf_47_clk),
    .D(_01170_),
    .Q(\brancher.imm13_b[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13555_ (.CLK(clknet_leaf_42_clk),
    .D(_01171_),
    .Q(\brancher.pc_return[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13556_ (.CLK(clknet_leaf_42_clk),
    .D(_01172_),
    .Q(\brancher.pc_return[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13557_ (.CLK(clknet_leaf_45_clk),
    .D(_01173_),
    .Q(\brancher.pc_return[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13558_ (.CLK(clknet_leaf_41_clk),
    .D(_01174_),
    .Q(\brancher.pc_return[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13559_ (.CLK(clknet_leaf_45_clk),
    .D(_01175_),
    .Q(\brancher.pc_return[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13560_ (.CLK(clknet_leaf_24_clk),
    .D(_01176_),
    .Q(\brancher.pc_return[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13561_ (.CLK(clknet_leaf_22_clk),
    .D(_01177_),
    .Q(\brancher.pc_return[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13562_ (.CLK(clknet_leaf_21_clk),
    .D(_01178_),
    .Q(\brancher.pc_return[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13563_ (.CLK(clknet_leaf_23_clk),
    .D(_01179_),
    .Q(\brancher.pc_return[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13564_ (.CLK(clknet_leaf_23_clk),
    .D(_01180_),
    .Q(\brancher.pc_return[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13565_ (.CLK(clknet_leaf_20_clk),
    .D(_01181_),
    .Q(\brancher.pc_return[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13566_ (.CLK(clknet_leaf_20_clk),
    .D(_01182_),
    .Q(\brancher.pc_return[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13567_ (.CLK(clknet_leaf_48_clk),
    .D(_01183_),
    .Q(\brancher.pc_return[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13568_ (.CLK(clknet_leaf_48_clk),
    .D(_01184_),
    .Q(\brancher.pc_return[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13569_ (.CLK(clknet_leaf_48_clk),
    .D(_01185_),
    .Q(\brancher.pc_return[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13570_ (.CLK(clknet_leaf_48_clk),
    .D(_01186_),
    .Q(\brancher.pc_return[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13571_ (.CLK(clknet_leaf_48_clk),
    .D(_01187_),
    .Q(\brancher.pc_return[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13572_ (.CLK(clknet_leaf_50_clk),
    .D(_01188_),
    .Q(\brancher.pc_return[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13573_ (.CLK(clknet_leaf_51_clk),
    .D(_01189_),
    .Q(\brancher.pc_return[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13574_ (.CLK(clknet_leaf_51_clk),
    .D(net1307),
    .Q(\brancher.pc_return[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13575_ (.CLK(clknet_leaf_51_clk),
    .D(_01191_),
    .Q(\brancher.pc_return[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13576_ (.CLK(clknet_leaf_73_clk),
    .D(_01192_),
    .Q(\brancher.pc_return[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13577_ (.CLK(clknet_leaf_73_clk),
    .D(_01193_),
    .Q(\brancher.pc_return[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13578_ (.CLK(clknet_leaf_73_clk),
    .D(_01194_),
    .Q(\brancher.pc_return[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13579_ (.CLK(clknet_leaf_73_clk),
    .D(_01195_),
    .Q(\brancher.pc_return[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13580_ (.CLK(clknet_leaf_73_clk),
    .D(_01196_),
    .Q(\brancher.pc_return[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13581_ (.CLK(clknet_leaf_72_clk),
    .D(_01197_),
    .Q(\brancher.pc_return[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13582_ (.CLK(clknet_leaf_73_clk),
    .D(_01198_),
    .Q(\brancher.pc_return[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13583_ (.CLK(clknet_leaf_72_clk),
    .D(_01199_),
    .Q(\brancher.pc_return[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13584_ (.CLK(clknet_leaf_72_clk),
    .D(_01200_),
    .Q(\brancher.pc_return[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13585_ (.CLK(clknet_leaf_72_clk),
    .D(_01201_),
    .Q(\brancher.pc_return[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13586_ (.CLK(clknet_leaf_52_clk),
    .D(_01202_),
    .Q(\brancher.pc_return[31] ));
 sky130_fd_sc_hd__clkbuf_1 _13587_ (.A(\brancher.funct3[2] ),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _13588_ (.A(wRamWordEn),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _13589_ (.A(wRamHalfEn),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _13590_ (.A(wRamByteEn),
    .X(net70));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_2821 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(clkEn),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(dataBusIn[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(dataBusIn[10]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(dataBusIn[11]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input5 (.A(dataBusIn[12]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(dataBusIn[13]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(dataBusIn[14]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(dataBusIn[15]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(dataBusIn[16]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(dataBusIn[17]),
    .X(net10));
 sky130_fd_sc_hd__dlymetal6s2s_1 input11 (.A(dataBusIn[18]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(dataBusIn[19]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(dataBusIn[1]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(dataBusIn[20]),
    .X(net14));
 sky130_fd_sc_hd__dlymetal6s2s_1 input15 (.A(dataBusIn[21]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(dataBusIn[22]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(dataBusIn[23]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(dataBusIn[24]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(dataBusIn[25]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(dataBusIn[26]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(dataBusIn[27]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(dataBusIn[28]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(dataBusIn[29]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(dataBusIn[2]),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(dataBusIn[30]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(dataBusIn[31]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(dataBusIn[3]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(dataBusIn[4]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(dataBusIn[5]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(dataBusIn[6]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(dataBusIn[7]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(dataBusIn[8]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(dataBusIn[9]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(inst_in[0]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(inst_in[10]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(inst_in[11]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(inst_in[12]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(inst_in[13]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(inst_in[14]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(inst_in[15]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(inst_in[16]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(inst_in[17]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(inst_in[18]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(inst_in[19]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(inst_in[1]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(inst_in[20]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(inst_in[21]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(inst_in[22]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(inst_in[23]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(inst_in[24]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(inst_in[25]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(inst_in[26]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(inst_in[27]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(inst_in[28]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(inst_in[29]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(inst_in[2]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(inst_in[30]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(inst_in[31]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(inst_in[3]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input60 (.A(inst_in[4]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(inst_in[5]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(inst_in[6]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(inst_in[7]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(inst_in[8]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(inst_in[9]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(rstB),
    .X(net66));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(RamMode[0]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(RamMode[1]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(RamMode[2]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(RamMode[3]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(addr[0]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(addr[10]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(addr[11]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(addr[12]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(addr[13]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(addr[14]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(addr[15]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(addr[16]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(addr[17]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(addr[18]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(addr[19]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(addr[1]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(addr[20]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(addr[21]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(addr[22]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(addr[23]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(addr[24]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(addr[25]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(addr[26]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(addr[27]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(addr[28]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(addr[29]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(addr[2]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(addr[30]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(addr[31]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(addr[3]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(addr[4]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(addr[5]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(addr[6]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(addr[7]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(addr[8]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(addr[9]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(dataBusOut[0]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(dataBusOut[10]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(dataBusOut[11]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(dataBusOut[12]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(dataBusOut[13]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(dataBusOut[14]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(dataBusOut[15]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(dataBusOut[16]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(dataBusOut[17]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(dataBusOut[18]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(dataBusOut[19]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(dataBusOut[1]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(dataBusOut[20]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(dataBusOut[21]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(dataBusOut[22]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(dataBusOut[23]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(dataBusOut[24]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(dataBusOut[25]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(dataBusOut[26]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(dataBusOut[27]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(dataBusOut[28]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(dataBusOut[29]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(dataBusOut[2]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(dataBusOut[30]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(dataBusOut[31]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(dataBusOut[3]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(dataBusOut[4]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(dataBusOut[5]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(dataBusOut[6]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(dataBusOut[7]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(dataBusOut[8]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(dataBusOut[9]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(pc[0]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(pc[10]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(pc[11]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(pc[12]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(pc[13]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(pc[14]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(pc[15]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(pc[16]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(pc[17]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(pc[18]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(pc[19]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(pc[1]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(pc[20]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(pc[21]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(pc[22]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(pc[23]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(pc[24]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(pc[25]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(pc[26]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(pc[27]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(pc[28]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(pc[29]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(pc[2]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(pc[30]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(pc[31]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(pc[3]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(pc[4]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(pc[5]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(pc[6]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(pc[7]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(pc[8]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(pc[9]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(rdEn));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(wrEn));
 sky130_fd_sc_hd__buf_2 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 fanout170 (.A(_04049_),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 fanout171 (.A(net173),
    .X(net171));
 sky130_fd_sc_hd__buf_1 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__buf_2 fanout173 (.A(_04048_),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_4 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_4 fanout175 (.A(net176),
    .X(net175));
 sky130_fd_sc_hd__buf_2 fanout176 (.A(_04045_),
    .X(net176));
 sky130_fd_sc_hd__buf_2 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_4 fanout178 (.A(_04045_),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 wire179 (.A(_04037_),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 wire180 (.A(_05870_),
    .X(net180));
 sky130_fd_sc_hd__buf_2 fanout181 (.A(_02949_),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 max_cap182 (.A(_02906_),
    .X(net182));
 sky130_fd_sc_hd__buf_1 max_cap183 (.A(_02753_),
    .X(net183));
 sky130_fd_sc_hd__buf_2 fanout184 (.A(_05456_),
    .X(net184));
 sky130_fd_sc_hd__buf_2 fanout185 (.A(_03507_),
    .X(net185));
 sky130_fd_sc_hd__buf_2 fanout186 (.A(_03178_),
    .X(net186));
 sky130_fd_sc_hd__buf_2 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_2 fanout188 (.A(net189),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 fanout189 (.A(_02694_),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(_02693_),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_4 fanout191 (.A(net193),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_4 fanout193 (.A(_02647_),
    .X(net193));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(_02646_),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 fanout195 (.A(_02646_),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_4 fanout196 (.A(_02646_),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 fanout197 (.A(_02646_),
    .X(net197));
 sky130_fd_sc_hd__buf_2 fanout198 (.A(_02589_),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 fanout199 (.A(_02589_),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_4 fanout200 (.A(_05453_),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_4 fanout201 (.A(_05453_),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_4 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__buf_2 fanout203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(_05452_),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_2 max_cap205 (.A(_02988_),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_4 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_2 fanout207 (.A(_02723_),
    .X(net207));
 sky130_fd_sc_hd__buf_2 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_4 fanout209 (.A(_02723_),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_4 fanout210 (.A(net215),
    .X(net210));
 sky130_fd_sc_hd__buf_2 fanout211 (.A(net214),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_4 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_2 fanout215 (.A(_02722_),
    .X(net215));
 sky130_fd_sc_hd__buf_2 fanout216 (.A(net221),
    .X(net216));
 sky130_fd_sc_hd__buf_2 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__buf_2 fanout218 (.A(net221),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_4 fanout219 (.A(net221),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__buf_2 fanout221 (.A(_02708_),
    .X(net221));
 sky130_fd_sc_hd__buf_2 fanout222 (.A(_02708_),
    .X(net222));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout223 (.A(_02708_),
    .X(net223));
 sky130_fd_sc_hd__buf_2 fanout224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__buf_2 fanout225 (.A(_02708_),
    .X(net225));
 sky130_fd_sc_hd__buf_2 fanout226 (.A(_02707_),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_4 fanout227 (.A(_02707_),
    .X(net227));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout228 (.A(_02707_),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 fanout229 (.A(net230),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 fanout230 (.A(net232),
    .X(net230));
 sky130_fd_sc_hd__buf_2 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__buf_2 fanout232 (.A(_02690_),
    .X(net232));
 sky130_fd_sc_hd__buf_2 fanout233 (.A(net235),
    .X(net233));
 sky130_fd_sc_hd__buf_2 fanout234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 fanout235 (.A(_02689_),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_4 fanout236 (.A(net238),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 fanout237 (.A(net238),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 fanout238 (.A(net244),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__buf_2 fanout240 (.A(net244),
    .X(net240));
 sky130_fd_sc_hd__buf_2 fanout241 (.A(net244),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 fanout242 (.A(net244),
    .X(net242));
 sky130_fd_sc_hd__buf_2 fanout243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__buf_2 fanout244 (.A(_02683_),
    .X(net244));
 sky130_fd_sc_hd__buf_2 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__buf_2 fanout246 (.A(_02682_),
    .X(net246));
 sky130_fd_sc_hd__buf_2 fanout247 (.A(_02682_),
    .X(net247));
 sky130_fd_sc_hd__buf_2 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 fanout249 (.A(_02682_),
    .X(net249));
 sky130_fd_sc_hd__buf_2 fanout250 (.A(net254),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_2 fanout251 (.A(net254),
    .X(net251));
 sky130_fd_sc_hd__buf_2 fanout252 (.A(net254),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 fanout253 (.A(net254),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_2 fanout254 (.A(net264),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_4 fanout255 (.A(net258),
    .X(net255));
 sky130_fd_sc_hd__buf_2 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__buf_2 fanout257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__buf_2 fanout258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 fanout259 (.A(net264),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_4 fanout260 (.A(net264),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_4 fanout261 (.A(net263),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_2 fanout262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__buf_2 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_4 fanout264 (.A(\brancher.stall ),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_4 fanout265 (.A(_03184_),
    .X(net265));
 sky130_fd_sc_hd__buf_2 fanout266 (.A(net268),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_2 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_4 fanout268 (.A(_01251_),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_8 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__buf_4 fanout270 (.A(_05406_),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_8 fanout271 (.A(net272),
    .X(net271));
 sky130_fd_sc_hd__buf_4 fanout272 (.A(_05406_),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_8 fanout273 (.A(net274),
    .X(net273));
 sky130_fd_sc_hd__buf_4 fanout274 (.A(_05373_),
    .X(net274));
 sky130_fd_sc_hd__buf_4 fanout275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__buf_4 fanout276 (.A(_05373_),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_8 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__buf_4 fanout278 (.A(_05340_),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_8 fanout279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__buf_4 fanout280 (.A(_05340_),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_8 fanout281 (.A(_05307_),
    .X(net281));
 sky130_fd_sc_hd__buf_2 fanout282 (.A(_05307_),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_8 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_8 fanout284 (.A(_05307_),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_8 fanout285 (.A(_05274_),
    .X(net285));
 sky130_fd_sc_hd__buf_2 fanout286 (.A(_05274_),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_8 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_8 fanout288 (.A(_05274_),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_8 fanout289 (.A(_05241_),
    .X(net289));
 sky130_fd_sc_hd__buf_2 fanout290 (.A(_05241_),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_8 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_8 fanout292 (.A(_05241_),
    .X(net292));
 sky130_fd_sc_hd__buf_4 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__buf_4 fanout294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__buf_4 fanout295 (.A(_05208_),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_4 fanout296 (.A(net298),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_4 fanout297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_4 fanout298 (.A(net299),
    .X(net298));
 sky130_fd_sc_hd__buf_4 fanout299 (.A(_05208_),
    .X(net299));
 sky130_fd_sc_hd__buf_4 fanout300 (.A(net301),
    .X(net300));
 sky130_fd_sc_hd__buf_4 fanout301 (.A(_05175_),
    .X(net301));
 sky130_fd_sc_hd__buf_4 fanout302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__buf_4 fanout303 (.A(_05175_),
    .X(net303));
 sky130_fd_sc_hd__buf_4 fanout304 (.A(net305),
    .X(net304));
 sky130_fd_sc_hd__buf_4 fanout305 (.A(_05142_),
    .X(net305));
 sky130_fd_sc_hd__buf_4 fanout306 (.A(net307),
    .X(net306));
 sky130_fd_sc_hd__buf_4 fanout307 (.A(_05142_),
    .X(net307));
 sky130_fd_sc_hd__buf_4 fanout308 (.A(net309),
    .X(net308));
 sky130_fd_sc_hd__buf_4 fanout309 (.A(_05109_),
    .X(net309));
 sky130_fd_sc_hd__buf_4 fanout310 (.A(net311),
    .X(net310));
 sky130_fd_sc_hd__buf_4 fanout311 (.A(_05109_),
    .X(net311));
 sky130_fd_sc_hd__buf_4 fanout312 (.A(net313),
    .X(net312));
 sky130_fd_sc_hd__buf_4 fanout313 (.A(_05076_),
    .X(net313));
 sky130_fd_sc_hd__buf_4 fanout314 (.A(net315),
    .X(net314));
 sky130_fd_sc_hd__buf_4 fanout315 (.A(_05076_),
    .X(net315));
 sky130_fd_sc_hd__buf_4 fanout316 (.A(net317),
    .X(net316));
 sky130_fd_sc_hd__buf_4 fanout317 (.A(_05043_),
    .X(net317));
 sky130_fd_sc_hd__buf_4 fanout318 (.A(net319),
    .X(net318));
 sky130_fd_sc_hd__buf_4 fanout319 (.A(_05043_),
    .X(net319));
 sky130_fd_sc_hd__buf_4 fanout320 (.A(net321),
    .X(net320));
 sky130_fd_sc_hd__buf_4 fanout321 (.A(_05010_),
    .X(net321));
 sky130_fd_sc_hd__buf_4 fanout322 (.A(net323),
    .X(net322));
 sky130_fd_sc_hd__buf_4 fanout323 (.A(_05010_),
    .X(net323));
 sky130_fd_sc_hd__buf_4 fanout324 (.A(net325),
    .X(net324));
 sky130_fd_sc_hd__buf_4 fanout325 (.A(_04977_),
    .X(net325));
 sky130_fd_sc_hd__buf_4 fanout326 (.A(net327),
    .X(net326));
 sky130_fd_sc_hd__buf_4 fanout327 (.A(_04977_),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_8 fanout328 (.A(_04909_),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_4 fanout329 (.A(_04909_),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_8 fanout330 (.A(net331),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_8 fanout331 (.A(_04909_),
    .X(net331));
 sky130_fd_sc_hd__buf_6 fanout332 (.A(net333),
    .X(net332));
 sky130_fd_sc_hd__buf_4 fanout333 (.A(_04844_),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_8 fanout334 (.A(_04844_),
    .X(net334));
 sky130_fd_sc_hd__buf_2 fanout335 (.A(_04844_),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_8 fanout336 (.A(net337),
    .X(net336));
 sky130_fd_sc_hd__buf_4 fanout337 (.A(_04778_),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_8 fanout338 (.A(_04778_),
    .X(net338));
 sky130_fd_sc_hd__buf_2 fanout339 (.A(_04778_),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_8 fanout340 (.A(net341),
    .X(net340));
 sky130_fd_sc_hd__buf_4 fanout341 (.A(_04712_),
    .X(net341));
 sky130_fd_sc_hd__buf_4 fanout342 (.A(_04712_),
    .X(net342));
 sky130_fd_sc_hd__buf_2 fanout343 (.A(_04712_),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_8 fanout344 (.A(net347),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_8 fanout345 (.A(net346),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_8 fanout346 (.A(net347),
    .X(net346));
 sky130_fd_sc_hd__buf_4 fanout347 (.A(_04646_),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_8 fanout348 (.A(_04580_),
    .X(net348));
 sky130_fd_sc_hd__buf_2 fanout349 (.A(_04580_),
    .X(net349));
 sky130_fd_sc_hd__buf_4 fanout350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_8 fanout351 (.A(_04580_),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_8 fanout352 (.A(net355),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_8 fanout353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_8 fanout354 (.A(net355),
    .X(net354));
 sky130_fd_sc_hd__buf_4 fanout355 (.A(_04514_),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_4 fanout356 (.A(net358),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_4 fanout357 (.A(net358),
    .X(net357));
 sky130_fd_sc_hd__buf_4 fanout358 (.A(_04480_),
    .X(net358));
 sky130_fd_sc_hd__buf_4 fanout359 (.A(net361),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_4 fanout360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_4 fanout361 (.A(net362),
    .X(net361));
 sky130_fd_sc_hd__buf_4 fanout362 (.A(_04480_),
    .X(net362));
 sky130_fd_sc_hd__buf_4 fanout363 (.A(net364),
    .X(net363));
 sky130_fd_sc_hd__buf_4 fanout364 (.A(_04447_),
    .X(net364));
 sky130_fd_sc_hd__buf_4 fanout365 (.A(net366),
    .X(net365));
 sky130_fd_sc_hd__buf_4 fanout366 (.A(_04447_),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_8 fanout367 (.A(net368),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_4 fanout368 (.A(_04382_),
    .X(net368));
 sky130_fd_sc_hd__buf_4 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__buf_4 fanout370 (.A(_04382_),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_8 fanout371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__buf_4 fanout372 (.A(_04348_),
    .X(net372));
 sky130_fd_sc_hd__buf_4 fanout373 (.A(_04348_),
    .X(net373));
 sky130_fd_sc_hd__buf_2 fanout374 (.A(_04348_),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_8 fanout375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__buf_4 fanout376 (.A(_04314_),
    .X(net376));
 sky130_fd_sc_hd__buf_4 fanout377 (.A(net378),
    .X(net377));
 sky130_fd_sc_hd__buf_4 fanout378 (.A(_04314_),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_8 fanout379 (.A(net380),
    .X(net379));
 sky130_fd_sc_hd__buf_4 fanout380 (.A(_04280_),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_8 fanout381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__buf_4 fanout382 (.A(_04280_),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_8 fanout383 (.A(net384),
    .X(net383));
 sky130_fd_sc_hd__buf_4 fanout384 (.A(_04246_),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_8 fanout385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__buf_4 fanout386 (.A(_04246_),
    .X(net386));
 sky130_fd_sc_hd__buf_2 fanout387 (.A(_04243_),
    .X(net387));
 sky130_fd_sc_hd__buf_2 fanout388 (.A(_04241_),
    .X(net388));
 sky130_fd_sc_hd__buf_2 fanout389 (.A(_04239_),
    .X(net389));
 sky130_fd_sc_hd__buf_2 fanout390 (.A(_04237_),
    .X(net390));
 sky130_fd_sc_hd__buf_2 fanout391 (.A(_04235_),
    .X(net391));
 sky130_fd_sc_hd__buf_2 fanout392 (.A(_04233_),
    .X(net392));
 sky130_fd_sc_hd__buf_2 fanout393 (.A(_04231_),
    .X(net393));
 sky130_fd_sc_hd__buf_2 fanout394 (.A(_04229_),
    .X(net394));
 sky130_fd_sc_hd__buf_2 fanout395 (.A(_04227_),
    .X(net395));
 sky130_fd_sc_hd__buf_2 fanout396 (.A(_04225_),
    .X(net396));
 sky130_fd_sc_hd__buf_2 fanout397 (.A(_04223_),
    .X(net397));
 sky130_fd_sc_hd__buf_2 fanout398 (.A(_04221_),
    .X(net398));
 sky130_fd_sc_hd__buf_2 fanout399 (.A(_04219_),
    .X(net399));
 sky130_fd_sc_hd__buf_2 fanout400 (.A(_04217_),
    .X(net400));
 sky130_fd_sc_hd__buf_2 fanout401 (.A(_04215_),
    .X(net401));
 sky130_fd_sc_hd__buf_2 fanout402 (.A(_04213_),
    .X(net402));
 sky130_fd_sc_hd__buf_2 fanout403 (.A(_04211_),
    .X(net403));
 sky130_fd_sc_hd__buf_2 fanout404 (.A(_04209_),
    .X(net404));
 sky130_fd_sc_hd__buf_2 fanout405 (.A(_04207_),
    .X(net405));
 sky130_fd_sc_hd__buf_2 fanout406 (.A(_04205_),
    .X(net406));
 sky130_fd_sc_hd__buf_2 fanout407 (.A(_04203_),
    .X(net407));
 sky130_fd_sc_hd__buf_2 fanout408 (.A(_04201_),
    .X(net408));
 sky130_fd_sc_hd__buf_2 fanout409 (.A(_04199_),
    .X(net409));
 sky130_fd_sc_hd__buf_2 fanout410 (.A(_04197_),
    .X(net410));
 sky130_fd_sc_hd__buf_2 fanout411 (.A(_04195_),
    .X(net411));
 sky130_fd_sc_hd__buf_2 fanout412 (.A(_04193_),
    .X(net412));
 sky130_fd_sc_hd__buf_2 fanout413 (.A(_04191_),
    .X(net413));
 sky130_fd_sc_hd__buf_2 fanout414 (.A(_04189_),
    .X(net414));
 sky130_fd_sc_hd__buf_2 fanout415 (.A(_04187_),
    .X(net415));
 sky130_fd_sc_hd__buf_2 fanout416 (.A(_04185_),
    .X(net416));
 sky130_fd_sc_hd__buf_2 fanout417 (.A(_04183_),
    .X(net417));
 sky130_fd_sc_hd__buf_2 fanout418 (.A(_04181_),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_8 fanout419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__buf_4 fanout420 (.A(_04177_),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_8 fanout421 (.A(net422),
    .X(net421));
 sky130_fd_sc_hd__buf_4 fanout422 (.A(_04177_),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_4 fanout423 (.A(net425),
    .X(net423));
 sky130_fd_sc_hd__buf_2 fanout424 (.A(net425),
    .X(net424));
 sky130_fd_sc_hd__buf_2 fanout425 (.A(_03266_),
    .X(net425));
 sky130_fd_sc_hd__buf_2 fanout426 (.A(_03260_),
    .X(net426));
 sky130_fd_sc_hd__clkbuf_2 fanout427 (.A(_03260_),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_4 fanout428 (.A(_03259_),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_2 fanout429 (.A(_03259_),
    .X(net429));
 sky130_fd_sc_hd__buf_4 fanout430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_4 fanout431 (.A(_03182_),
    .X(net431));
 sky130_fd_sc_hd__clkbuf_1 max_cap432 (.A(_05995_),
    .X(net432));
 sky130_fd_sc_hd__buf_2 fanout433 (.A(net436),
    .X(net433));
 sky130_fd_sc_hd__buf_2 fanout434 (.A(net436),
    .X(net434));
 sky130_fd_sc_hd__buf_2 fanout435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__buf_2 fanout436 (.A(net442),
    .X(net436));
 sky130_fd_sc_hd__buf_2 fanout437 (.A(net442),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_2 fanout438 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_4 fanout439 (.A(net442),
    .X(net439));
 sky130_fd_sc_hd__buf_2 fanout440 (.A(net442),
    .X(net440));
 sky130_fd_sc_hd__buf_2 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_2 fanout442 (.A(net488),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_4 fanout443 (.A(net451),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_2 fanout444 (.A(net451),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_4 fanout445 (.A(net451),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_2 fanout446 (.A(net451),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_4 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_4 fanout448 (.A(net451),
    .X(net448));
 sky130_fd_sc_hd__buf_2 fanout449 (.A(net451),
    .X(net449));
 sky130_fd_sc_hd__buf_2 fanout450 (.A(net451),
    .X(net450));
 sky130_fd_sc_hd__buf_2 fanout451 (.A(net488),
    .X(net451));
 sky130_fd_sc_hd__clkbuf_4 fanout452 (.A(net454),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_4 fanout453 (.A(net454),
    .X(net453));
 sky130_fd_sc_hd__clkbuf_4 fanout454 (.A(net459),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_4 fanout455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__buf_2 fanout456 (.A(net458),
    .X(net456));
 sky130_fd_sc_hd__buf_4 fanout457 (.A(net458),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_2 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__buf_2 fanout459 (.A(net488),
    .X(net459));
 sky130_fd_sc_hd__buf_2 fanout460 (.A(net461),
    .X(net460));
 sky130_fd_sc_hd__buf_2 fanout461 (.A(net469),
    .X(net461));
 sky130_fd_sc_hd__buf_2 fanout462 (.A(net464),
    .X(net462));
 sky130_fd_sc_hd__buf_2 fanout463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_2 fanout464 (.A(net469),
    .X(net464));
 sky130_fd_sc_hd__buf_2 fanout465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_4 fanout466 (.A(net469),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_4 fanout467 (.A(net469),
    .X(net467));
 sky130_fd_sc_hd__clkbuf_2 fanout468 (.A(net469),
    .X(net468));
 sky130_fd_sc_hd__buf_2 fanout469 (.A(net488),
    .X(net469));
 sky130_fd_sc_hd__buf_2 fanout470 (.A(net472),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_2 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_4 fanout472 (.A(net474),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_4 fanout473 (.A(net474),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_2 fanout474 (.A(net488),
    .X(net474));
 sky130_fd_sc_hd__buf_2 fanout475 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_4 fanout476 (.A(net479),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_4 fanout477 (.A(net479),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_2 fanout478 (.A(net479),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_2 fanout479 (.A(net488),
    .X(net479));
 sky130_fd_sc_hd__clkbuf_4 fanout480 (.A(net487),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_2 fanout481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__buf_2 fanout482 (.A(net487),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_4 fanout483 (.A(net486),
    .X(net483));
 sky130_fd_sc_hd__buf_2 fanout484 (.A(net486),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_4 fanout485 (.A(net486),
    .X(net485));
 sky130_fd_sc_hd__buf_2 fanout486 (.A(net487),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_4 fanout487 (.A(net488),
    .X(net487));
 sky130_fd_sc_hd__buf_4 fanout488 (.A(_04975_),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_8 fanout489 (.A(net490),
    .X(net489));
 sky130_fd_sc_hd__buf_4 fanout490 (.A(_04942_),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_8 fanout491 (.A(net492),
    .X(net491));
 sky130_fd_sc_hd__buf_4 fanout492 (.A(_04942_),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_8 fanout493 (.A(net494),
    .X(net493));
 sky130_fd_sc_hd__buf_4 fanout494 (.A(_04777_),
    .X(net494));
 sky130_fd_sc_hd__buf_4 fanout495 (.A(net496),
    .X(net495));
 sky130_fd_sc_hd__buf_4 fanout496 (.A(_04777_),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_8 fanout497 (.A(_04711_),
    .X(net497));
 sky130_fd_sc_hd__buf_4 fanout498 (.A(_04711_),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_8 fanout499 (.A(net500),
    .X(net499));
 sky130_fd_sc_hd__buf_4 fanout500 (.A(_04711_),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_8 fanout501 (.A(_04513_),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_4 fanout502 (.A(_04513_),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_8 fanout503 (.A(net504),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_8 fanout504 (.A(_04513_),
    .X(net504));
 sky130_fd_sc_hd__buf_4 fanout505 (.A(net506),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_4 fanout506 (.A(_04180_),
    .X(net506));
 sky130_fd_sc_hd__buf_4 fanout507 (.A(net508),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_4 fanout508 (.A(_04180_),
    .X(net508));
 sky130_fd_sc_hd__buf_2 fanout509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_2 fanout510 (.A(net517),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_4 fanout511 (.A(net517),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_2 fanout512 (.A(net517),
    .X(net512));
 sky130_fd_sc_hd__buf_2 fanout513 (.A(net517),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_2 fanout514 (.A(net517),
    .X(net514));
 sky130_fd_sc_hd__buf_2 fanout515 (.A(net517),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_2 fanout516 (.A(net517),
    .X(net516));
 sky130_fd_sc_hd__buf_2 fanout517 (.A(net528),
    .X(net517));
 sky130_fd_sc_hd__buf_2 fanout518 (.A(net519),
    .X(net518));
 sky130_fd_sc_hd__buf_2 fanout519 (.A(net523),
    .X(net519));
 sky130_fd_sc_hd__buf_2 fanout520 (.A(net522),
    .X(net520));
 sky130_fd_sc_hd__buf_2 fanout521 (.A(net522),
    .X(net521));
 sky130_fd_sc_hd__clkbuf_2 fanout522 (.A(net523),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_2 fanout523 (.A(net528),
    .X(net523));
 sky130_fd_sc_hd__buf_2 fanout524 (.A(net528),
    .X(net524));
 sky130_fd_sc_hd__clkbuf_2 fanout525 (.A(net528),
    .X(net525));
 sky130_fd_sc_hd__buf_2 fanout526 (.A(net527),
    .X(net526));
 sky130_fd_sc_hd__buf_2 fanout527 (.A(net528),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_2 fanout528 (.A(net537),
    .X(net528));
 sky130_fd_sc_hd__buf_2 fanout529 (.A(net531),
    .X(net529));
 sky130_fd_sc_hd__buf_2 fanout530 (.A(net531),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_2 fanout531 (.A(net532),
    .X(net531));
 sky130_fd_sc_hd__buf_2 fanout532 (.A(net537),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_4 fanout533 (.A(net535),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_2 fanout534 (.A(net535),
    .X(net534));
 sky130_fd_sc_hd__buf_2 fanout535 (.A(net536),
    .X(net535));
 sky130_fd_sc_hd__clkbuf_8 fanout536 (.A(net537),
    .X(net536));
 sky130_fd_sc_hd__buf_2 fanout537 (.A(_04174_),
    .X(net537));
 sky130_fd_sc_hd__buf_2 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_4 fanout539 (.A(net542),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_4 fanout540 (.A(net542),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_2 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_2 fanout542 (.A(net556),
    .X(net542));
 sky130_fd_sc_hd__buf_2 fanout543 (.A(net556),
    .X(net543));
 sky130_fd_sc_hd__buf_2 fanout544 (.A(net556),
    .X(net544));
 sky130_fd_sc_hd__buf_2 fanout545 (.A(net546),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_4 fanout546 (.A(net556),
    .X(net546));
 sky130_fd_sc_hd__buf_2 fanout547 (.A(net548),
    .X(net547));
 sky130_fd_sc_hd__buf_2 fanout548 (.A(net555),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_4 fanout549 (.A(net555),
    .X(net549));
 sky130_fd_sc_hd__buf_2 fanout550 (.A(net555),
    .X(net550));
 sky130_fd_sc_hd__buf_2 fanout551 (.A(net555),
    .X(net551));
 sky130_fd_sc_hd__buf_2 fanout552 (.A(net554),
    .X(net552));
 sky130_fd_sc_hd__clkbuf_2 fanout553 (.A(net554),
    .X(net553));
 sky130_fd_sc_hd__buf_2 fanout554 (.A(net555),
    .X(net554));
 sky130_fd_sc_hd__buf_2 fanout555 (.A(net556),
    .X(net555));
 sky130_fd_sc_hd__buf_2 fanout556 (.A(_04174_),
    .X(net556));
 sky130_fd_sc_hd__buf_2 fanout557 (.A(net564),
    .X(net557));
 sky130_fd_sc_hd__buf_2 fanout558 (.A(net564),
    .X(net558));
 sky130_fd_sc_hd__buf_2 fanout559 (.A(net563),
    .X(net559));
 sky130_fd_sc_hd__buf_2 fanout560 (.A(net562),
    .X(net560));
 sky130_fd_sc_hd__buf_2 fanout561 (.A(net562),
    .X(net561));
 sky130_fd_sc_hd__buf_2 fanout562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_2 fanout563 (.A(net564),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_2 fanout564 (.A(net565),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_4 fanout565 (.A(_04174_),
    .X(net565));
 sky130_fd_sc_hd__clkbuf_4 fanout566 (.A(net567),
    .X(net566));
 sky130_fd_sc_hd__buf_2 fanout567 (.A(_03219_),
    .X(net567));
 sky130_fd_sc_hd__buf_2 fanout568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__buf_2 fanout569 (.A(_03219_),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_4 fanout570 (.A(net572),
    .X(net570));
 sky130_fd_sc_hd__buf_1 fanout571 (.A(net572),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_4 fanout572 (.A(_03169_),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_4 fanout573 (.A(_03138_),
    .X(net573));
 sky130_fd_sc_hd__clkbuf_4 fanout574 (.A(_02585_),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_4 fanout575 (.A(net582),
    .X(net575));
 sky130_fd_sc_hd__buf_2 fanout576 (.A(net582),
    .X(net576));
 sky130_fd_sc_hd__buf_4 fanout577 (.A(net582),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_4 fanout578 (.A(net579),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_4 fanout579 (.A(net582),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_4 fanout580 (.A(net581),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_4 fanout581 (.A(net582),
    .X(net581));
 sky130_fd_sc_hd__buf_4 fanout582 (.A(_01986_),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_8 fanout583 (.A(net584),
    .X(net583));
 sky130_fd_sc_hd__buf_4 fanout584 (.A(_01985_),
    .X(net584));
 sky130_fd_sc_hd__buf_4 fanout585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__buf_4 fanout586 (.A(_01985_),
    .X(net586));
 sky130_fd_sc_hd__buf_2 fanout587 (.A(net588),
    .X(net587));
 sky130_fd_sc_hd__buf_2 fanout588 (.A(net589),
    .X(net588));
 sky130_fd_sc_hd__buf_2 fanout589 (.A(_01264_),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_4 fanout590 (.A(net592),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_2 fanout591 (.A(net592),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_2 fanout592 (.A(net593),
    .X(net592));
 sky130_fd_sc_hd__buf_2 fanout593 (.A(net594),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_4 fanout594 (.A(_01264_),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_4 fanout595 (.A(net597),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_4 fanout596 (.A(net597),
    .X(net596));
 sky130_fd_sc_hd__buf_2 fanout597 (.A(net600),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_4 fanout598 (.A(net599),
    .X(net598));
 sky130_fd_sc_hd__buf_4 fanout599 (.A(net600),
    .X(net599));
 sky130_fd_sc_hd__buf_4 fanout600 (.A(_01263_),
    .X(net600));
 sky130_fd_sc_hd__buf_4 fanout601 (.A(net604),
    .X(net601));
 sky130_fd_sc_hd__buf_4 fanout602 (.A(net603),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_4 fanout603 (.A(net604),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_4 fanout604 (.A(_01250_),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_4 fanout605 (.A(net608),
    .X(net605));
 sky130_fd_sc_hd__buf_2 fanout606 (.A(net608),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_4 fanout607 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_4 fanout608 (.A(_01250_),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_4 fanout609 (.A(net611),
    .X(net609));
 sky130_fd_sc_hd__buf_4 fanout610 (.A(net611),
    .X(net610));
 sky130_fd_sc_hd__buf_4 fanout611 (.A(_01249_),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_4 fanout612 (.A(net615),
    .X(net612));
 sky130_fd_sc_hd__clkbuf_4 fanout613 (.A(net615),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_4 fanout614 (.A(net615),
    .X(net614));
 sky130_fd_sc_hd__buf_4 fanout615 (.A(_01249_),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_4 fanout616 (.A(net618),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_4 fanout617 (.A(net618),
    .X(net617));
 sky130_fd_sc_hd__clkbuf_4 fanout618 (.A(_01238_),
    .X(net618));
 sky130_fd_sc_hd__buf_2 fanout619 (.A(net621),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_4 fanout620 (.A(net621),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_4 fanout621 (.A(_01238_),
    .X(net621));
 sky130_fd_sc_hd__clkbuf_4 fanout622 (.A(net623),
    .X(net622));
 sky130_fd_sc_hd__buf_4 fanout623 (.A(_01237_),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_2 fanout624 (.A(_01237_),
    .X(net624));
 sky130_fd_sc_hd__buf_2 fanout625 (.A(net626),
    .X(net625));
 sky130_fd_sc_hd__buf_2 fanout626 (.A(net627),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_4 fanout627 (.A(_01237_),
    .X(net627));
 sky130_fd_sc_hd__buf_4 fanout628 (.A(_05455_),
    .X(net628));
 sky130_fd_sc_hd__buf_2 fanout629 (.A(_05455_),
    .X(net629));
 sky130_fd_sc_hd__buf_4 fanout630 (.A(_05454_),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_8 fanout631 (.A(net632),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_8 fanout632 (.A(_04843_),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_8 fanout633 (.A(net634),
    .X(net633));
 sky130_fd_sc_hd__buf_4 fanout634 (.A(_04843_),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_8 fanout635 (.A(_04645_),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_4 fanout636 (.A(_04645_),
    .X(net636));
 sky130_fd_sc_hd__buf_4 fanout637 (.A(net638),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_8 fanout638 (.A(_04645_),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_8 fanout639 (.A(_04579_),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_4 fanout640 (.A(_04579_),
    .X(net640));
 sky130_fd_sc_hd__buf_4 fanout641 (.A(net642),
    .X(net641));
 sky130_fd_sc_hd__clkbuf_8 fanout642 (.A(_04579_),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_8 fanout643 (.A(net644),
    .X(net643));
 sky130_fd_sc_hd__buf_4 fanout644 (.A(_04381_),
    .X(net644));
 sky130_fd_sc_hd__clkbuf_8 fanout645 (.A(net646),
    .X(net645));
 sky130_fd_sc_hd__buf_4 fanout646 (.A(_04381_),
    .X(net646));
 sky130_fd_sc_hd__buf_4 fanout647 (.A(net649),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_4 fanout648 (.A(net649),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_4 fanout649 (.A(net654),
    .X(net649));
 sky130_fd_sc_hd__buf_4 fanout650 (.A(net654),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_4 fanout651 (.A(net653),
    .X(net651));
 sky130_fd_sc_hd__clkbuf_4 fanout652 (.A(net653),
    .X(net652));
 sky130_fd_sc_hd__buf_4 fanout653 (.A(net654),
    .X(net653));
 sky130_fd_sc_hd__buf_4 fanout654 (.A(_04347_),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_4 fanout655 (.A(net657),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_4 fanout656 (.A(net657),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_4 fanout657 (.A(net658),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_8 fanout658 (.A(_04313_),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_4 fanout659 (.A(net661),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_4 fanout660 (.A(net661),
    .X(net660));
 sky130_fd_sc_hd__buf_2 fanout661 (.A(net662),
    .X(net661));
 sky130_fd_sc_hd__buf_4 fanout662 (.A(_04313_),
    .X(net662));
 sky130_fd_sc_hd__buf_4 fanout663 (.A(net665),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_4 fanout664 (.A(net665),
    .X(net664));
 sky130_fd_sc_hd__clkbuf_4 fanout665 (.A(net666),
    .X(net665));
 sky130_fd_sc_hd__buf_4 fanout666 (.A(_04279_),
    .X(net666));
 sky130_fd_sc_hd__buf_4 fanout667 (.A(net668),
    .X(net667));
 sky130_fd_sc_hd__buf_4 fanout668 (.A(net670),
    .X(net668));
 sky130_fd_sc_hd__buf_4 fanout669 (.A(net670),
    .X(net669));
 sky130_fd_sc_hd__clkbuf_4 fanout670 (.A(_04279_),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_4 fanout671 (.A(net673),
    .X(net671));
 sky130_fd_sc_hd__clkbuf_4 fanout672 (.A(net679),
    .X(net672));
 sky130_fd_sc_hd__buf_2 fanout673 (.A(net679),
    .X(net673));
 sky130_fd_sc_hd__clkbuf_8 fanout674 (.A(net679),
    .X(net674));
 sky130_fd_sc_hd__clkbuf_4 fanout675 (.A(net678),
    .X(net675));
 sky130_fd_sc_hd__buf_4 fanout676 (.A(net678),
    .X(net676));
 sky130_fd_sc_hd__buf_4 fanout677 (.A(net678),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_4 fanout678 (.A(net679),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_4 fanout679 (.A(_04176_),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_4 fanout680 (.A(net682),
    .X(net680));
 sky130_fd_sc_hd__clkbuf_4 fanout681 (.A(net683),
    .X(net681));
 sky130_fd_sc_hd__clkbuf_2 fanout682 (.A(net683),
    .X(net682));
 sky130_fd_sc_hd__buf_4 fanout683 (.A(net687),
    .X(net683));
 sky130_fd_sc_hd__clkbuf_4 fanout684 (.A(net685),
    .X(net684));
 sky130_fd_sc_hd__buf_4 fanout685 (.A(net686),
    .X(net685));
 sky130_fd_sc_hd__buf_4 fanout686 (.A(net687),
    .X(net686));
 sky130_fd_sc_hd__buf_4 fanout687 (.A(_04140_),
    .X(net687));
 sky130_fd_sc_hd__buf_2 fanout688 (.A(_03131_),
    .X(net688));
 sky130_fd_sc_hd__buf_2 fanout689 (.A(_03077_),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_4 fanout690 (.A(_03061_),
    .X(net690));
 sky130_fd_sc_hd__buf_2 fanout691 (.A(_03044_),
    .X(net691));
 sky130_fd_sc_hd__buf_2 fanout692 (.A(_03030_),
    .X(net692));
 sky130_fd_sc_hd__buf_2 fanout693 (.A(_03014_),
    .X(net693));
 sky130_fd_sc_hd__buf_2 fanout694 (.A(_03000_),
    .X(net694));
 sky130_fd_sc_hd__buf_2 fanout695 (.A(_02984_),
    .X(net695));
 sky130_fd_sc_hd__clkbuf_4 fanout696 (.A(_02969_),
    .X(net696));
 sky130_fd_sc_hd__buf_2 fanout697 (.A(_02951_),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_4 fanout698 (.A(_02938_),
    .X(net698));
 sky130_fd_sc_hd__buf_2 fanout699 (.A(_02923_),
    .X(net699));
 sky130_fd_sc_hd__buf_2 fanout700 (.A(_02909_),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_4 fanout701 (.A(_02894_),
    .X(net701));
 sky130_fd_sc_hd__buf_2 fanout702 (.A(_02881_),
    .X(net702));
 sky130_fd_sc_hd__buf_2 fanout703 (.A(_02864_),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_4 fanout704 (.A(_02850_),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_4 fanout705 (.A(_02832_),
    .X(net705));
 sky130_fd_sc_hd__buf_2 fanout706 (.A(_02816_),
    .X(net706));
 sky130_fd_sc_hd__buf_2 fanout707 (.A(_02800_),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_4 fanout708 (.A(_02786_),
    .X(net708));
 sky130_fd_sc_hd__buf_2 fanout709 (.A(_02770_),
    .X(net709));
 sky130_fd_sc_hd__buf_2 fanout710 (.A(_02756_),
    .X(net710));
 sky130_fd_sc_hd__buf_2 fanout711 (.A(_02742_),
    .X(net711));
 sky130_fd_sc_hd__buf_2 fanout712 (.A(_02717_),
    .X(net712));
 sky130_fd_sc_hd__buf_2 fanout713 (.A(_02703_),
    .X(net713));
 sky130_fd_sc_hd__clkbuf_2 fanout714 (.A(net715),
    .X(net714));
 sky130_fd_sc_hd__clkbuf_2 fanout715 (.A(net717),
    .X(net715));
 sky130_fd_sc_hd__buf_2 fanout716 (.A(net717),
    .X(net716));
 sky130_fd_sc_hd__buf_2 fanout717 (.A(_02692_),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_4 fanout718 (.A(net720),
    .X(net718));
 sky130_fd_sc_hd__buf_2 fanout719 (.A(net720),
    .X(net719));
 sky130_fd_sc_hd__clkbuf_2 fanout720 (.A(_02691_),
    .X(net720));
 sky130_fd_sc_hd__buf_2 fanout721 (.A(_02673_),
    .X(net721));
 sky130_fd_sc_hd__buf_2 fanout722 (.A(_02654_),
    .X(net722));
 sky130_fd_sc_hd__clkbuf_4 fanout723 (.A(_02642_),
    .X(net723));
 sky130_fd_sc_hd__buf_2 fanout724 (.A(_02623_),
    .X(net724));
 sky130_fd_sc_hd__buf_2 fanout725 (.A(_02604_),
    .X(net725));
 sky130_fd_sc_hd__buf_2 fanout726 (.A(net727),
    .X(net726));
 sky130_fd_sc_hd__buf_2 fanout727 (.A(_02590_),
    .X(net727));
 sky130_fd_sc_hd__clkbuf_8 fanout728 (.A(net729),
    .X(net728));
 sky130_fd_sc_hd__buf_4 fanout729 (.A(net730),
    .X(net729));
 sky130_fd_sc_hd__clkbuf_8 fanout730 (.A(_02581_),
    .X(net730));
 sky130_fd_sc_hd__clkbuf_8 fanout731 (.A(net732),
    .X(net731));
 sky130_fd_sc_hd__buf_4 fanout732 (.A(net733),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_4 fanout733 (.A(_02581_),
    .X(net733));
 sky130_fd_sc_hd__buf_4 fanout734 (.A(net736),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_4 fanout735 (.A(net736),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_8 fanout736 (.A(net739),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_8 fanout737 (.A(net738),
    .X(net737));
 sky130_fd_sc_hd__buf_4 fanout738 (.A(net739),
    .X(net738));
 sky130_fd_sc_hd__buf_4 fanout739 (.A(_02580_),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_4 fanout740 (.A(net742),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_4 fanout741 (.A(net742),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_4 fanout742 (.A(_02576_),
    .X(net742));
 sky130_fd_sc_hd__buf_2 wire743 (.A(_02575_),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_1 max_cap744 (.A(_01259_),
    .X(net744));
 sky130_fd_sc_hd__buf_4 fanout745 (.A(net747),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_4 fanout746 (.A(net747),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_4 fanout747 (.A(net748),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_8 fanout748 (.A(_04245_),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_4 fanout749 (.A(net750),
    .X(net749));
 sky130_fd_sc_hd__buf_4 fanout750 (.A(net752),
    .X(net750));
 sky130_fd_sc_hd__buf_4 fanout751 (.A(net752),
    .X(net751));
 sky130_fd_sc_hd__buf_4 fanout752 (.A(_04245_),
    .X(net752));
 sky130_fd_sc_hd__buf_2 fanout753 (.A(net755),
    .X(net753));
 sky130_fd_sc_hd__buf_2 fanout754 (.A(net755),
    .X(net754));
 sky130_fd_sc_hd__buf_2 fanout755 (.A(net756),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_4 fanout756 (.A(_04050_),
    .X(net756));
 sky130_fd_sc_hd__buf_2 fanout757 (.A(_03612_),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_4 fanout758 (.A(_02578_),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_4 fanout759 (.A(_02578_),
    .X(net759));
 sky130_fd_sc_hd__buf_4 fanout760 (.A(net761),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_4 fanout761 (.A(_02577_),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_4 fanout762 (.A(net763),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_4 fanout763 (.A(_02577_),
    .X(net763));
 sky130_fd_sc_hd__buf_4 fanout764 (.A(_02574_),
    .X(net764));
 sky130_fd_sc_hd__clkbuf_2 fanout765 (.A(_02574_),
    .X(net765));
 sky130_fd_sc_hd__buf_2 fanout766 (.A(net770),
    .X(net766));
 sky130_fd_sc_hd__buf_2 fanout767 (.A(net769),
    .X(net767));
 sky130_fd_sc_hd__buf_2 fanout768 (.A(net769),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_2 fanout769 (.A(net770),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_2 fanout770 (.A(_02573_),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_2 fanout771 (.A(net772),
    .X(net771));
 sky130_fd_sc_hd__buf_4 fanout772 (.A(_01285_),
    .X(net772));
 sky130_fd_sc_hd__buf_4 fanout773 (.A(_01284_),
    .X(net773));
 sky130_fd_sc_hd__clkbuf_4 fanout774 (.A(net776),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_4 fanout775 (.A(net776),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_4 fanout776 (.A(net777),
    .X(net776));
 sky130_fd_sc_hd__buf_4 fanout777 (.A(_01253_),
    .X(net777));
 sky130_fd_sc_hd__buf_4 fanout778 (.A(net780),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_4 fanout779 (.A(net780),
    .X(net779));
 sky130_fd_sc_hd__buf_2 fanout780 (.A(net781),
    .X(net780));
 sky130_fd_sc_hd__buf_4 fanout781 (.A(net782),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_2 max_cap782 (.A(_01253_),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_8 fanout783 (.A(net784),
    .X(net783));
 sky130_fd_sc_hd__buf_4 fanout784 (.A(_01222_),
    .X(net784));
 sky130_fd_sc_hd__buf_4 fanout785 (.A(net786),
    .X(net785));
 sky130_fd_sc_hd__buf_4 fanout786 (.A(_01222_),
    .X(net786));
 sky130_fd_sc_hd__buf_4 fanout787 (.A(net789),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_2 fanout788 (.A(net789),
    .X(net788));
 sky130_fd_sc_hd__buf_4 fanout789 (.A(net790),
    .X(net789));
 sky130_fd_sc_hd__buf_4 fanout790 (.A(net794),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_4 fanout791 (.A(net793),
    .X(net791));
 sky130_fd_sc_hd__buf_4 fanout792 (.A(net793),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_8 fanout793 (.A(net794),
    .X(net793));
 sky130_fd_sc_hd__buf_8 fanout794 (.A(_01221_),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_4 fanout795 (.A(net798),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_2 fanout796 (.A(net798),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_4 fanout797 (.A(net798),
    .X(net797));
 sky130_fd_sc_hd__clkbuf_2 fanout798 (.A(net803),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_4 fanout799 (.A(net803),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_4 fanout800 (.A(net803),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_4 fanout801 (.A(net803),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_2 fanout802 (.A(net803),
    .X(net802));
 sky130_fd_sc_hd__buf_4 fanout803 (.A(_01220_),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_4 fanout804 (.A(net806),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_2 fanout805 (.A(net806),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_4 fanout806 (.A(net811),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_4 fanout807 (.A(net808),
    .X(net807));
 sky130_fd_sc_hd__buf_4 fanout808 (.A(net811),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_4 fanout809 (.A(net810),
    .X(net809));
 sky130_fd_sc_hd__buf_4 fanout810 (.A(net811),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_4 fanout811 (.A(_01220_),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_4 fanout812 (.A(_01219_),
    .X(net812));
 sky130_fd_sc_hd__clkbuf_4 fanout813 (.A(_01217_),
    .X(net813));
 sky130_fd_sc_hd__buf_4 fanout814 (.A(net815),
    .X(net814));
 sky130_fd_sc_hd__buf_4 fanout815 (.A(_01212_),
    .X(net815));
 sky130_fd_sc_hd__buf_4 fanout816 (.A(net817),
    .X(net816));
 sky130_fd_sc_hd__buf_4 fanout817 (.A(_01212_),
    .X(net817));
 sky130_fd_sc_hd__buf_4 fanout818 (.A(net820),
    .X(net818));
 sky130_fd_sc_hd__buf_2 fanout819 (.A(net820),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_4 fanout820 (.A(_01211_),
    .X(net820));
 sky130_fd_sc_hd__buf_4 fanout821 (.A(net822),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_8 fanout822 (.A(_01211_),
    .X(net822));
 sky130_fd_sc_hd__buf_4 fanout823 (.A(net828),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_4 fanout824 (.A(net828),
    .X(net824));
 sky130_fd_sc_hd__buf_4 fanout825 (.A(net828),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_4 fanout826 (.A(net828),
    .X(net826));
 sky130_fd_sc_hd__buf_4 fanout827 (.A(net828),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_4 fanout828 (.A(_01210_),
    .X(net828));
 sky130_fd_sc_hd__buf_4 fanout829 (.A(net835),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_2 fanout830 (.A(net835),
    .X(net830));
 sky130_fd_sc_hd__buf_4 fanout831 (.A(net832),
    .X(net831));
 sky130_fd_sc_hd__buf_4 fanout832 (.A(net835),
    .X(net832));
 sky130_fd_sc_hd__buf_4 fanout833 (.A(net835),
    .X(net833));
 sky130_fd_sc_hd__clkbuf_2 fanout834 (.A(net835),
    .X(net834));
 sky130_fd_sc_hd__buf_4 fanout835 (.A(_01210_),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_4 fanout836 (.A(net839),
    .X(net836));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout837 (.A(net839),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_4 fanout838 (.A(net839),
    .X(net838));
 sky130_fd_sc_hd__buf_2 fanout839 (.A(_01207_),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_4 fanout840 (.A(\brancher.imm13_b[12] ),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_4 fanout841 (.A(net843),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_2 fanout842 (.A(net843),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_2 fanout843 (.A(net844),
    .X(net843));
 sky130_fd_sc_hd__buf_2 fanout844 (.A(\brancher.imm13_b[12] ),
    .X(net844));
 sky130_fd_sc_hd__clkbuf_4 fanout845 (.A(net846),
    .X(net845));
 sky130_fd_sc_hd__buf_4 fanout846 (.A(\brancher.funct3[1] ),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_4 fanout847 (.A(\brancher.funct3[0] ),
    .X(net847));
 sky130_fd_sc_hd__buf_4 fanout848 (.A(net850),
    .X(net848));
 sky130_fd_sc_hd__buf_4 fanout849 (.A(net850),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_4 fanout850 (.A(\brancher.imm21_j[3] ),
    .X(net850));
 sky130_fd_sc_hd__clkbuf_4 fanout851 (.A(net852),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_2 fanout852 (.A(\brancher.imm21_j[3] ),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_4 fanout853 (.A(net856),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_4 fanout854 (.A(net856),
    .X(net854));
 sky130_fd_sc_hd__buf_4 fanout855 (.A(net856),
    .X(net855));
 sky130_fd_sc_hd__buf_4 fanout856 (.A(\brancher.imm21_j[3] ),
    .X(net856));
 sky130_fd_sc_hd__buf_4 fanout857 (.A(net859),
    .X(net857));
 sky130_fd_sc_hd__buf_2 fanout858 (.A(net859),
    .X(net858));
 sky130_fd_sc_hd__buf_4 fanout859 (.A(net861),
    .X(net859));
 sky130_fd_sc_hd__buf_4 fanout860 (.A(net861),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_4 fanout861 (.A(\brancher.imm21_j[2] ),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_4 fanout862 (.A(net863),
    .X(net862));
 sky130_fd_sc_hd__buf_4 fanout863 (.A(net864),
    .X(net863));
 sky130_fd_sc_hd__buf_4 fanout864 (.A(\brancher.imm21_j[2] ),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_4 fanout865 (.A(net866),
    .X(net865));
 sky130_fd_sc_hd__clkbuf_4 fanout866 (.A(net870),
    .X(net866));
 sky130_fd_sc_hd__clkbuf_4 fanout867 (.A(net869),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_4 fanout868 (.A(net869),
    .X(net868));
 sky130_fd_sc_hd__buf_2 fanout869 (.A(net870),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_2 fanout870 (.A(net901),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_4 fanout871 (.A(net873),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_4 fanout872 (.A(net873),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_2 fanout873 (.A(net876),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_4 fanout874 (.A(net876),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_4 fanout875 (.A(net876),
    .X(net875));
 sky130_fd_sc_hd__buf_2 fanout876 (.A(net901),
    .X(net876));
 sky130_fd_sc_hd__clkbuf_4 fanout877 (.A(net878),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_4 fanout878 (.A(net881),
    .X(net878));
 sky130_fd_sc_hd__clkbuf_4 fanout879 (.A(net880),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_4 fanout880 (.A(net881),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_2 fanout881 (.A(net882),
    .X(net881));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout882 (.A(net901),
    .X(net882));
 sky130_fd_sc_hd__clkbuf_4 fanout883 (.A(net885),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_4 fanout884 (.A(net885),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_2 fanout885 (.A(net894),
    .X(net885));
 sky130_fd_sc_hd__clkbuf_4 fanout886 (.A(net887),
    .X(net886));
 sky130_fd_sc_hd__clkbuf_4 fanout887 (.A(net894),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_4 fanout888 (.A(net893),
    .X(net888));
 sky130_fd_sc_hd__clkbuf_4 fanout889 (.A(net893),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_4 fanout890 (.A(net892),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_4 fanout891 (.A(net893),
    .X(net891));
 sky130_fd_sc_hd__clkbuf_2 fanout892 (.A(net893),
    .X(net892));
 sky130_fd_sc_hd__clkbuf_4 fanout893 (.A(net894),
    .X(net893));
 sky130_fd_sc_hd__buf_2 fanout894 (.A(net901),
    .X(net894));
 sky130_fd_sc_hd__clkbuf_4 fanout895 (.A(net900),
    .X(net895));
 sky130_fd_sc_hd__clkbuf_2 fanout896 (.A(net900),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_4 fanout897 (.A(net899),
    .X(net897));
 sky130_fd_sc_hd__clkbuf_2 fanout898 (.A(net899),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_4 fanout899 (.A(net900),
    .X(net899));
 sky130_fd_sc_hd__clkbuf_4 fanout900 (.A(net901),
    .X(net900));
 sky130_fd_sc_hd__buf_4 fanout901 (.A(\brancher.imm21_j[1] ),
    .X(net901));
 sky130_fd_sc_hd__buf_4 fanout902 (.A(net903),
    .X(net902));
 sky130_fd_sc_hd__buf_4 fanout903 (.A(net907),
    .X(net903));
 sky130_fd_sc_hd__buf_4 fanout904 (.A(net906),
    .X(net904));
 sky130_fd_sc_hd__buf_4 fanout905 (.A(net906),
    .X(net905));
 sky130_fd_sc_hd__buf_2 fanout906 (.A(net907),
    .X(net906));
 sky130_fd_sc_hd__buf_2 fanout907 (.A(net937),
    .X(net907));
 sky130_fd_sc_hd__buf_4 fanout908 (.A(net910),
    .X(net908));
 sky130_fd_sc_hd__buf_4 fanout909 (.A(net910),
    .X(net909));
 sky130_fd_sc_hd__buf_2 fanout910 (.A(net913),
    .X(net910));
 sky130_fd_sc_hd__buf_4 fanout911 (.A(net913),
    .X(net911));
 sky130_fd_sc_hd__buf_4 fanout912 (.A(net913),
    .X(net912));
 sky130_fd_sc_hd__clkbuf_4 fanout913 (.A(net937),
    .X(net913));
 sky130_fd_sc_hd__buf_4 fanout914 (.A(net915),
    .X(net914));
 sky130_fd_sc_hd__clkbuf_4 fanout915 (.A(net918),
    .X(net915));
 sky130_fd_sc_hd__buf_4 fanout916 (.A(net917),
    .X(net916));
 sky130_fd_sc_hd__buf_4 fanout917 (.A(net918),
    .X(net917));
 sky130_fd_sc_hd__clkbuf_4 fanout918 (.A(net937),
    .X(net918));
 sky130_fd_sc_hd__buf_4 fanout919 (.A(net921),
    .X(net919));
 sky130_fd_sc_hd__buf_4 fanout920 (.A(net921),
    .X(net920));
 sky130_fd_sc_hd__buf_2 fanout921 (.A(net930),
    .X(net921));
 sky130_fd_sc_hd__buf_4 fanout922 (.A(net923),
    .X(net922));
 sky130_fd_sc_hd__buf_4 fanout923 (.A(net930),
    .X(net923));
 sky130_fd_sc_hd__buf_4 fanout924 (.A(net929),
    .X(net924));
 sky130_fd_sc_hd__buf_4 fanout925 (.A(net929),
    .X(net925));
 sky130_fd_sc_hd__buf_4 fanout926 (.A(net928),
    .X(net926));
 sky130_fd_sc_hd__buf_4 fanout927 (.A(net929),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_2 fanout928 (.A(net929),
    .X(net928));
 sky130_fd_sc_hd__clkbuf_4 fanout929 (.A(net930),
    .X(net929));
 sky130_fd_sc_hd__buf_2 fanout930 (.A(net937),
    .X(net930));
 sky130_fd_sc_hd__buf_4 fanout931 (.A(net936),
    .X(net931));
 sky130_fd_sc_hd__clkbuf_2 fanout932 (.A(net936),
    .X(net932));
 sky130_fd_sc_hd__buf_4 fanout933 (.A(net935),
    .X(net933));
 sky130_fd_sc_hd__buf_2 fanout934 (.A(net935),
    .X(net934));
 sky130_fd_sc_hd__buf_4 fanout935 (.A(net936),
    .X(net935));
 sky130_fd_sc_hd__buf_4 fanout936 (.A(net937),
    .X(net936));
 sky130_fd_sc_hd__buf_4 fanout937 (.A(\brancher.imm21_j[11] ),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_8 fanout938 (.A(net939),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_8 fanout939 (.A(\brancher.imm21_j[4] ),
    .X(net939));
 sky130_fd_sc_hd__buf_2 fanout940 (.A(\brancher.imm21_j[4] ),
    .X(net940));
 sky130_fd_sc_hd__buf_4 fanout941 (.A(net942),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_8 fanout942 (.A(\brancher.imm21_j[4] ),
    .X(net942));
 sky130_fd_sc_hd__clkbuf_4 fanout943 (.A(\brancher.funct3[2] ),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_4 fanout944 (.A(\brancher.imm12_i_s[11] ),
    .X(net944));
 sky130_fd_sc_hd__clkbuf_2 fanout945 (.A(\brancher.imm12_i_s[11] ),
    .X(net945));
 sky130_fd_sc_hd__buf_2 fanout946 (.A(net947),
    .X(net946));
 sky130_fd_sc_hd__buf_2 fanout947 (.A(\brancher.imm12_i_s[11] ),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_4 fanout948 (.A(net951),
    .X(net948));
 sky130_fd_sc_hd__buf_2 fanout949 (.A(net950),
    .X(net949));
 sky130_fd_sc_hd__clkbuf_2 fanout950 (.A(net951),
    .X(net950));
 sky130_fd_sc_hd__clkbuf_4 fanout951 (.A(\dec.op_auipc ),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_4 fanout952 (.A(net953),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_4 fanout953 (.A(\brancher.op_jal ),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_4 fanout954 (.A(\brancher.op_jal ),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_2 fanout955 (.A(\brancher.op_jal ),
    .X(net955));
 sky130_fd_sc_hd__buf_4 fanout956 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__buf_4 fanout957 (.A(\brancher.op_jalr ),
    .X(net957));
 sky130_fd_sc_hd__buf_2 fanout958 (.A(net959),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_2 fanout959 (.A(net960),
    .X(net959));
 sky130_fd_sc_hd__buf_2 fanout960 (.A(\brancher.op_jalr ),
    .X(net960));
 sky130_fd_sc_hd__buf_2 fanout961 (.A(\dec.rStall ),
    .X(net961));
 sky130_fd_sc_hd__buf_2 fanout962 (.A(net963),
    .X(net962));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout963 (.A(\dec.rStall ),
    .X(net963));
 sky130_fd_sc_hd__clkbuf_4 fanout964 (.A(\dec.rStall ),
    .X(net964));
 sky130_fd_sc_hd__buf_4 fanout965 (.A(net966),
    .X(net965));
 sky130_fd_sc_hd__buf_2 fanout966 (.A(net967),
    .X(net966));
 sky130_fd_sc_hd__buf_4 fanout967 (.A(\rReg_d2[3] ),
    .X(net967));
 sky130_fd_sc_hd__buf_2 fanout968 (.A(\rReg_d2[2] ),
    .X(net968));
 sky130_fd_sc_hd__buf_2 fanout969 (.A(\rReg_d2[1] ),
    .X(net969));
 sky130_fd_sc_hd__buf_1 fanout970 (.A(\rReg_d2[1] ),
    .X(net970));
 sky130_fd_sc_hd__clkbuf_4 fanout971 (.A(net972),
    .X(net971));
 sky130_fd_sc_hd__buf_4 fanout972 (.A(net983),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_4 fanout973 (.A(net975),
    .X(net973));
 sky130_fd_sc_hd__buf_2 fanout974 (.A(net975),
    .X(net974));
 sky130_fd_sc_hd__buf_2 fanout975 (.A(net983),
    .X(net975));
 sky130_fd_sc_hd__clkbuf_4 fanout976 (.A(net979),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_4 fanout977 (.A(net979),
    .X(net977));
 sky130_fd_sc_hd__clkbuf_2 fanout978 (.A(net979),
    .X(net978));
 sky130_fd_sc_hd__clkbuf_2 fanout979 (.A(net983),
    .X(net979));
 sky130_fd_sc_hd__clkbuf_4 fanout980 (.A(net981),
    .X(net980));
 sky130_fd_sc_hd__clkbuf_4 fanout981 (.A(net982),
    .X(net981));
 sky130_fd_sc_hd__clkbuf_4 fanout982 (.A(net983),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_4 fanout983 (.A(rOp_memLd2),
    .X(net983));
 sky130_fd_sc_hd__clkbuf_4 fanout984 (.A(net985),
    .X(net984));
 sky130_fd_sc_hd__buf_4 fanout985 (.A(net987),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_4 fanout986 (.A(net987),
    .X(net986));
 sky130_fd_sc_hd__buf_4 fanout987 (.A(\brancher.imm21_j[18] ),
    .X(net987));
 sky130_fd_sc_hd__buf_4 fanout988 (.A(net991),
    .X(net988));
 sky130_fd_sc_hd__buf_4 fanout989 (.A(net991),
    .X(net989));
 sky130_fd_sc_hd__buf_4 fanout990 (.A(net991),
    .X(net990));
 sky130_fd_sc_hd__buf_4 fanout991 (.A(\brancher.imm21_j[18] ),
    .X(net991));
 sky130_fd_sc_hd__buf_4 fanout992 (.A(net993),
    .X(net992));
 sky130_fd_sc_hd__buf_4 fanout993 (.A(net994),
    .X(net993));
 sky130_fd_sc_hd__clkbuf_8 fanout994 (.A(\brancher.imm21_j[17] ),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_8 fanout995 (.A(net997),
    .X(net995));
 sky130_fd_sc_hd__buf_2 fanout996 (.A(net997),
    .X(net996));
 sky130_fd_sc_hd__buf_4 fanout997 (.A(\brancher.imm21_j[17] ),
    .X(net997));
 sky130_fd_sc_hd__clkbuf_4 fanout998 (.A(net1002),
    .X(net998));
 sky130_fd_sc_hd__clkbuf_4 fanout999 (.A(net1002),
    .X(net999));
 sky130_fd_sc_hd__clkbuf_4 fanout1000 (.A(net1002),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_4 fanout1001 (.A(net1002),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_4 fanout1002 (.A(net1013),
    .X(net1002));
 sky130_fd_sc_hd__clkbuf_4 fanout1003 (.A(net1005),
    .X(net1003));
 sky130_fd_sc_hd__clkbuf_4 fanout1004 (.A(net1005),
    .X(net1004));
 sky130_fd_sc_hd__clkbuf_2 fanout1005 (.A(net1008),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_4 fanout1006 (.A(net1008),
    .X(net1006));
 sky130_fd_sc_hd__clkbuf_4 fanout1007 (.A(net1008),
    .X(net1007));
 sky130_fd_sc_hd__buf_2 fanout1008 (.A(net1013),
    .X(net1008));
 sky130_fd_sc_hd__clkbuf_4 fanout1009 (.A(net1010),
    .X(net1009));
 sky130_fd_sc_hd__clkbuf_4 fanout1010 (.A(net1013),
    .X(net1010));
 sky130_fd_sc_hd__clkbuf_4 fanout1011 (.A(net1012),
    .X(net1011));
 sky130_fd_sc_hd__clkbuf_4 fanout1012 (.A(net1013),
    .X(net1012));
 sky130_fd_sc_hd__buf_2 fanout1013 (.A(\brancher.imm21_j[16] ),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_4 fanout1014 (.A(net1016),
    .X(net1014));
 sky130_fd_sc_hd__clkbuf_4 fanout1015 (.A(net1016),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_2 fanout1016 (.A(net1031),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_4 fanout1017 (.A(net1018),
    .X(net1017));
 sky130_fd_sc_hd__clkbuf_4 fanout1018 (.A(net1031),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_4 fanout1019 (.A(net1024),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_4 fanout1020 (.A(net1024),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_4 fanout1021 (.A(net1023),
    .X(net1021));
 sky130_fd_sc_hd__clkbuf_4 fanout1022 (.A(net1024),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_2 fanout1023 (.A(net1024),
    .X(net1023));
 sky130_fd_sc_hd__clkbuf_4 fanout1024 (.A(net1031),
    .X(net1024));
 sky130_fd_sc_hd__clkbuf_4 fanout1025 (.A(net1030),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_2 fanout1026 (.A(net1030),
    .X(net1026));
 sky130_fd_sc_hd__clkbuf_4 fanout1027 (.A(net1029),
    .X(net1027));
 sky130_fd_sc_hd__clkbuf_2 fanout1028 (.A(net1029),
    .X(net1028));
 sky130_fd_sc_hd__clkbuf_4 fanout1029 (.A(net1030),
    .X(net1029));
 sky130_fd_sc_hd__buf_4 fanout1030 (.A(net1031),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_4 fanout1031 (.A(\brancher.imm21_j[16] ),
    .X(net1031));
 sky130_fd_sc_hd__buf_4 fanout1032 (.A(net1036),
    .X(net1032));
 sky130_fd_sc_hd__buf_4 fanout1033 (.A(net1036),
    .X(net1033));
 sky130_fd_sc_hd__buf_4 fanout1034 (.A(net1036),
    .X(net1034));
 sky130_fd_sc_hd__buf_4 fanout1035 (.A(net1036),
    .X(net1035));
 sky130_fd_sc_hd__buf_4 fanout1036 (.A(net1047),
    .X(net1036));
 sky130_fd_sc_hd__buf_4 fanout1037 (.A(net1039),
    .X(net1037));
 sky130_fd_sc_hd__buf_4 fanout1038 (.A(net1039),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_2 fanout1039 (.A(net1042),
    .X(net1039));
 sky130_fd_sc_hd__buf_4 fanout1040 (.A(net1042),
    .X(net1040));
 sky130_fd_sc_hd__buf_4 fanout1041 (.A(net1042),
    .X(net1041));
 sky130_fd_sc_hd__buf_2 fanout1042 (.A(net1047),
    .X(net1042));
 sky130_fd_sc_hd__buf_4 fanout1043 (.A(net1044),
    .X(net1043));
 sky130_fd_sc_hd__clkbuf_4 fanout1044 (.A(net1047),
    .X(net1044));
 sky130_fd_sc_hd__buf_4 fanout1045 (.A(net1046),
    .X(net1045));
 sky130_fd_sc_hd__buf_4 fanout1046 (.A(net1047),
    .X(net1046));
 sky130_fd_sc_hd__clkbuf_4 fanout1047 (.A(\brancher.imm21_j[15] ),
    .X(net1047));
 sky130_fd_sc_hd__buf_4 fanout1048 (.A(net1050),
    .X(net1048));
 sky130_fd_sc_hd__buf_4 fanout1049 (.A(net1050),
    .X(net1049));
 sky130_fd_sc_hd__buf_2 fanout1050 (.A(net1065),
    .X(net1050));
 sky130_fd_sc_hd__buf_4 fanout1051 (.A(net1052),
    .X(net1051));
 sky130_fd_sc_hd__buf_4 fanout1052 (.A(net1065),
    .X(net1052));
 sky130_fd_sc_hd__buf_4 fanout1053 (.A(net1058),
    .X(net1053));
 sky130_fd_sc_hd__buf_4 fanout1054 (.A(net1058),
    .X(net1054));
 sky130_fd_sc_hd__buf_4 fanout1055 (.A(net1057),
    .X(net1055));
 sky130_fd_sc_hd__buf_4 fanout1056 (.A(net1058),
    .X(net1056));
 sky130_fd_sc_hd__clkbuf_2 fanout1057 (.A(net1058),
    .X(net1057));
 sky130_fd_sc_hd__clkbuf_4 fanout1058 (.A(net1065),
    .X(net1058));
 sky130_fd_sc_hd__buf_4 fanout1059 (.A(net1064),
    .X(net1059));
 sky130_fd_sc_hd__buf_2 fanout1060 (.A(net1064),
    .X(net1060));
 sky130_fd_sc_hd__buf_4 fanout1061 (.A(net1063),
    .X(net1061));
 sky130_fd_sc_hd__buf_2 fanout1062 (.A(net1063),
    .X(net1062));
 sky130_fd_sc_hd__buf_4 fanout1063 (.A(net1064),
    .X(net1063));
 sky130_fd_sc_hd__buf_4 fanout1064 (.A(net1065),
    .X(net1064));
 sky130_fd_sc_hd__clkbuf_4 fanout1065 (.A(\brancher.imm21_j[15] ),
    .X(net1065));
 sky130_fd_sc_hd__clkbuf_8 fanout1066 (.A(net1067),
    .X(net1066));
 sky130_fd_sc_hd__clkbuf_8 fanout1067 (.A(net1070),
    .X(net1067));
 sky130_fd_sc_hd__buf_4 fanout1068 (.A(net1069),
    .X(net1068));
 sky130_fd_sc_hd__buf_4 fanout1069 (.A(net1070),
    .X(net1069));
 sky130_fd_sc_hd__buf_4 fanout1070 (.A(\brancher.imm21_j[19] ),
    .X(net1070));
 sky130_fd_sc_hd__clkbuf_2 fanout1071 (.A(net1072),
    .X(net1071));
 sky130_fd_sc_hd__clkbuf_2 fanout1072 (.A(net1073),
    .X(net1072));
 sky130_fd_sc_hd__buf_2 fanout1073 (.A(net1093),
    .X(net1073));
 sky130_fd_sc_hd__clkbuf_2 fanout1074 (.A(net1080),
    .X(net1074));
 sky130_fd_sc_hd__clkbuf_2 fanout1075 (.A(net1080),
    .X(net1075));
 sky130_fd_sc_hd__buf_1 fanout1076 (.A(net1080),
    .X(net1076));
 sky130_fd_sc_hd__clkbuf_2 fanout1077 (.A(net1079),
    .X(net1077));
 sky130_fd_sc_hd__clkbuf_2 fanout1078 (.A(net1079),
    .X(net1078));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1079 (.A(net1080),
    .X(net1079));
 sky130_fd_sc_hd__clkbuf_2 fanout1080 (.A(net1093),
    .X(net1080));
 sky130_fd_sc_hd__clkbuf_2 fanout1081 (.A(net1083),
    .X(net1081));
 sky130_fd_sc_hd__clkbuf_2 fanout1082 (.A(net1083),
    .X(net1082));
 sky130_fd_sc_hd__clkbuf_2 fanout1083 (.A(net1093),
    .X(net1083));
 sky130_fd_sc_hd__clkbuf_2 fanout1084 (.A(net1086),
    .X(net1084));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1085 (.A(net1086),
    .X(net1085));
 sky130_fd_sc_hd__clkbuf_2 fanout1086 (.A(net1093),
    .X(net1086));
 sky130_fd_sc_hd__clkbuf_2 fanout1087 (.A(net1092),
    .X(net1087));
 sky130_fd_sc_hd__clkbuf_2 fanout1088 (.A(net1092),
    .X(net1088));
 sky130_fd_sc_hd__clkbuf_2 fanout1089 (.A(net1091),
    .X(net1089));
 sky130_fd_sc_hd__clkbuf_2 fanout1090 (.A(net1091),
    .X(net1090));
 sky130_fd_sc_hd__clkbuf_2 fanout1091 (.A(net1092),
    .X(net1091));
 sky130_fd_sc_hd__clkbuf_2 fanout1092 (.A(net1093),
    .X(net1092));
 sky130_fd_sc_hd__buf_2 fanout1093 (.A(net1138),
    .X(net1093));
 sky130_fd_sc_hd__clkbuf_2 fanout1094 (.A(net1096),
    .X(net1094));
 sky130_fd_sc_hd__clkbuf_2 fanout1095 (.A(net1096),
    .X(net1095));
 sky130_fd_sc_hd__clkbuf_2 fanout1096 (.A(net1105),
    .X(net1096));
 sky130_fd_sc_hd__clkbuf_2 fanout1097 (.A(net1098),
    .X(net1097));
 sky130_fd_sc_hd__clkbuf_2 fanout1098 (.A(net1105),
    .X(net1098));
 sky130_fd_sc_hd__clkbuf_2 fanout1099 (.A(net1100),
    .X(net1099));
 sky130_fd_sc_hd__clkbuf_2 fanout1100 (.A(net1105),
    .X(net1100));
 sky130_fd_sc_hd__buf_1 fanout1101 (.A(net1105),
    .X(net1101));
 sky130_fd_sc_hd__clkbuf_2 fanout1102 (.A(net1104),
    .X(net1102));
 sky130_fd_sc_hd__clkbuf_2 fanout1103 (.A(net1104),
    .X(net1103));
 sky130_fd_sc_hd__clkbuf_2 fanout1104 (.A(net1105),
    .X(net1104));
 sky130_fd_sc_hd__buf_2 fanout1105 (.A(net1138),
    .X(net1105));
 sky130_fd_sc_hd__clkbuf_2 fanout1106 (.A(net1112),
    .X(net1106));
 sky130_fd_sc_hd__buf_1 fanout1107 (.A(net1112),
    .X(net1107));
 sky130_fd_sc_hd__clkbuf_2 fanout1108 (.A(net1112),
    .X(net1108));
 sky130_fd_sc_hd__buf_1 fanout1109 (.A(net1112),
    .X(net1109));
 sky130_fd_sc_hd__clkbuf_2 fanout1110 (.A(net1111),
    .X(net1110));
 sky130_fd_sc_hd__clkbuf_2 fanout1111 (.A(net1112),
    .X(net1111));
 sky130_fd_sc_hd__clkbuf_2 fanout1112 (.A(net1138),
    .X(net1112));
 sky130_fd_sc_hd__clkbuf_2 fanout1113 (.A(net1117),
    .X(net1113));
 sky130_fd_sc_hd__clkbuf_2 fanout1114 (.A(net1117),
    .X(net1114));
 sky130_fd_sc_hd__clkbuf_2 fanout1115 (.A(net1116),
    .X(net1115));
 sky130_fd_sc_hd__clkbuf_2 fanout1116 (.A(net1117),
    .X(net1116));
 sky130_fd_sc_hd__clkbuf_2 fanout1117 (.A(net1138),
    .X(net1117));
 sky130_fd_sc_hd__clkbuf_2 fanout1118 (.A(net1123),
    .X(net1118));
 sky130_fd_sc_hd__buf_1 fanout1119 (.A(net1123),
    .X(net1119));
 sky130_fd_sc_hd__clkbuf_2 fanout1120 (.A(net1123),
    .X(net1120));
 sky130_fd_sc_hd__clkbuf_2 fanout1121 (.A(net1122),
    .X(net1121));
 sky130_fd_sc_hd__clkbuf_2 fanout1122 (.A(net1123),
    .X(net1122));
 sky130_fd_sc_hd__buf_2 fanout1123 (.A(net1134),
    .X(net1123));
 sky130_fd_sc_hd__clkbuf_2 fanout1124 (.A(net1125),
    .X(net1124));
 sky130_fd_sc_hd__buf_2 fanout1125 (.A(net1134),
    .X(net1125));
 sky130_fd_sc_hd__clkbuf_2 fanout1126 (.A(net1128),
    .X(net1126));
 sky130_fd_sc_hd__buf_1 fanout1127 (.A(net1128),
    .X(net1127));
 sky130_fd_sc_hd__clkbuf_2 fanout1128 (.A(net1131),
    .X(net1128));
 sky130_fd_sc_hd__clkbuf_2 fanout1129 (.A(net1131),
    .X(net1129));
 sky130_fd_sc_hd__clkbuf_2 fanout1130 (.A(net1131),
    .X(net1130));
 sky130_fd_sc_hd__clkbuf_2 fanout1131 (.A(net1134),
    .X(net1131));
 sky130_fd_sc_hd__clkbuf_2 fanout1132 (.A(net1133),
    .X(net1132));
 sky130_fd_sc_hd__clkbuf_2 fanout1133 (.A(net1134),
    .X(net1133));
 sky130_fd_sc_hd__clkbuf_2 fanout1134 (.A(net1138),
    .X(net1134));
 sky130_fd_sc_hd__clkbuf_4 fanout1135 (.A(net1137),
    .X(net1135));
 sky130_fd_sc_hd__clkbuf_2 fanout1136 (.A(net1137),
    .X(net1136));
 sky130_fd_sc_hd__buf_2 fanout1137 (.A(net1138),
    .X(net1137));
 sky130_fd_sc_hd__buf_4 fanout1138 (.A(net1210),
    .X(net1138));
 sky130_fd_sc_hd__clkbuf_2 fanout1139 (.A(net1141),
    .X(net1139));
 sky130_fd_sc_hd__clkbuf_2 fanout1140 (.A(net1141),
    .X(net1140));
 sky130_fd_sc_hd__clkbuf_2 fanout1141 (.A(net1151),
    .X(net1141));
 sky130_fd_sc_hd__clkbuf_2 fanout1142 (.A(net1144),
    .X(net1142));
 sky130_fd_sc_hd__clkbuf_2 fanout1143 (.A(net1151),
    .X(net1143));
 sky130_fd_sc_hd__buf_1 fanout1144 (.A(net1151),
    .X(net1144));
 sky130_fd_sc_hd__clkbuf_2 fanout1145 (.A(net1147),
    .X(net1145));
 sky130_fd_sc_hd__clkbuf_2 fanout1146 (.A(net1147),
    .X(net1146));
 sky130_fd_sc_hd__clkbuf_2 fanout1147 (.A(net1151),
    .X(net1147));
 sky130_fd_sc_hd__clkbuf_2 fanout1148 (.A(net1150),
    .X(net1148));
 sky130_fd_sc_hd__clkbuf_2 fanout1149 (.A(net1150),
    .X(net1149));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1150 (.A(net1151),
    .X(net1150));
 sky130_fd_sc_hd__clkbuf_2 fanout1151 (.A(net1187),
    .X(net1151));
 sky130_fd_sc_hd__clkbuf_2 fanout1152 (.A(net1154),
    .X(net1152));
 sky130_fd_sc_hd__clkbuf_2 fanout1153 (.A(net1154),
    .X(net1153));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1154 (.A(net1187),
    .X(net1154));
 sky130_fd_sc_hd__clkbuf_2 fanout1155 (.A(net1157),
    .X(net1155));
 sky130_fd_sc_hd__clkbuf_2 fanout1156 (.A(net1157),
    .X(net1156));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1157 (.A(net1187),
    .X(net1157));
 sky130_fd_sc_hd__clkbuf_2 fanout1158 (.A(net1160),
    .X(net1158));
 sky130_fd_sc_hd__clkbuf_2 fanout1159 (.A(net1160),
    .X(net1159));
 sky130_fd_sc_hd__clkbuf_2 fanout1160 (.A(net1163),
    .X(net1160));
 sky130_fd_sc_hd__clkbuf_2 fanout1161 (.A(net1162),
    .X(net1161));
 sky130_fd_sc_hd__buf_2 fanout1162 (.A(net1163),
    .X(net1162));
 sky130_fd_sc_hd__clkbuf_2 fanout1163 (.A(net1187),
    .X(net1163));
 sky130_fd_sc_hd__clkbuf_2 fanout1164 (.A(net1166),
    .X(net1164));
 sky130_fd_sc_hd__clkbuf_2 fanout1165 (.A(net1166),
    .X(net1165));
 sky130_fd_sc_hd__clkbuf_2 fanout1166 (.A(net1186),
    .X(net1166));
 sky130_fd_sc_hd__clkbuf_2 fanout1167 (.A(net1169),
    .X(net1167));
 sky130_fd_sc_hd__clkbuf_2 fanout1168 (.A(net1169),
    .X(net1168));
 sky130_fd_sc_hd__clkbuf_2 fanout1169 (.A(net1186),
    .X(net1169));
 sky130_fd_sc_hd__clkbuf_2 fanout1170 (.A(net1174),
    .X(net1170));
 sky130_fd_sc_hd__clkbuf_2 fanout1171 (.A(net1173),
    .X(net1171));
 sky130_fd_sc_hd__clkbuf_2 fanout1172 (.A(net1173),
    .X(net1172));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1173 (.A(net1174),
    .X(net1173));
 sky130_fd_sc_hd__clkbuf_2 fanout1174 (.A(net1186),
    .X(net1174));
 sky130_fd_sc_hd__clkbuf_2 fanout1175 (.A(net1177),
    .X(net1175));
 sky130_fd_sc_hd__clkbuf_2 fanout1176 (.A(net1177),
    .X(net1176));
 sky130_fd_sc_hd__clkbuf_2 fanout1177 (.A(net1186),
    .X(net1177));
 sky130_fd_sc_hd__clkbuf_2 fanout1178 (.A(net1186),
    .X(net1178));
 sky130_fd_sc_hd__buf_1 fanout1179 (.A(net1186),
    .X(net1179));
 sky130_fd_sc_hd__clkbuf_2 fanout1180 (.A(net1181),
    .X(net1180));
 sky130_fd_sc_hd__clkbuf_2 fanout1181 (.A(net1185),
    .X(net1181));
 sky130_fd_sc_hd__clkbuf_2 fanout1182 (.A(net1184),
    .X(net1182));
 sky130_fd_sc_hd__clkbuf_2 fanout1183 (.A(net1184),
    .X(net1183));
 sky130_fd_sc_hd__buf_1 fanout1184 (.A(net1185),
    .X(net1184));
 sky130_fd_sc_hd__clkbuf_2 fanout1185 (.A(net1186),
    .X(net1185));
 sky130_fd_sc_hd__buf_2 fanout1186 (.A(net1187),
    .X(net1186));
 sky130_fd_sc_hd__clkbuf_2 fanout1187 (.A(net1210),
    .X(net1187));
 sky130_fd_sc_hd__buf_2 fanout1188 (.A(net1210),
    .X(net1188));
 sky130_fd_sc_hd__clkbuf_2 fanout1189 (.A(net1210),
    .X(net1189));
 sky130_fd_sc_hd__buf_2 fanout1190 (.A(net1191),
    .X(net1190));
 sky130_fd_sc_hd__buf_2 fanout1191 (.A(net1209),
    .X(net1191));
 sky130_fd_sc_hd__clkbuf_2 fanout1192 (.A(net1194),
    .X(net1192));
 sky130_fd_sc_hd__clkbuf_2 fanout1193 (.A(net1194),
    .X(net1193));
 sky130_fd_sc_hd__clkbuf_2 fanout1194 (.A(net1198),
    .X(net1194));
 sky130_fd_sc_hd__clkbuf_2 fanout1195 (.A(net1198),
    .X(net1195));
 sky130_fd_sc_hd__clkbuf_2 fanout1196 (.A(net1198),
    .X(net1196));
 sky130_fd_sc_hd__buf_1 fanout1197 (.A(net1198),
    .X(net1197));
 sky130_fd_sc_hd__clkbuf_2 fanout1198 (.A(net1209),
    .X(net1198));
 sky130_fd_sc_hd__clkbuf_2 fanout1199 (.A(net1200),
    .X(net1199));
 sky130_fd_sc_hd__clkbuf_2 fanout1200 (.A(net1203),
    .X(net1200));
 sky130_fd_sc_hd__clkbuf_2 fanout1201 (.A(net1203),
    .X(net1201));
 sky130_fd_sc_hd__clkbuf_2 fanout1202 (.A(net1203),
    .X(net1202));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1203 (.A(net1209),
    .X(net1203));
 sky130_fd_sc_hd__clkbuf_2 fanout1204 (.A(net1206),
    .X(net1204));
 sky130_fd_sc_hd__clkbuf_2 fanout1205 (.A(net1206),
    .X(net1205));
 sky130_fd_sc_hd__buf_1 fanout1206 (.A(net1208),
    .X(net1206));
 sky130_fd_sc_hd__clkbuf_2 fanout1207 (.A(net1208),
    .X(net1207));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1208 (.A(net1209),
    .X(net1208));
 sky130_fd_sc_hd__buf_2 fanout1209 (.A(net1210),
    .X(net1209));
 sky130_fd_sc_hd__buf_4 fanout1210 (.A(net66),
    .X(net1210));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_4_1_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_4_4_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_4_5_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_44_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_45_clk (.A(clknet_4_7_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_46_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_47_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_48_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_49_clk (.A(clknet_4_6_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_50_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_51_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_52_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_53_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_54_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_55_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_56_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_57_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_58_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_59_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_60_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_61_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_62_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_63_clk (.A(clknet_4_15_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_64_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_65_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_66_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_67_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_68_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_69_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_70_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_71_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_72_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_73_clk (.A(clknet_4_13_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_74_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_75_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_76_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_77_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_78_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_79_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_80_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_81_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_82_clk (.A(clknet_4_12_0_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_83_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_84_clk (.A(clknet_4_14_0_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_85_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_86_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_87_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_88_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_89_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_90_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_91_clk (.A(clknet_4_11_0_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_92_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_93_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_94_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_95_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_96_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_97_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_98_clk (.A(clknet_4_10_0_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_99_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_100_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_101_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_102_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_103_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_104_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_105_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_106_clk (.A(clknet_4_8_0_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_107_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_108_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_109_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_110_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_111_clk (.A(clknet_4_9_0_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_112_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_113_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_114_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_115_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_116_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_117_clk (.A(clknet_4_3_0_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_118_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_119_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_120_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_121_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_122_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_123_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_124_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_125_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_126_clk (.A(clknet_4_2_0_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_127_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_128_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_129_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_130_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_131_clk (.A(clknet_4_0_0_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_4_0_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_4_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload2 (.A(clknet_4_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload3 (.A(clknet_4_4_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload4 (.A(clknet_4_5_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload5 (.A(clknet_4_7_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload6 (.A(clknet_4_8_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload7 (.A(clknet_4_9_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload8 (.A(clknet_4_10_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload9 (.A(clknet_4_11_0_clk));
 sky130_fd_sc_hd__inv_8 clkload10 (.A(clknet_4_12_0_clk));
 sky130_fd_sc_hd__inv_8 clkload11 (.A(clknet_4_13_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload12 (.A(clknet_4_14_0_clk));
 sky130_fd_sc_hd__inv_8 clkload13 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload14 (.A(clknet_leaf_1_clk));
 sky130_fd_sc_hd__inv_6 clkload15 (.A(clknet_leaf_127_clk));
 sky130_fd_sc_hd__bufinv_16 clkload16 (.A(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload17 (.A(clknet_leaf_129_clk));
 sky130_fd_sc_hd__inv_8 clkload18 (.A(clknet_leaf_130_clk));
 sky130_fd_sc_hd__inv_8 clkload19 (.A(clknet_leaf_131_clk));
 sky130_fd_sc_hd__bufinv_16 clkload20 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload21 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__bufinv_16 clkload22 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload23 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload24 (.A(clknet_leaf_13_clk));
 sky130_fd_sc_hd__bufinv_16 clkload25 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__inv_8 clkload26 (.A(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload27 (.A(clknet_leaf_120_clk));
 sky130_fd_sc_hd__bufinv_16 clkload28 (.A(clknet_leaf_121_clk));
 sky130_fd_sc_hd__inv_6 clkload29 (.A(clknet_leaf_122_clk));
 sky130_fd_sc_hd__inv_8 clkload30 (.A(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload31 (.A(clknet_leaf_124_clk));
 sky130_fd_sc_hd__inv_8 clkload32 (.A(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload33 (.A(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload34 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload35 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload36 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkinv_2 clkload37 (.A(clknet_leaf_112_clk));
 sky130_fd_sc_hd__bufinv_16 clkload38 (.A(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload39 (.A(clknet_leaf_114_clk));
 sky130_fd_sc_hd__bufinv_16 clkload40 (.A(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload41 (.A(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload42 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkinv_4 clkload43 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkinv_4 clkload44 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkinv_4 clkload45 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkinv_2 clkload46 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__bufinv_16 clkload47 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkinv_2 clkload48 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload49 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkinv_4 clkload50 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__bufinv_16 clkload51 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload52 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkinv_4 clkload53 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkinv_2 clkload54 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__bufinv_16 clkload55 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__inv_6 clkload56 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkinv_4 clkload57 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkinv_2 clkload58 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__inv_8 clkload59 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload60 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__inv_6 clkload61 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__inv_8 clkload62 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload63 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkinv_4 clkload64 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__inv_6 clkload65 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__inv_8 clkload66 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload67 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__inv_6 clkload68 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__inv_8 clkload69 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkinv_4 clkload70 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__inv_8 clkload71 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload72 (.A(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload73 (.A(clknet_leaf_102_clk));
 sky130_fd_sc_hd__bufinv_16 clkload74 (.A(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload75 (.A(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkinv_2 clkload76 (.A(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload77 (.A(clknet_leaf_106_clk));
 sky130_fd_sc_hd__inv_6 clkload78 (.A(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkinv_2 clkload79 (.A(clknet_leaf_78_clk));
 sky130_fd_sc_hd__inv_8 clkload80 (.A(clknet_leaf_79_clk));
 sky130_fd_sc_hd__inv_8 clkload81 (.A(clknet_leaf_107_clk));
 sky130_fd_sc_hd__inv_6 clkload82 (.A(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload83 (.A(clknet_leaf_110_clk));
 sky130_fd_sc_hd__inv_6 clkload84 (.A(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkinv_4 clkload85 (.A(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload86 (.A(clknet_leaf_93_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload87 (.A(clknet_leaf_94_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload88 (.A(clknet_leaf_95_clk));
 sky130_fd_sc_hd__bufinv_16 clkload89 (.A(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload90 (.A(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload91 (.A(clknet_leaf_98_clk));
 sky130_fd_sc_hd__bufinv_16 clkload92 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload93 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__inv_6 clkload94 (.A(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload95 (.A(clknet_leaf_87_clk));
 sky130_fd_sc_hd__inv_6 clkload96 (.A(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkinv_2 clkload97 (.A(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkinv_4 clkload98 (.A(clknet_leaf_91_clk));
 sky130_fd_sc_hd__inv_4 clkload99 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload100 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__inv_6 clkload101 (.A(clknet_leaf_74_clk));
 sky130_fd_sc_hd__inv_6 clkload102 (.A(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload103 (.A(clknet_leaf_82_clk));
 sky130_fd_sc_hd__inv_8 clkload104 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload105 (.A(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkinv_4 clkload106 (.A(clknet_leaf_70_clk));
 sky130_fd_sc_hd__inv_6 clkload107 (.A(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkinv_2 clkload108 (.A(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload109 (.A(clknet_leaf_64_clk));
 sky130_fd_sc_hd__inv_6 clkload110 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload111 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__inv_8 clkload112 (.A(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload113 (.A(clknet_leaf_68_clk));
 sky130_fd_sc_hd__inv_8 clkload114 (.A(clknet_leaf_69_clk));
 sky130_fd_sc_hd__inv_6 clkload115 (.A(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkinv_8 clkload116 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__inv_12 clkload117 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkinv_8 clkload118 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkinv_4 clkload119 (.A(clknet_leaf_58_clk));
 sky130_fd_sc_hd__inv_6 clkload120 (.A(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload121 (.A(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload122 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__inv_6 clkload123 (.A(clknet_leaf_63_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\rWrData[24] ),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\rWrData[28] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(rOp_memLd),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\rWrData[12] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\rWrData[16] ),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\rWrData[1] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\rWrData[25] ),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\rWrData[2] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\rWrData[14] ),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\rWrData[22] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\rWrData[21] ),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\rWrData[13] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\rWrData[9] ),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\rWrData[19] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\rWrData[8] ),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\rWrData[20] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\rWrData[15] ),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(rRegWrEn),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\rWrData[0] ),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\rWrData[29] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\rWrData[31] ),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\brancher.imm13_b[2] ),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\rWrData[26] ),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\rWrData[4] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\rReg_d[0] ),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\rWrData[27] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\rReg_d[4] ),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\rWrData[11] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\rWrData[7] ),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\rWrData[18] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\rWrData[5] ),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\brancher.imm13_b[3] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\rWrData[6] ),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\rReg_d[3] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\rReg_d[1] ),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\rWrData[17] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\rWrData[10] ),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\rWrData[3] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\brancher.imm13_b[1] ),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\brancher.imm13_b[11] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\brancher.pc_return[31] ),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\brancher.imm13_b[4] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\reg_module.gprf[1018] ),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\reg_module.gprf[999] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\brancher.pc_return[30] ),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\rReg_d[2] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\reg_module.gprf[1017] ),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\reg_module.gprf[992] ),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\dec.op_memLd ),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\reg_module.gprf[1015] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\reg_module.gprf[1014] ),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\reg_module.gprf[1001] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\reg_module.gprf[1019] ),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\reg_module.gprf[1022] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\reg_module.gprf[1023] ),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\reg_module.gprf[997] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\reg_module.gprf[1013] ),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\reg_module.gprf[1005] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\reg_module.gprf[995] ),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\reg_module.gprf[1003] ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\reg_module.gprf[1012] ),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\reg_module.gprf[1009] ),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\reg_module.gprf[1010] ),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\reg_module.gprf[1006] ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\reg_module.gprf[1021] ),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\reg_module.gprf[1004] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\brancher.rPc_current_reg2[0] ),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_00070_),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\reg_module.gprf[993] ),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\reg_module.gprf[1002] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\brancher.rPc_current_reg2[7] ),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_00077_),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\reg_module.gprf[994] ),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\brancher.rPc_current_reg2[1] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_00071_),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\reg_module.gprf[1008] ),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\reg_module.gprf[1020] ),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\reg_module.gprf[1011] ),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\reg_module.gprf[998] ),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\reg_module.gprf[1000] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\reg_module.gprf[1007] ),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\reg_module.gprf[996] ),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\brancher.rPc_current_reg2[31] ),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\brancher.pc_return[14] ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\brancher.pc_return[17] ),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\brancher.pc_return[13] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_00083_),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\reg_module.gprf[1016] ),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\brancher.pc_return[15] ),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\brancher.pc_return[16] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\brancher.rPc_current_reg2[11] ),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(_00081_),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\brancher.pc_return[9] ),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_00079_),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\brancher.rPc_current_reg2[30] ),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\brancher.pc_return[19] ),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_01190_),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\brancher.pc_return[23] ),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\brancher.pc_return[6] ),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(_00076_),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\brancher.pc_return[12] ),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_00082_),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\brancher.pc_return[18] ),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\brancher.pc_return[11] ),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\brancher.rPc_current_reg2[25] ),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(_00095_),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\brancher.pc_return[22] ),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(_00092_),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\brancher.pc_return[10] ),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_00080_),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\rWrData[30] ),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\rWrData[23] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\brancher.pc_return[2] ),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\brancher.pc_return[4] ),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_00074_),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\brancher.pc_return[5] ),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_00075_),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\brancher.pc_return[8] ),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(_00078_),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\brancher.pc_return[28] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_00098_),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\brancher.pc_return[29] ),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_00099_),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\brancher.rPc_current_reg2[21] ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_00091_),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\brancher.pc_return[24] ),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_00094_),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\brancher.pc_return[25] ),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\dec.op_lui ),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(net156),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\brancher.pc_return[20] ),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_00090_),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\brancher.pc_return[3] ),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\brancher.pc_return[27] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\brancher.pc_return[21] ),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\reg_module.gprf[258] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\brancher.pc_return[1] ),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\reg_module.gprf[269] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\brancher.pc_return[7] ),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\reg_module.gprf[770] ),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\reg_module.gprf[20] ),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\reg_module.gprf[5] ),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\reg_module.gprf[274] ),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\reg_module.gprf[789] ),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\reg_module.gprf[266] ),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\reg_module.gprf[780] ),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\reg_module.gprf[782] ),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\reg_module.gprf[799] ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\reg_module.gprf[772] ),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\reg_module.gprf[284] ),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\reg_module.gprf[796] ),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\reg_module.gprf[263] ),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\reg_module.gprf[797] ),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\reg_module.gprf[774] ),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\reg_module.gprf[30] ),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\reg_module.gprf[790] ),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\reg_module.gprf[8] ),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\reg_module.gprf[283] ),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\reg_module.gprf[279] ),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\reg_module.gprf[785] ),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\reg_module.gprf[28] ),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\reg_module.gprf[25] ),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\reg_module.gprf[775] ),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\brancher.rPc_current_reg2[3] ),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\reg_module.gprf[278] ),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\reg_module.gprf[27] ),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\reg_module.gprf[788] ),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\reg_module.gprf[14] ),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\reg_module.gprf[270] ),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\reg_module.gprf[268] ),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\reg_module.gprf[7] ),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\reg_module.gprf[3] ),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\reg_module.gprf[277] ),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\reg_module.gprf[264] ),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\reg_module.gprf[261] ),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\reg_module.gprf[260] ),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\reg_module.gprf[257] ),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\reg_module.gprf[4] ),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\reg_module.gprf[794] ),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\reg_module.gprf[781] ),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\reg_module.gprf[771] ),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\reg_module.gprf[259] ),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\reg_module.gprf[2] ),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\reg_module.gprf[11] ),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\reg_module.gprf[792] ),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\reg_module.gprf[275] ),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\reg_module.gprf[784] ),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\reg_module.gprf[285] ),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\reg_module.gprf[286] ),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\reg_module.gprf[793] ),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\reg_module.gprf[1] ),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\reg_module.gprf[24] ),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\reg_module.gprf[281] ),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\reg_module.gprf[262] ),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\reg_module.gprf[23] ),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\reg_module.gprf[267] ),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\reg_module.gprf[10] ),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\reg_module.gprf[280] ),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\reg_module.gprf[273] ),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\reg_module.gprf[791] ),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\reg_module.gprf[12] ),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\reg_module.gprf[17] ),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\reg_module.gprf[26] ),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\reg_module.gprf[31] ),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\reg_module.gprf[16] ),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\reg_module.gprf[787] ),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\reg_module.gprf[272] ),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\dec.op_intRegImm ),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\reg_module.gprf[6] ),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\reg_module.gprf[13] ),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\reg_module.gprf[769] ),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\reg_module.gprf[276] ),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\reg_module.gprf[282] ),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\reg_module.gprf[287] ),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\reg_module.gprf[786] ),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\reg_module.gprf[29] ),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\reg_module.gprf[783] ),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\reg_module.gprf[265] ),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\reg_module.gprf[773] ),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\reg_module.gprf[18] ),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\reg_module.gprf[9] ),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\reg_module.gprf[798] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\brancher.pc_return[26] ),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\reg_module.gprf[21] ),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\reg_module.gprf[271] ),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\reg_module.gprf[777] ),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\reg_module.gprf[795] ),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\reg_module.gprf[776] ),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\brancher.pc_return[0] ),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\reg_module.gprf[15] ),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\reg_module.gprf[19] ),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\reg_module.gprf[22] ),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\reg_module.gprf[779] ),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\reg_module.gprf[778] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\brancher.rPc_current_reg2[26] ),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\reg_module.gprf[0] ),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\alu.op_consShf ),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\brancher.imm13_b[6] ),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\brancher.imm13_b[8] ),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\brancher.imm13_b[9] ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\dec.rInstrustion[14] ),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\brancher.pc_return[27] ),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\brancher.pc_return[26] ),
    .X(net1453));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_01237_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_01237_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_01238_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_01985_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_03184_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_03219_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_03612_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_04177_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_04177_));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(_04245_));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(_04245_));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_04280_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(_04348_));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(_04579_));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(_04580_));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(_04712_));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(_04712_));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(_04843_));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(_05043_));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(_05076_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(_05109_));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(_05142_));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(_05274_));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(_05307_));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(_05307_));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(_05340_));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(_05373_));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(_05406_));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\brancher.imm21_j[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\brancher.imm21_j[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\brancher.imm21_j[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\brancher.op_jalr ));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(net380));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(net382));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(net585));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(net631));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(net820));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(net856));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(net937));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(net1070));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(_02581_));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(_02682_));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(_02854_));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(_04279_));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(_04314_));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(_04382_));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(_04645_));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(_04711_));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(_05274_));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(_05406_));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(_05453_));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(_05453_));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(\rWrDataWB[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(net370));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(net379));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(net383));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(net939));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(net942));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(net987));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(net995));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(net1065));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(_05142_));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(net378));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(net817));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(net835));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_854 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_914 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_16 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_24 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_777 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_915 ();
endmodule
