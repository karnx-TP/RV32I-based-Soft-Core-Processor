module uart_tb ();

localparam CLK_PERIOD = 10;

//Wire
logic			clk;
logic			rstB;
logic			rx;
logic		dataEn;
logic[7:0]	dataOut;

logic		FfRdEn;
logic[7:0]  dataFFOut;
logic       FfEmpty;
logic       FfFull;
logic		tx;

//Module
uart_rx #(
	.BAUD_CYCLE(868), //BAUD_RATE = 115200 for clk=10n
	.LSB_FIRST(1'b1)
) rx_module (
    .clk(clk),
    .rstB(rstB),

    .rx(rx),
    
    .dataEn(dataEn),
    .dataOut(dataOut),
	.FfFull(FfFull)
);

sync_fifo #(
    .WIDTH(8),
    .DEPTH(256)
) ff (
    .clk(clk),
    .rst(rstB),

    .data_in(dataOut),
    .FfWrEn(dataEn),
    .FfRdEn(FfRdEn),

    .data_out(dataFFOut),
    .FfEmpty(FfEmpty),
    .FfFull(FfFull)
);

uart_tx_ff #(
    parameter BAUD_CYCLE = 868, //BAUD_RATE = 115200 for clk=10n
	parameter LSB_FIRST = 1'b1
) tx_module (
    .clk(clk),
    .rstB(rstB),

    .ffEmpty(FfEmpty),
    .rdEn(FfRdEn),
    .rdData(dataFFOut),
    
    .tx(tx)
);


//Test Signal
int TM = 0;
logic[7:0]	data;
logic[9:0] data_ss;


//Task
    always 
    begin : clock
      #(CLK_PERIOD / 2) 
      clk = 0;
      #(CLK_PERIOD / 2) 
      clk = 1;
    end

    task init;
    begin
        rstB = 0;
		rx = 1;
        #(CLK_PERIOD + 0.5*CLK_PERIOD);
        rstB = 1;
        #(2 * CLK_PERIOD);
    end
    endtask

    initial begin
        init();
        data = 8'h5C;
		data_ss = {1'b1,data,1'b0};
		for(int i=0;i<10;i++)
		begin
			rx = data_ss[i];
			#(868*CLK_PERIOD);
		end

		data = 8'hCC;
		data_ss = {1'b1,data,1'b0};
		for(int i=0;i<10;i++)
		begin
			rx = data_ss[i];
			#(868*CLK_PERIOD);
		end

		data = 8'h00;
		data_ss = {1'b1,data,1'b0};
		for(int i=0;i<10;i++)
		begin
			rx = data_ss[i];
			#(865*CLK_PERIOD);
		end

		data = 8'hFF;
		data_ss = {1'b1,data,1'b0};
		for(int i=0;i<10;i++)
		begin
			rx = data_ss[i];
			#(872*CLK_PERIOD);
		end

		$display("test end");
        $stop;
    end


endmodule
