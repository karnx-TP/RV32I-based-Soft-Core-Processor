module rv32i_core (clk,
    clkEn,
    dataBusInEn,
    rdEn,
    rstB,
    wrEn,
    RamMode,
    addr,
    dataBusIn,
    dataBusOut,
    inst_in,
    pc);
 input clk;
 input clkEn;
 input dataBusInEn;
 output rdEn;
 input rstB;
 output wrEn;
 output [3:0] RamMode;
 output [31:0] addr;
 input [31:0] dataBusIn;
 output [31:0] dataBusOut;
 input [31:0] inst_in;
 output [31:0] pc;

 wire \Op_code[0] ;
 wire \Op_code[1] ;
 wire \Op_code[2] ;
 wire \Op_code[3] ;
 wire \Op_code[4] ;
 wire \Op_code[5] ;
 wire \Op_code[6] ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire b_type;
 wire \funct3[0] ;
 wire \funct3[1] ;
 wire \funct7[0] ;
 wire \funct7[1] ;
 wire \funct7[2] ;
 wire \funct7[3] ;
 wire \funct7[4] ;
 wire \funct7[5] ;
 wire \funct7[6] ;
 wire i_type;
 wire \imm12_i_s[0] ;
 wire \imm12_i_s[10] ;
 wire \imm12_i_s[11] ;
 wire \imm12_i_s[1] ;
 wire \imm12_i_s[2] ;
 wire \imm12_i_s[3] ;
 wire \imm12_i_s[4] ;
 wire \imm12_i_s[5] ;
 wire \imm12_i_s[6] ;
 wire \imm12_i_s[7] ;
 wire \imm12_i_s[8] ;
 wire \imm12_i_s[9] ;
 wire net1075;
 wire \imm13_b[10] ;
 wire \imm13_b[11] ;
 wire \imm13_b[12] ;
 wire \imm13_b[1] ;
 wire \imm13_b[2] ;
 wire \imm13_b[3] ;
 wire \imm13_b[4] ;
 wire \imm13_b[5] ;
 wire \imm13_b[6] ;
 wire \imm13_b[7] ;
 wire \imm13_b[8] ;
 wire \imm13_b[9] ;
 wire net1076;
 wire \imm21_j[10] ;
 wire \imm21_j[11] ;
 wire \imm21_j[12] ;
 wire \imm21_j[13] ;
 wire \imm21_j[14] ;
 wire \imm21_j[15] ;
 wire \imm21_j[16] ;
 wire \imm21_j[17] ;
 wire \imm21_j[18] ;
 wire \imm21_j[19] ;
 wire \imm21_j[1] ;
 wire \imm21_j[20] ;
 wire \imm21_j[2] ;
 wire \imm21_j[3] ;
 wire \imm21_j[4] ;
 wire \imm21_j[5] ;
 wire \imm21_j[6] ;
 wire \imm21_j[7] ;
 wire \imm21_j[8] ;
 wire \imm21_j[9] ;
 wire net1078;
 wire net1098;
 wire clknet_leaf_0_clk;
 wire \imm32_u[12] ;
 wire \imm32_u[13] ;
 wire \imm32_u[14] ;
 wire \imm32_u[15] ;
 wire \imm32_u[16] ;
 wire \imm32_u[17] ;
 wire \imm32_u[18] ;
 wire \imm32_u[19] ;
 wire net1080;
 wire \imm32_u[20] ;
 wire \imm32_u[21] ;
 wire \imm32_u[22] ;
 wire \imm32_u[23] ;
 wire \imm32_u[24] ;
 wire \imm32_u[25] ;
 wire \imm32_u[26] ;
 wire \imm32_u[27] ;
 wire \imm32_u[28] ;
 wire \imm32_u[29] ;
 wire net1082;
 wire \imm32_u[30] ;
 wire \imm32_u[31] ;
 wire net1084;
 wire net1086;
 wire net1088;
 wire net1090;
 wire net1092;
 wire net1094;
 wire net1096;
 wire j_type;
 wire op_auipc;
 wire op_branch;
 wire op_consShf;
 wire op_ecb;
 wire op_efence;
 wire op_intRegImm;
 wire op_intRegReg;
 wire op_jal;
 wire op_jalr;
 wire op_lui;
 wire op_memLd;
 wire op_memSt;
 wire rCond;
 wire rHazardStallRs1;
 wire rHazardStallRs2;
 wire rJumping1;
 wire rJumping2;
 wire rOp_memLd;
 wire rOp_memLd2;
 wire rRegWrEn;
 wire rRegWrEn2;
 wire \rReg_d2[0] ;
 wire \rReg_d2[1] ;
 wire \rReg_d2[2] ;
 wire \rReg_d2[3] ;
 wire \rReg_d2[4] ;
 wire \rReg_d[0] ;
 wire \rReg_d[1] ;
 wire \rReg_d[2] ;
 wire \rReg_d[3] ;
 wire \rReg_d[4] ;
 wire rStall2;
 wire \rWrDataWB[0] ;
 wire \rWrDataWB[10] ;
 wire \rWrDataWB[11] ;
 wire \rWrDataWB[12] ;
 wire \rWrDataWB[13] ;
 wire \rWrDataWB[14] ;
 wire \rWrDataWB[15] ;
 wire \rWrDataWB[16] ;
 wire \rWrDataWB[17] ;
 wire \rWrDataWB[18] ;
 wire \rWrDataWB[19] ;
 wire \rWrDataWB[1] ;
 wire \rWrDataWB[20] ;
 wire \rWrDataWB[21] ;
 wire \rWrDataWB[22] ;
 wire \rWrDataWB[23] ;
 wire \rWrDataWB[24] ;
 wire \rWrDataWB[25] ;
 wire \rWrDataWB[26] ;
 wire \rWrDataWB[27] ;
 wire \rWrDataWB[28] ;
 wire \rWrDataWB[29] ;
 wire \rWrDataWB[2] ;
 wire \rWrDataWB[30] ;
 wire \rWrDataWB[31] ;
 wire \rWrDataWB[3] ;
 wire \rWrDataWB[4] ;
 wire \rWrDataWB[5] ;
 wire \rWrDataWB[6] ;
 wire \rWrDataWB[7] ;
 wire \rWrDataWB[8] ;
 wire \rWrDataWB[9] ;
 wire \rWrData[0] ;
 wire \rWrData[10] ;
 wire \rWrData[11] ;
 wire \rWrData[12] ;
 wire \rWrData[13] ;
 wire \rWrData[14] ;
 wire \rWrData[15] ;
 wire \rWrData[16] ;
 wire \rWrData[17] ;
 wire \rWrData[18] ;
 wire \rWrData[19] ;
 wire \rWrData[1] ;
 wire \rWrData[20] ;
 wire \rWrData[21] ;
 wire \rWrData[22] ;
 wire \rWrData[23] ;
 wire \rWrData[24] ;
 wire \rWrData[25] ;
 wire \rWrData[26] ;
 wire \rWrData[27] ;
 wire \rWrData[28] ;
 wire \rWrData[29] ;
 wire \rWrData[2] ;
 wire \rWrData[30] ;
 wire \rWrData[31] ;
 wire \rWrData[3] ;
 wire \rWrData[4] ;
 wire \rWrData[5] ;
 wire \rWrData[6] ;
 wire \rWrData[7] ;
 wire \rWrData[8] ;
 wire \rWrData[9] ;
 wire r_type;
 wire \reg_d[0] ;
 wire \reg_d[1] ;
 wire \reg_d[2] ;
 wire \reg_d[3] ;
 wire \reg_d[4] ;
 wire \reg_s1[0] ;
 wire \reg_s1[1] ;
 wire \reg_s1[2] ;
 wire \reg_s1[3] ;
 wire \reg_s1[4] ;
 wire \reg_s2[0] ;
 wire \reg_s2[1] ;
 wire \reg_s2[2] ;
 wire \reg_s2[3] ;
 wire \reg_s2[4] ;
 wire s_type;
 wire u_type;
 wire \wAluA[0] ;
 wire \wAluA[10] ;
 wire \wAluA[11] ;
 wire \wAluA[12] ;
 wire \wAluA[13] ;
 wire \wAluA[14] ;
 wire \wAluA[15] ;
 wire \wAluA[16] ;
 wire \wAluA[17] ;
 wire \wAluA[18] ;
 wire \wAluA[19] ;
 wire \wAluA[1] ;
 wire \wAluA[20] ;
 wire \wAluA[21] ;
 wire \wAluA[22] ;
 wire \wAluA[23] ;
 wire \wAluA[24] ;
 wire \wAluA[25] ;
 wire \wAluA[26] ;
 wire \wAluA[27] ;
 wire \wAluA[28] ;
 wire \wAluA[29] ;
 wire \wAluA[2] ;
 wire \wAluA[30] ;
 wire \wAluA[31] ;
 wire \wAluA[3] ;
 wire \wAluA[4] ;
 wire \wAluA[5] ;
 wire \wAluA[6] ;
 wire \wAluA[7] ;
 wire \wAluA[8] ;
 wire \wAluA[9] ;
 wire \wAluB[0] ;
 wire \wAluB[10] ;
 wire \wAluB[11] ;
 wire \wAluB[12] ;
 wire \wAluB[13] ;
 wire \wAluB[14] ;
 wire \wAluB[15] ;
 wire \wAluB[16] ;
 wire \wAluB[17] ;
 wire \wAluB[18] ;
 wire \wAluB[19] ;
 wire \wAluB[1] ;
 wire \wAluB[20] ;
 wire \wAluB[21] ;
 wire \wAluB[22] ;
 wire \wAluB[23] ;
 wire \wAluB[24] ;
 wire \wAluB[25] ;
 wire \wAluB[26] ;
 wire \wAluB[27] ;
 wire \wAluB[28] ;
 wire \wAluB[29] ;
 wire \wAluB[2] ;
 wire \wAluB[30] ;
 wire \wAluB[31] ;
 wire \wAluB[3] ;
 wire \wAluB[4] ;
 wire \wAluB[5] ;
 wire \wAluB[6] ;
 wire \wAluB[7] ;
 wire \wAluB[8] ;
 wire \wAluB[9] ;
 wire wAluFlag;
 wire \wAluOut[0] ;
 wire \wAluOut[10] ;
 wire \wAluOut[11] ;
 wire \wAluOut[12] ;
 wire \wAluOut[13] ;
 wire \wAluOut[14] ;
 wire \wAluOut[15] ;
 wire \wAluOut[16] ;
 wire \wAluOut[17] ;
 wire \wAluOut[18] ;
 wire \wAluOut[19] ;
 wire \wAluOut[1] ;
 wire \wAluOut[20] ;
 wire \wAluOut[21] ;
 wire \wAluOut[22] ;
 wire \wAluOut[23] ;
 wire \wAluOut[24] ;
 wire \wAluOut[25] ;
 wire \wAluOut[26] ;
 wire \wAluOut[27] ;
 wire \wAluOut[28] ;
 wire \wAluOut[29] ;
 wire \wAluOut[2] ;
 wire \wAluOut[30] ;
 wire \wAluOut[31] ;
 wire \wAluOut[3] ;
 wire \wAluOut[4] ;
 wire \wAluOut[5] ;
 wire \wAluOut[6] ;
 wire \wAluOut[7] ;
 wire \wAluOut[8] ;
 wire \wAluOut[9] ;
 wire wAluSextEn;
 wire wCond;
 wire \wFunct3_aluIn[0] ;
 wire \wFunct3_aluIn[1] ;
 wire \wFunct3_aluIn[2] ;
 wire \wFunct7_aluIn[0] ;
 wire \wFunct7_aluIn[1] ;
 wire \wFunct7_aluIn[2] ;
 wire \wFunct7_aluIn[3] ;
 wire \wFunct7_aluIn[4] ;
 wire \wFunct7_aluIn[5] ;
 wire \wFunct7_aluIn[6] ;
 wire wJmp;
 wire wJumping;
 wire \wPcNextCond[0] ;
 wire \wPcNextCond[10] ;
 wire \wPcNextCond[11] ;
 wire \wPcNextCond[12] ;
 wire \wPcNextCond[13] ;
 wire \wPcNextCond[14] ;
 wire \wPcNextCond[15] ;
 wire \wPcNextCond[16] ;
 wire \wPcNextCond[17] ;
 wire \wPcNextCond[18] ;
 wire \wPcNextCond[19] ;
 wire \wPcNextCond[1] ;
 wire \wPcNextCond[20] ;
 wire \wPcNextCond[21] ;
 wire \wPcNextCond[22] ;
 wire \wPcNextCond[23] ;
 wire \wPcNextCond[24] ;
 wire \wPcNextCond[25] ;
 wire \wPcNextCond[26] ;
 wire \wPcNextCond[27] ;
 wire \wPcNextCond[28] ;
 wire \wPcNextCond[29] ;
 wire \wPcNextCond[2] ;
 wire \wPcNextCond[30] ;
 wire \wPcNextCond[31] ;
 wire \wPcNextCond[3] ;
 wire \wPcNextCond[4] ;
 wire \wPcNextCond[5] ;
 wire \wPcNextCond[6] ;
 wire \wPcNextCond[7] ;
 wire \wPcNextCond[8] ;
 wire \wPcNextCond[9] ;
 wire \wPcReturn[0] ;
 wire \wPcReturn[10] ;
 wire \wPcReturn[11] ;
 wire \wPcReturn[12] ;
 wire \wPcReturn[13] ;
 wire \wPcReturn[14] ;
 wire \wPcReturn[15] ;
 wire \wPcReturn[16] ;
 wire \wPcReturn[17] ;
 wire \wPcReturn[18] ;
 wire \wPcReturn[19] ;
 wire \wPcReturn[1] ;
 wire \wPcReturn[20] ;
 wire \wPcReturn[21] ;
 wire \wPcReturn[22] ;
 wire \wPcReturn[23] ;
 wire \wPcReturn[24] ;
 wire \wPcReturn[25] ;
 wire \wPcReturn[26] ;
 wire \wPcReturn[27] ;
 wire \wPcReturn[28] ;
 wire \wPcReturn[29] ;
 wire \wPcReturn[2] ;
 wire \wPcReturn[30] ;
 wire \wPcReturn[31] ;
 wire \wPcReturn[3] ;
 wire \wPcReturn[4] ;
 wire \wPcReturn[5] ;
 wire \wPcReturn[6] ;
 wire \wPcReturn[7] ;
 wire \wPcReturn[8] ;
 wire \wPcReturn[9] ;
 wire wRamByteEn;
 wire wRamHalfEn;
 wire wRamWordEn;
 wire \wRegWrData[0] ;
 wire \wRegWrData[10] ;
 wire \wRegWrData[11] ;
 wire \wRegWrData[12] ;
 wire \wRegWrData[13] ;
 wire \wRegWrData[14] ;
 wire \wRegWrData[15] ;
 wire \wRegWrData[16] ;
 wire \wRegWrData[17] ;
 wire \wRegWrData[18] ;
 wire \wRegWrData[19] ;
 wire \wRegWrData[1] ;
 wire \wRegWrData[20] ;
 wire \wRegWrData[21] ;
 wire \wRegWrData[22] ;
 wire \wRegWrData[23] ;
 wire \wRegWrData[24] ;
 wire \wRegWrData[25] ;
 wire \wRegWrData[26] ;
 wire \wRegWrData[27] ;
 wire \wRegWrData[28] ;
 wire \wRegWrData[29] ;
 wire \wRegWrData[2] ;
 wire \wRegWrData[30] ;
 wire \wRegWrData[31] ;
 wire \wRegWrData[3] ;
 wire \wRegWrData[4] ;
 wire \wRegWrData[5] ;
 wire \wRegWrData[6] ;
 wire \wRegWrData[7] ;
 wire \wRegWrData[8] ;
 wire \wRegWrData[9] ;
 wire \wReg_s1_out[0] ;
 wire \wReg_s1_out[1] ;
 wire \wReg_s1_out[2] ;
 wire \wReg_s1_out[3] ;
 wire \wReg_s1_out[4] ;
 wire \wReg_s2_out[0] ;
 wire \wReg_s2_out[1] ;
 wire \wReg_s2_out[2] ;
 wire \wReg_s2_out[3] ;
 wire \wReg_s2_out[4] ;
 wire \wRs1Data[0] ;
 wire \wRs1Data[10] ;
 wire \wRs1Data[11] ;
 wire \wRs1Data[12] ;
 wire \wRs1Data[13] ;
 wire \wRs1Data[14] ;
 wire \wRs1Data[15] ;
 wire \wRs1Data[16] ;
 wire \wRs1Data[17] ;
 wire \wRs1Data[18] ;
 wire \wRs1Data[19] ;
 wire \wRs1Data[1] ;
 wire \wRs1Data[20] ;
 wire \wRs1Data[21] ;
 wire \wRs1Data[22] ;
 wire \wRs1Data[23] ;
 wire \wRs1Data[24] ;
 wire \wRs1Data[25] ;
 wire \wRs1Data[26] ;
 wire \wRs1Data[27] ;
 wire \wRs1Data[28] ;
 wire \wRs1Data[29] ;
 wire \wRs1Data[2] ;
 wire \wRs1Data[30] ;
 wire \wRs1Data[31] ;
 wire \wRs1Data[3] ;
 wire \wRs1Data[4] ;
 wire \wRs1Data[5] ;
 wire \wRs1Data[6] ;
 wire \wRs1Data[7] ;
 wire \wRs1Data[8] ;
 wire \wRs1Data[9] ;
 wire \wRs2Data[0] ;
 wire \wRs2Data[10] ;
 wire \wRs2Data[11] ;
 wire \wRs2Data[12] ;
 wire \wRs2Data[13] ;
 wire \wRs2Data[14] ;
 wire \wRs2Data[15] ;
 wire \wRs2Data[16] ;
 wire \wRs2Data[17] ;
 wire \wRs2Data[18] ;
 wire \wRs2Data[19] ;
 wire \wRs2Data[1] ;
 wire \wRs2Data[20] ;
 wire \wRs2Data[21] ;
 wire \wRs2Data[22] ;
 wire \wRs2Data[23] ;
 wire \wRs2Data[24] ;
 wire \wRs2Data[25] ;
 wire \wRs2Data[26] ;
 wire \wRs2Data[27] ;
 wire \wRs2Data[28] ;
 wire \wRs2Data[29] ;
 wire \wRs2Data[2] ;
 wire \wRs2Data[30] ;
 wire \wRs2Data[31] ;
 wire \wRs2Data[3] ;
 wire \wRs2Data[4] ;
 wire \wRs2Data[5] ;
 wire \wRs2Data[6] ;
 wire \wRs2Data[7] ;
 wire \wRs2Data[8] ;
 wire \wRs2Data[9] ;
 wire wStall;
 wire wStall1;
 wire \alu/_0000_ ;
 wire \alu/_0001_ ;
 wire \alu/_0002_ ;
 wire \alu/_0003_ ;
 wire \alu/_0004_ ;
 wire \alu/_0005_ ;
 wire \alu/_0006_ ;
 wire \alu/_0007_ ;
 wire \alu/_0008_ ;
 wire \alu/_0009_ ;
 wire \alu/_0010_ ;
 wire \alu/_0011_ ;
 wire \alu/_0012_ ;
 wire \alu/_0013_ ;
 wire \alu/_0014_ ;
 wire \alu/_0015_ ;
 wire \alu/_0016_ ;
 wire \alu/_0017_ ;
 wire \alu/_0018_ ;
 wire \alu/_0019_ ;
 wire \alu/_0020_ ;
 wire \alu/_0021_ ;
 wire \alu/_0022_ ;
 wire \alu/_0023_ ;
 wire \alu/_0024_ ;
 wire \alu/_0025_ ;
 wire \alu/_0026_ ;
 wire \alu/_0027_ ;
 wire \alu/_0028_ ;
 wire \alu/_0029_ ;
 wire \alu/_0030_ ;
 wire \alu/_0031_ ;
 wire \alu/_0032_ ;
 wire \alu/_0033_ ;
 wire \alu/_0034_ ;
 wire \alu/_0035_ ;
 wire \alu/_0036_ ;
 wire \alu/_0037_ ;
 wire \alu/_0038_ ;
 wire \alu/_0039_ ;
 wire \alu/_0040_ ;
 wire \alu/_0041_ ;
 wire \alu/_0042_ ;
 wire \alu/_0043_ ;
 wire \alu/_0044_ ;
 wire \alu/_0045_ ;
 wire \alu/_0046_ ;
 wire \alu/_0047_ ;
 wire \alu/_0048_ ;
 wire \alu/_0049_ ;
 wire \alu/_0050_ ;
 wire \alu/_0051_ ;
 wire \alu/_0052_ ;
 wire \alu/_0053_ ;
 wire \alu/_0054_ ;
 wire \alu/_0055_ ;
 wire \alu/_0056_ ;
 wire \alu/_0057_ ;
 wire \alu/_0058_ ;
 wire \alu/_0059_ ;
 wire \alu/_0060_ ;
 wire \alu/_0061_ ;
 wire \alu/_0062_ ;
 wire \alu/_0063_ ;
 wire \alu/_0064_ ;
 wire \alu/_0065_ ;
 wire \alu/_0066_ ;
 wire \alu/_0067_ ;
 wire \alu/_0068_ ;
 wire \alu/_0069_ ;
 wire \alu/_0070_ ;
 wire \alu/_0071_ ;
 wire \alu/_0072_ ;
 wire \alu/_0073_ ;
 wire \alu/_0074_ ;
 wire \alu/_0075_ ;
 wire \alu/_0076_ ;
 wire \alu/_0077_ ;
 wire \alu/_0078_ ;
 wire \alu/_0079_ ;
 wire \alu/_0080_ ;
 wire \alu/_0081_ ;
 wire \alu/_0082_ ;
 wire \alu/_0083_ ;
 wire \alu/_0084_ ;
 wire \alu/_0085_ ;
 wire \alu/_0086_ ;
 wire \alu/_0087_ ;
 wire \alu/_0088_ ;
 wire \alu/_0089_ ;
 wire \alu/_0090_ ;
 wire \alu/_0091_ ;
 wire \alu/_0092_ ;
 wire \alu/_0093_ ;
 wire \alu/_0094_ ;
 wire \alu/_0095_ ;
 wire \alu/_0096_ ;
 wire \alu/_0097_ ;
 wire \alu/_0098_ ;
 wire \alu/_0099_ ;
 wire \alu/_0100_ ;
 wire \alu/_0101_ ;
 wire \alu/_0102_ ;
 wire \alu/_0103_ ;
 wire \alu/_0104_ ;
 wire \alu/_0105_ ;
 wire \alu/_0106_ ;
 wire \alu/_0107_ ;
 wire \alu/_0108_ ;
 wire \alu/_0109_ ;
 wire \alu/_0110_ ;
 wire \alu/_0111_ ;
 wire \alu/_0112_ ;
 wire \alu/_0113_ ;
 wire \alu/_0114_ ;
 wire \alu/_0115_ ;
 wire \alu/_0116_ ;
 wire \alu/_0117_ ;
 wire \alu/_0118_ ;
 wire \alu/_0119_ ;
 wire \alu/_0120_ ;
 wire \alu/_0121_ ;
 wire \alu/_0122_ ;
 wire \alu/_0123_ ;
 wire \alu/_0124_ ;
 wire \alu/_0125_ ;
 wire \alu/_0126_ ;
 wire \alu/_0127_ ;
 wire \alu/_0128_ ;
 wire \alu/_0129_ ;
 wire \alu/_0130_ ;
 wire \alu/_0131_ ;
 wire \alu/_0132_ ;
 wire \alu/_0133_ ;
 wire \alu/_0134_ ;
 wire \alu/_0135_ ;
 wire \alu/_0136_ ;
 wire \alu/_0137_ ;
 wire \alu/_0138_ ;
 wire \alu/_0139_ ;
 wire \alu/_0140_ ;
 wire \alu/_0141_ ;
 wire \alu/_0142_ ;
 wire \alu/_0143_ ;
 wire \alu/_0144_ ;
 wire \alu/_0145_ ;
 wire \alu/_0146_ ;
 wire \alu/_0147_ ;
 wire \alu/_0148_ ;
 wire \alu/_0149_ ;
 wire \alu/_0150_ ;
 wire \alu/_0151_ ;
 wire \alu/_0152_ ;
 wire \alu/_0153_ ;
 wire \alu/_0154_ ;
 wire \alu/_0155_ ;
 wire \alu/_0156_ ;
 wire \alu/_0157_ ;
 wire \alu/_0158_ ;
 wire \alu/_0159_ ;
 wire \alu/_0160_ ;
 wire \alu/_0161_ ;
 wire \alu/_0162_ ;
 wire \alu/_0163_ ;
 wire \alu/_0164_ ;
 wire \alu/_0165_ ;
 wire \alu/_0166_ ;
 wire \alu/_0167_ ;
 wire \alu/_0168_ ;
 wire \alu/_0169_ ;
 wire \alu/_0170_ ;
 wire \alu/_0171_ ;
 wire \alu/_0172_ ;
 wire \alu/_0173_ ;
 wire \alu/_0174_ ;
 wire \alu/_0175_ ;
 wire \alu/_0176_ ;
 wire \alu/_0177_ ;
 wire \alu/_0178_ ;
 wire \alu/_0179_ ;
 wire \alu/_0180_ ;
 wire \alu/_0181_ ;
 wire \alu/_0182_ ;
 wire \alu/_0183_ ;
 wire \alu/_0184_ ;
 wire \alu/_0185_ ;
 wire \alu/_0186_ ;
 wire \alu/_0187_ ;
 wire \alu/_0188_ ;
 wire \alu/_0189_ ;
 wire \alu/_0190_ ;
 wire \alu/_0191_ ;
 wire \alu/_0192_ ;
 wire \alu/_0193_ ;
 wire \alu/_0194_ ;
 wire \alu/_0195_ ;
 wire \alu/_0196_ ;
 wire \alu/_0197_ ;
 wire \alu/_0198_ ;
 wire \alu/_0199_ ;
 wire \alu/_0200_ ;
 wire \alu/_0201_ ;
 wire \alu/_0202_ ;
 wire \alu/_0203_ ;
 wire \alu/_0204_ ;
 wire \alu/_0205_ ;
 wire \alu/_0206_ ;
 wire \alu/_0207_ ;
 wire \alu/_0208_ ;
 wire \alu/_0209_ ;
 wire \alu/_0210_ ;
 wire \alu/_0211_ ;
 wire \alu/_0212_ ;
 wire \alu/_0213_ ;
 wire \alu/_0214_ ;
 wire \alu/_0215_ ;
 wire \alu/_0216_ ;
 wire \alu/_0217_ ;
 wire \alu/_0218_ ;
 wire \alu/_0219_ ;
 wire \alu/_0220_ ;
 wire \alu/_0221_ ;
 wire \alu/_0222_ ;
 wire \alu/_0223_ ;
 wire \alu/_0224_ ;
 wire \alu/_0225_ ;
 wire \alu/_0226_ ;
 wire \alu/_0227_ ;
 wire \alu/_0228_ ;
 wire \alu/_0229_ ;
 wire \alu/_0230_ ;
 wire \alu/_0231_ ;
 wire \alu/_0232_ ;
 wire \alu/_0233_ ;
 wire \alu/_0234_ ;
 wire \alu/_0235_ ;
 wire \alu/_0236_ ;
 wire \alu/_0237_ ;
 wire \alu/_0238_ ;
 wire \alu/_0239_ ;
 wire \alu/_0240_ ;
 wire \alu/_0241_ ;
 wire \alu/_0242_ ;
 wire \alu/_0243_ ;
 wire \alu/_0244_ ;
 wire \alu/_0245_ ;
 wire \alu/_0246_ ;
 wire \alu/_0247_ ;
 wire \alu/_0248_ ;
 wire \alu/_0249_ ;
 wire \alu/_0250_ ;
 wire \alu/_0251_ ;
 wire \alu/_0252_ ;
 wire \alu/_0253_ ;
 wire \alu/_0254_ ;
 wire \alu/_0255_ ;
 wire \alu/_0256_ ;
 wire \alu/_0257_ ;
 wire \alu/_0258_ ;
 wire \alu/_0259_ ;
 wire \alu/_0260_ ;
 wire \alu/_0261_ ;
 wire \alu/_0262_ ;
 wire \alu/_0263_ ;
 wire \alu/_0264_ ;
 wire \alu/_0265_ ;
 wire \alu/_0266_ ;
 wire \alu/_0267_ ;
 wire \alu/_0268_ ;
 wire \alu/_0269_ ;
 wire \alu/_0270_ ;
 wire \alu/_0271_ ;
 wire \alu/_0272_ ;
 wire \alu/_0273_ ;
 wire \alu/_0274_ ;
 wire \alu/_0275_ ;
 wire \alu/_0276_ ;
 wire \alu/_0277_ ;
 wire \alu/_0278_ ;
 wire \alu/_0279_ ;
 wire \alu/_0280_ ;
 wire \alu/_0281_ ;
 wire \alu/_0282_ ;
 wire \alu/_0283_ ;
 wire \alu/_0284_ ;
 wire \alu/_0285_ ;
 wire \alu/_0286_ ;
 wire \alu/_0287_ ;
 wire \alu/_0288_ ;
 wire \alu/_0289_ ;
 wire \alu/_0290_ ;
 wire \alu/_0291_ ;
 wire \alu/_0292_ ;
 wire \alu/_0293_ ;
 wire \alu/_0294_ ;
 wire \alu/_0295_ ;
 wire \alu/_0296_ ;
 wire \alu/_0297_ ;
 wire \alu/_0298_ ;
 wire \alu/_0299_ ;
 wire \alu/_0300_ ;
 wire \alu/_0301_ ;
 wire \alu/_0302_ ;
 wire \alu/_0303_ ;
 wire \alu/_0304_ ;
 wire \alu/_0305_ ;
 wire \alu/_0306_ ;
 wire \alu/_0307_ ;
 wire \alu/_0308_ ;
 wire \alu/_0309_ ;
 wire \alu/_0310_ ;
 wire \alu/_0311_ ;
 wire \alu/_0312_ ;
 wire \alu/_0313_ ;
 wire \alu/_0314_ ;
 wire \alu/_0315_ ;
 wire \alu/_0316_ ;
 wire \alu/_0317_ ;
 wire \alu/_0318_ ;
 wire \alu/_0319_ ;
 wire \alu/_0320_ ;
 wire \alu/_0321_ ;
 wire \alu/_0322_ ;
 wire \alu/_0323_ ;
 wire \alu/_0324_ ;
 wire \alu/_0325_ ;
 wire \alu/_0326_ ;
 wire \alu/_0327_ ;
 wire \alu/_0328_ ;
 wire \alu/_0329_ ;
 wire \alu/_0330_ ;
 wire \alu/_0331_ ;
 wire \alu/_0332_ ;
 wire \alu/_0333_ ;
 wire \alu/_0334_ ;
 wire \alu/_0335_ ;
 wire \alu/_0336_ ;
 wire \alu/_0337_ ;
 wire \alu/_0338_ ;
 wire \alu/_0339_ ;
 wire \alu/_0340_ ;
 wire \alu/_0341_ ;
 wire \alu/_0342_ ;
 wire \alu/_0343_ ;
 wire \alu/_0344_ ;
 wire \alu/_0345_ ;
 wire \alu/_0346_ ;
 wire \alu/_0347_ ;
 wire \alu/_0348_ ;
 wire \alu/_0349_ ;
 wire \alu/_0350_ ;
 wire \alu/_0351_ ;
 wire \alu/_0352_ ;
 wire \alu/_0353_ ;
 wire \alu/_0354_ ;
 wire \alu/_0355_ ;
 wire \alu/_0356_ ;
 wire \alu/_0357_ ;
 wire \alu/_0358_ ;
 wire \alu/_0359_ ;
 wire \alu/_0360_ ;
 wire \alu/_0361_ ;
 wire \alu/_0362_ ;
 wire \alu/_0363_ ;
 wire \alu/_0364_ ;
 wire \alu/_0365_ ;
 wire \alu/_0366_ ;
 wire \alu/_0367_ ;
 wire \alu/_0368_ ;
 wire \alu/_0369_ ;
 wire \alu/_0370_ ;
 wire \alu/_0371_ ;
 wire \alu/_0372_ ;
 wire \alu/_0373_ ;
 wire \alu/_0374_ ;
 wire \alu/_0375_ ;
 wire \alu/_0376_ ;
 wire \alu/_0377_ ;
 wire \alu/_0378_ ;
 wire \alu/_0379_ ;
 wire \alu/_0380_ ;
 wire \alu/_0381_ ;
 wire \alu/_0382_ ;
 wire \alu/_0383_ ;
 wire \alu/_0384_ ;
 wire \alu/_0385_ ;
 wire \alu/_0386_ ;
 wire \alu/_0387_ ;
 wire \alu/_0388_ ;
 wire \alu/_0389_ ;
 wire \alu/_0390_ ;
 wire \alu/_0391_ ;
 wire \alu/_0392_ ;
 wire \alu/_0393_ ;
 wire \alu/_0394_ ;
 wire \alu/_0395_ ;
 wire \alu/_0396_ ;
 wire \alu/_0397_ ;
 wire \alu/_0398_ ;
 wire \alu/_0399_ ;
 wire \alu/_0400_ ;
 wire \alu/_0401_ ;
 wire \alu/_0402_ ;
 wire \alu/_0403_ ;
 wire \alu/_0404_ ;
 wire \alu/_0405_ ;
 wire \alu/_0406_ ;
 wire \alu/_0407_ ;
 wire \alu/_0408_ ;
 wire \alu/_0409_ ;
 wire \alu/_0410_ ;
 wire \alu/_0411_ ;
 wire \alu/_0412_ ;
 wire \alu/_0413_ ;
 wire \alu/_0414_ ;
 wire \alu/_0415_ ;
 wire \alu/_0416_ ;
 wire \alu/_0417_ ;
 wire \alu/_0418_ ;
 wire \alu/_0419_ ;
 wire \alu/_0420_ ;
 wire \alu/_0421_ ;
 wire \alu/_0422_ ;
 wire \alu/_0423_ ;
 wire \alu/_0424_ ;
 wire \alu/_0425_ ;
 wire \alu/_0426_ ;
 wire \alu/_0427_ ;
 wire \alu/_0428_ ;
 wire \alu/_0429_ ;
 wire \alu/_0430_ ;
 wire \alu/_0431_ ;
 wire \alu/_0432_ ;
 wire \alu/_0433_ ;
 wire \alu/_0434_ ;
 wire \alu/_0435_ ;
 wire \alu/_0436_ ;
 wire \alu/_0437_ ;
 wire \alu/_0438_ ;
 wire \alu/_0439_ ;
 wire \alu/_0440_ ;
 wire \alu/_0441_ ;
 wire \alu/_0442_ ;
 wire \alu/_0443_ ;
 wire \alu/_0444_ ;
 wire \alu/_0445_ ;
 wire \alu/_0446_ ;
 wire \alu/_0447_ ;
 wire \alu/_0448_ ;
 wire \alu/_0449_ ;
 wire \alu/_0450_ ;
 wire \alu/_0451_ ;
 wire \alu/_0452_ ;
 wire \alu/_0453_ ;
 wire \alu/_0454_ ;
 wire \alu/_0455_ ;
 wire \alu/_0456_ ;
 wire \alu/_0457_ ;
 wire \alu/_0458_ ;
 wire \alu/_0459_ ;
 wire \alu/_0460_ ;
 wire \alu/_0461_ ;
 wire \alu/_0462_ ;
 wire \alu/_0463_ ;
 wire \alu/_0464_ ;
 wire \alu/_0465_ ;
 wire \alu/_0466_ ;
 wire \alu/_0467_ ;
 wire \alu/_0468_ ;
 wire \alu/_0469_ ;
 wire \alu/_0470_ ;
 wire \alu/_0471_ ;
 wire \alu/_0472_ ;
 wire \alu/_0473_ ;
 wire \alu/_0474_ ;
 wire \alu/_0475_ ;
 wire \alu/_0476_ ;
 wire \alu/_0477_ ;
 wire \alu/_0478_ ;
 wire \alu/_0479_ ;
 wire \alu/_0480_ ;
 wire \alu/_0481_ ;
 wire \alu/_0482_ ;
 wire \alu/_0483_ ;
 wire \alu/_0484_ ;
 wire \alu/_0485_ ;
 wire \alu/_0486_ ;
 wire \alu/_0487_ ;
 wire \alu/_0488_ ;
 wire \alu/_0489_ ;
 wire \alu/_0490_ ;
 wire \alu/_0491_ ;
 wire \alu/_0492_ ;
 wire \alu/_0493_ ;
 wire \alu/_0494_ ;
 wire \alu/_0495_ ;
 wire \alu/_0496_ ;
 wire \alu/_0497_ ;
 wire \alu/_0498_ ;
 wire \alu/_0499_ ;
 wire \alu/_0500_ ;
 wire \alu/_0501_ ;
 wire \alu/_0502_ ;
 wire \alu/_0503_ ;
 wire \alu/_0504_ ;
 wire \alu/_0505_ ;
 wire \alu/_0506_ ;
 wire \alu/_0507_ ;
 wire \alu/_0508_ ;
 wire \alu/_0509_ ;
 wire \alu/_0510_ ;
 wire \alu/_0511_ ;
 wire \alu/_0512_ ;
 wire \alu/_0513_ ;
 wire \alu/_0514_ ;
 wire \alu/_0515_ ;
 wire \alu/_0516_ ;
 wire \alu/_0517_ ;
 wire \alu/_0518_ ;
 wire \alu/_0519_ ;
 wire \alu/_0520_ ;
 wire \alu/_0521_ ;
 wire \alu/_0522_ ;
 wire \alu/_0523_ ;
 wire \alu/_0524_ ;
 wire \alu/_0525_ ;
 wire \alu/_0526_ ;
 wire \alu/_0527_ ;
 wire \alu/_0528_ ;
 wire \alu/_0529_ ;
 wire \alu/_0530_ ;
 wire \alu/_0531_ ;
 wire \alu/_0532_ ;
 wire \alu/_0533_ ;
 wire \alu/_0534_ ;
 wire \alu/_0535_ ;
 wire \alu/_0536_ ;
 wire \alu/_0537_ ;
 wire \alu/_0538_ ;
 wire \alu/_0539_ ;
 wire \alu/_0540_ ;
 wire \alu/_0541_ ;
 wire \alu/_0542_ ;
 wire \alu/_0543_ ;
 wire \alu/_0544_ ;
 wire \alu/_0545_ ;
 wire \alu/_0546_ ;
 wire \alu/_0547_ ;
 wire \alu/_0548_ ;
 wire \alu/_0549_ ;
 wire \alu/_0550_ ;
 wire \alu/_0551_ ;
 wire \alu/_0552_ ;
 wire \alu/_0553_ ;
 wire \alu/_0554_ ;
 wire \alu/_0555_ ;
 wire \alu/_0556_ ;
 wire \alu/_0557_ ;
 wire \alu/_0558_ ;
 wire \alu/_0559_ ;
 wire \alu/_0560_ ;
 wire \alu/_0561_ ;
 wire \alu/_0562_ ;
 wire \alu/_0563_ ;
 wire \alu/_0564_ ;
 wire \alu/_0565_ ;
 wire \alu/_0566_ ;
 wire \alu/_0567_ ;
 wire \alu/_0568_ ;
 wire \alu/_0569_ ;
 wire \alu/_0570_ ;
 wire \alu/_0571_ ;
 wire \alu/_0572_ ;
 wire \alu/_0573_ ;
 wire \alu/_0574_ ;
 wire \alu/_0575_ ;
 wire \alu/_0576_ ;
 wire \alu/_0577_ ;
 wire \alu/_0578_ ;
 wire \alu/_0579_ ;
 wire \alu/_0580_ ;
 wire \alu/_0581_ ;
 wire \alu/_0582_ ;
 wire \alu/_0583_ ;
 wire \alu/_0584_ ;
 wire \alu/_0585_ ;
 wire \alu/_0586_ ;
 wire \alu/_0587_ ;
 wire \alu/_0588_ ;
 wire \alu/_0589_ ;
 wire \alu/_0590_ ;
 wire \alu/_0591_ ;
 wire \alu/_0592_ ;
 wire \alu/_0593_ ;
 wire \alu/_0594_ ;
 wire \alu/_0595_ ;
 wire \alu/_0596_ ;
 wire \alu/_0597_ ;
 wire \alu/_0598_ ;
 wire \alu/_0599_ ;
 wire \alu/_0600_ ;
 wire \alu/_0601_ ;
 wire \alu/_0602_ ;
 wire \alu/_0603_ ;
 wire \alu/_0604_ ;
 wire \alu/_0605_ ;
 wire \alu/_0606_ ;
 wire \alu/_0607_ ;
 wire \alu/_0608_ ;
 wire \alu/_0609_ ;
 wire \alu/_0610_ ;
 wire \alu/_0611_ ;
 wire \alu/_0612_ ;
 wire \alu/_0613_ ;
 wire \alu/_0614_ ;
 wire \alu/_0615_ ;
 wire \alu/_0616_ ;
 wire \alu/_0617_ ;
 wire \alu/_0618_ ;
 wire \alu/_0619_ ;
 wire \alu/_0620_ ;
 wire \alu/_0621_ ;
 wire \alu/_0622_ ;
 wire \alu/_0623_ ;
 wire \alu/_0624_ ;
 wire \alu/_0625_ ;
 wire \alu/_0626_ ;
 wire \alu/_0627_ ;
 wire \alu/_0628_ ;
 wire \alu/_0629_ ;
 wire \alu/_0630_ ;
 wire \alu/_0631_ ;
 wire \alu/_0632_ ;
 wire \alu/_0633_ ;
 wire \alu/_0634_ ;
 wire \alu/_0635_ ;
 wire \alu/_0636_ ;
 wire \alu/_0637_ ;
 wire \alu/_0638_ ;
 wire \alu/_0639_ ;
 wire \alu/_0640_ ;
 wire \alu/_0641_ ;
 wire \alu/_0642_ ;
 wire \alu/_0643_ ;
 wire \alu/_0644_ ;
 wire \alu/_0645_ ;
 wire \alu/_0646_ ;
 wire \alu/_0647_ ;
 wire \alu/_0648_ ;
 wire \alu/_0649_ ;
 wire \alu/_0650_ ;
 wire \alu/_0651_ ;
 wire \alu/_0652_ ;
 wire \alu/_0653_ ;
 wire \alu/_0654_ ;
 wire \alu/_0655_ ;
 wire \alu/_0656_ ;
 wire \alu/_0657_ ;
 wire \alu/_0658_ ;
 wire \alu/_0659_ ;
 wire \alu/_0660_ ;
 wire \alu/_0661_ ;
 wire \alu/_0662_ ;
 wire \alu/_0663_ ;
 wire \alu/_0664_ ;
 wire \alu/_0665_ ;
 wire \alu/_0666_ ;
 wire \alu/_0667_ ;
 wire \alu/_0668_ ;
 wire \alu/_0669_ ;
 wire \alu/_0670_ ;
 wire \alu/_0671_ ;
 wire \alu/_0672_ ;
 wire \alu/_0673_ ;
 wire \alu/_0674_ ;
 wire \alu/_0675_ ;
 wire \alu/_0676_ ;
 wire \alu/_0677_ ;
 wire \alu/_0678_ ;
 wire \alu/_0679_ ;
 wire \alu/_0680_ ;
 wire \alu/_0681_ ;
 wire \alu/_0682_ ;
 wire \alu/_0683_ ;
 wire \alu/_0684_ ;
 wire \alu/_0685_ ;
 wire \alu/_0686_ ;
 wire \alu/_0687_ ;
 wire \alu/_0688_ ;
 wire \alu/_0689_ ;
 wire \alu/_0690_ ;
 wire \alu/_0691_ ;
 wire \alu/_0692_ ;
 wire \alu/_0693_ ;
 wire \alu/_0694_ ;
 wire \alu/_0695_ ;
 wire \alu/_0696_ ;
 wire \alu/_0697_ ;
 wire \alu/_0698_ ;
 wire \alu/_0699_ ;
 wire \alu/_0700_ ;
 wire \alu/_0701_ ;
 wire \alu/_0702_ ;
 wire \alu/_0703_ ;
 wire \alu/_0704_ ;
 wire \alu/_0705_ ;
 wire \alu/_0706_ ;
 wire \alu/_0707_ ;
 wire \alu/_0708_ ;
 wire \alu/_0709_ ;
 wire \alu/_0710_ ;
 wire \alu/_0711_ ;
 wire \alu/_0712_ ;
 wire \alu/_0713_ ;
 wire \alu/_0714_ ;
 wire \alu/_0715_ ;
 wire \alu/_0716_ ;
 wire \alu/_0717_ ;
 wire \alu/_0718_ ;
 wire \alu/_0719_ ;
 wire \alu/_0720_ ;
 wire \alu/_0721_ ;
 wire \alu/_0722_ ;
 wire \alu/_0723_ ;
 wire \alu/_0724_ ;
 wire \alu/_0725_ ;
 wire \alu/_0726_ ;
 wire \alu/_0727_ ;
 wire \alu/_0728_ ;
 wire \alu/_0729_ ;
 wire \alu/_0730_ ;
 wire \alu/_0731_ ;
 wire \alu/_0732_ ;
 wire \alu/_0733_ ;
 wire \alu/_0734_ ;
 wire \alu/_0735_ ;
 wire \alu/_0736_ ;
 wire \alu/_0737_ ;
 wire \alu/_0738_ ;
 wire \alu/_0739_ ;
 wire \alu/_0740_ ;
 wire \alu/_0741_ ;
 wire \alu/_0742_ ;
 wire \alu/_0743_ ;
 wire \alu/_0744_ ;
 wire \alu/_0745_ ;
 wire \alu/_0746_ ;
 wire \alu/_0747_ ;
 wire \alu/_0748_ ;
 wire \alu/_0749_ ;
 wire \alu/_0750_ ;
 wire \alu/_0751_ ;
 wire \alu/_0752_ ;
 wire \alu/_0753_ ;
 wire \alu/_0754_ ;
 wire \alu/_0755_ ;
 wire \alu/_0756_ ;
 wire \alu/_0757_ ;
 wire \alu/_0758_ ;
 wire \alu/_0759_ ;
 wire \alu/_0760_ ;
 wire \alu/_0761_ ;
 wire \alu/_0762_ ;
 wire \alu/_0763_ ;
 wire \alu/_0764_ ;
 wire \alu/_0765_ ;
 wire \alu/_0766_ ;
 wire \alu/_0767_ ;
 wire \alu/_0768_ ;
 wire \alu/_0769_ ;
 wire \alu/_0770_ ;
 wire \alu/_0771_ ;
 wire \alu/_0772_ ;
 wire \alu/_0773_ ;
 wire \alu/_0774_ ;
 wire \alu/_0775_ ;
 wire \alu/_0776_ ;
 wire \alu/_0777_ ;
 wire \alu/_0778_ ;
 wire \alu/_0779_ ;
 wire \alu/_0780_ ;
 wire \alu/_0781_ ;
 wire \alu/_0782_ ;
 wire \alu/_0783_ ;
 wire \alu/_0784_ ;
 wire \alu/_0785_ ;
 wire \alu/_0786_ ;
 wire \alu/_0787_ ;
 wire \alu/_0788_ ;
 wire \alu/_0789_ ;
 wire \alu/_0790_ ;
 wire \alu/_0791_ ;
 wire \alu/_0792_ ;
 wire \alu/_0793_ ;
 wire \alu/_0794_ ;
 wire \alu/_0795_ ;
 wire \alu/_0796_ ;
 wire \alu/_0797_ ;
 wire \alu/_0798_ ;
 wire \alu/_0799_ ;
 wire \alu/_0800_ ;
 wire \alu/_0801_ ;
 wire \alu/_0802_ ;
 wire \alu/_0803_ ;
 wire \alu/_0804_ ;
 wire \alu/_0805_ ;
 wire \alu/_0806_ ;
 wire \alu/_0807_ ;
 wire \alu/_0808_ ;
 wire \alu/_0809_ ;
 wire \alu/_0810_ ;
 wire \alu/_0811_ ;
 wire \alu/_0812_ ;
 wire \alu/_0813_ ;
 wire \alu/_0814_ ;
 wire \alu/_0815_ ;
 wire \alu/_0816_ ;
 wire \alu/_0817_ ;
 wire \alu/_0818_ ;
 wire \alu/_0819_ ;
 wire \alu/_0820_ ;
 wire \alu/_0821_ ;
 wire \alu/_0822_ ;
 wire \alu/_0823_ ;
 wire \alu/_0824_ ;
 wire \alu/_0825_ ;
 wire \alu/_0826_ ;
 wire \alu/_0827_ ;
 wire \alu/_0828_ ;
 wire \alu/_0829_ ;
 wire \alu/_0830_ ;
 wire \alu/_0831_ ;
 wire \alu/_0832_ ;
 wire \alu/_0833_ ;
 wire \alu/_0834_ ;
 wire \alu/_0835_ ;
 wire \alu/_0836_ ;
 wire \alu/_0837_ ;
 wire \alu/_0838_ ;
 wire \alu/_0839_ ;
 wire \alu/_0840_ ;
 wire \alu/_0841_ ;
 wire \alu/_0842_ ;
 wire \alu/_0843_ ;
 wire \alu/_0844_ ;
 wire \alu/_0845_ ;
 wire \alu/_0846_ ;
 wire \alu/_0847_ ;
 wire \alu/_0848_ ;
 wire \alu/_0849_ ;
 wire \alu/_0850_ ;
 wire \alu/_0851_ ;
 wire \alu/_0852_ ;
 wire \alu/_0853_ ;
 wire \alu/_0854_ ;
 wire \alu/_0855_ ;
 wire \alu/_0856_ ;
 wire \alu/_0857_ ;
 wire \alu/_0858_ ;
 wire \alu/_0859_ ;
 wire \alu/_0860_ ;
 wire \alu/_0861_ ;
 wire \alu/_0862_ ;
 wire \alu/_0863_ ;
 wire \alu/_0864_ ;
 wire \alu/_0865_ ;
 wire \alu/_0866_ ;
 wire \alu/_0867_ ;
 wire \alu/_0868_ ;
 wire \alu/_0869_ ;
 wire \alu/_0870_ ;
 wire \alu/_0871_ ;
 wire \alu/_0872_ ;
 wire \alu/_0873_ ;
 wire \alu/_0874_ ;
 wire \alu/_0875_ ;
 wire \alu/_0876_ ;
 wire \alu/_0877_ ;
 wire \alu/_0878_ ;
 wire \alu/_0879_ ;
 wire \alu/_0880_ ;
 wire \alu/_0881_ ;
 wire \alu/_0882_ ;
 wire \alu/_0883_ ;
 wire \alu/_0884_ ;
 wire \alu/_0885_ ;
 wire \alu/_0886_ ;
 wire \alu/_0887_ ;
 wire \alu/_0888_ ;
 wire \alu/_0889_ ;
 wire \alu/_0890_ ;
 wire \alu/_0891_ ;
 wire \alu/_0892_ ;
 wire \alu/_0893_ ;
 wire \alu/_0894_ ;
 wire \alu/_0895_ ;
 wire \alu/_0896_ ;
 wire \alu/_0897_ ;
 wire \alu/_0898_ ;
 wire \alu/_0899_ ;
 wire \alu/_0900_ ;
 wire \alu/_0901_ ;
 wire \alu/_0902_ ;
 wire \alu/_0903_ ;
 wire \alu/_0904_ ;
 wire \alu/_0905_ ;
 wire \alu/_0906_ ;
 wire \alu/_0907_ ;
 wire \alu/_0908_ ;
 wire \alu/_0909_ ;
 wire \alu/_0910_ ;
 wire \alu/_0911_ ;
 wire \alu/_0912_ ;
 wire \alu/_0913_ ;
 wire \alu/_0914_ ;
 wire \alu/_0915_ ;
 wire \alu/_0916_ ;
 wire \alu/_0917_ ;
 wire \alu/_0918_ ;
 wire \alu/_0919_ ;
 wire \alu/_0920_ ;
 wire \alu/_0921_ ;
 wire \alu/_0922_ ;
 wire \alu/_0923_ ;
 wire \alu/_0924_ ;
 wire \alu/_0925_ ;
 wire \alu/_0926_ ;
 wire \alu/_0927_ ;
 wire \alu/_0928_ ;
 wire \alu/_0929_ ;
 wire \alu/_0930_ ;
 wire \alu/_0931_ ;
 wire \alu/_0932_ ;
 wire \alu/_0933_ ;
 wire \alu/_0934_ ;
 wire \alu/_0935_ ;
 wire \alu/_0936_ ;
 wire \alu/_0937_ ;
 wire \alu/_0938_ ;
 wire \alu/_0939_ ;
 wire \alu/_0940_ ;
 wire \alu/_0941_ ;
 wire \alu/_0942_ ;
 wire \alu/_0943_ ;
 wire \alu/_0944_ ;
 wire \alu/_0945_ ;
 wire \alu/_0946_ ;
 wire \alu/_0947_ ;
 wire \alu/_0948_ ;
 wire \alu/_0949_ ;
 wire \alu/_0950_ ;
 wire \alu/_0951_ ;
 wire \alu/_0952_ ;
 wire \alu/_0953_ ;
 wire \alu/_0954_ ;
 wire \alu/_0955_ ;
 wire \alu/_0956_ ;
 wire \alu/_0957_ ;
 wire \alu/_0958_ ;
 wire \alu/_0959_ ;
 wire \alu/_0960_ ;
 wire \alu/_0961_ ;
 wire \alu/_0962_ ;
 wire \alu/_0963_ ;
 wire \alu/_0964_ ;
 wire \alu/_0965_ ;
 wire \alu/_0966_ ;
 wire \alu/_0967_ ;
 wire \alu/_0968_ ;
 wire \alu/_0969_ ;
 wire \alu/_0970_ ;
 wire \alu/_0971_ ;
 wire \alu/_0972_ ;
 wire \alu/_0973_ ;
 wire \alu/_0974_ ;
 wire \alu/_0975_ ;
 wire \alu/_0976_ ;
 wire \alu/_0977_ ;
 wire \alu/_0978_ ;
 wire \alu/_0979_ ;
 wire \alu/_0980_ ;
 wire \alu/_0981_ ;
 wire \alu/_0982_ ;
 wire \alu/_0983_ ;
 wire \alu/_0984_ ;
 wire \alu/_0985_ ;
 wire \alu/_0986_ ;
 wire \alu/_0987_ ;
 wire \alu/_0988_ ;
 wire \alu/_0989_ ;
 wire \alu/_0990_ ;
 wire \alu/_0991_ ;
 wire \alu/_0992_ ;
 wire \alu/_0993_ ;
 wire \alu/_0994_ ;
 wire \alu/_0995_ ;
 wire \alu/_0996_ ;
 wire \alu/_0997_ ;
 wire \alu/_0998_ ;
 wire \alu/_0999_ ;
 wire \alu/_1000_ ;
 wire \alu/_1001_ ;
 wire \alu/_1002_ ;
 wire \alu/_1003_ ;
 wire \alu/_1004_ ;
 wire \alu/_1005_ ;
 wire \alu/_1006_ ;
 wire \alu/_1007_ ;
 wire \alu/_1008_ ;
 wire \alu/_1009_ ;
 wire \alu/_1010_ ;
 wire \alu/_1011_ ;
 wire \alu/_1012_ ;
 wire \alu/_1013_ ;
 wire \alu/_1014_ ;
 wire \alu/_1015_ ;
 wire \alu/_1016_ ;
 wire \alu/_1017_ ;
 wire \alu/_1018_ ;
 wire \alu/_1019_ ;
 wire \alu/_1020_ ;
 wire \alu/_1021_ ;
 wire \alu/_1022_ ;
 wire \alu/_1023_ ;
 wire \alu/_1024_ ;
 wire \alu/_1025_ ;
 wire \alu/_1026_ ;
 wire \alu/_1027_ ;
 wire \alu/_1028_ ;
 wire \alu/_1029_ ;
 wire \alu/_1030_ ;
 wire \alu/_1031_ ;
 wire \alu/_1032_ ;
 wire \alu/_1033_ ;
 wire \alu/_1034_ ;
 wire \alu/_1035_ ;
 wire \alu/_1036_ ;
 wire \alu/_1037_ ;
 wire \alu/_1038_ ;
 wire \alu/_1039_ ;
 wire \alu/_1040_ ;
 wire \alu/_1041_ ;
 wire \alu/_1042_ ;
 wire \alu/_1043_ ;
 wire \alu/_1044_ ;
 wire \alu/_1045_ ;
 wire \alu/_1046_ ;
 wire \alu/_1047_ ;
 wire \alu/_1048_ ;
 wire \alu/_1049_ ;
 wire \alu/_1050_ ;
 wire \alu/_1051_ ;
 wire \alu/_1052_ ;
 wire \alu/_1053_ ;
 wire \alu/_1054_ ;
 wire \alu/_1055_ ;
 wire \alu/_1056_ ;
 wire \alu/_1057_ ;
 wire \alu/_1058_ ;
 wire \alu/_1059_ ;
 wire \alu/_1060_ ;
 wire \alu/_1061_ ;
 wire \alu/_1062_ ;
 wire \alu/_1063_ ;
 wire \alu/_1064_ ;
 wire \alu/_1065_ ;
 wire \alu/_1066_ ;
 wire \alu/_1067_ ;
 wire \alu/_1068_ ;
 wire \alu/_1069_ ;
 wire \alu/_1070_ ;
 wire \alu/_1071_ ;
 wire \alu/_1072_ ;
 wire \alu/_1073_ ;
 wire \alu/_1074_ ;
 wire \alu/_1075_ ;
 wire \alu/_1076_ ;
 wire \alu/_1077_ ;
 wire \alu/_1078_ ;
 wire \alu/_1079_ ;
 wire \alu/_1080_ ;
 wire \alu/_1081_ ;
 wire \alu/_1082_ ;
 wire \alu/_1083_ ;
 wire \alu/_1084_ ;
 wire \alu/_1085_ ;
 wire \alu/_1086_ ;
 wire \alu/_1087_ ;
 wire \alu/_1088_ ;
 wire \alu/_1089_ ;
 wire \alu/_1090_ ;
 wire \alu/_1091_ ;
 wire \alu/_1092_ ;
 wire \alu/_1093_ ;
 wire \alu/_1094_ ;
 wire \alu/_1095_ ;
 wire \alu/_1096_ ;
 wire \alu/_1097_ ;
 wire \alu/_1098_ ;
 wire \alu/_1099_ ;
 wire \alu/_1100_ ;
 wire \alu/_1101_ ;
 wire \alu/_1102_ ;
 wire \alu/_1103_ ;
 wire \alu/_1104_ ;
 wire \alu/_1105_ ;
 wire \alu/_1106_ ;
 wire \alu/_1107_ ;
 wire \alu/_1108_ ;
 wire \alu/_1109_ ;
 wire \alu/_1110_ ;
 wire \alu/_1111_ ;
 wire \alu/_1112_ ;
 wire \alu/_1113_ ;
 wire \alu/_1114_ ;
 wire \alu/_1115_ ;
 wire \alu/_1116_ ;
 wire \alu/_1117_ ;
 wire \alu/_1118_ ;
 wire \alu/_1119_ ;
 wire \alu/_1120_ ;
 wire \alu/_1121_ ;
 wire \alu/_1122_ ;
 wire \alu/_1123_ ;
 wire \alu/_1124_ ;
 wire \alu/_1125_ ;
 wire \alu/_1126_ ;
 wire \alu/_1127_ ;
 wire \alu/_1128_ ;
 wire \alu/_1129_ ;
 wire \alu/_1130_ ;
 wire \alu/_1131_ ;
 wire \alu/_1132_ ;
 wire \alu/_1133_ ;
 wire \alu/_1134_ ;
 wire \alu/_1135_ ;
 wire \alu/_1136_ ;
 wire \alu/_1137_ ;
 wire \alu/_1138_ ;
 wire \alu/_1139_ ;
 wire \alu/_1140_ ;
 wire \alu/_1141_ ;
 wire \alu/_1142_ ;
 wire \alu/_1143_ ;
 wire \alu/_1144_ ;
 wire \alu/_1145_ ;
 wire \alu/_1146_ ;
 wire \alu/_1147_ ;
 wire \alu/_1148_ ;
 wire \alu/_1149_ ;
 wire \alu/_1150_ ;
 wire \alu/_1151_ ;
 wire \alu/_1152_ ;
 wire \alu/_1153_ ;
 wire \alu/_1154_ ;
 wire \alu/_1155_ ;
 wire \alu/_1156_ ;
 wire \alu/_1157_ ;
 wire \alu/_1158_ ;
 wire \alu/_1159_ ;
 wire \alu/_1160_ ;
 wire \alu/_1161_ ;
 wire \alu/_1162_ ;
 wire \alu/_1163_ ;
 wire \alu/_1164_ ;
 wire \alu/_1165_ ;
 wire \alu/_1166_ ;
 wire \alu/_1167_ ;
 wire \alu/_1168_ ;
 wire \alu/_1169_ ;
 wire \alu/_1170_ ;
 wire \alu/_1171_ ;
 wire \alu/_1172_ ;
 wire \alu/_1173_ ;
 wire \alu/_1174_ ;
 wire \alu/_1175_ ;
 wire \alu/_1176_ ;
 wire \alu/_1177_ ;
 wire \alu/_1178_ ;
 wire \alu/_1179_ ;
 wire \alu/_1180_ ;
 wire \alu/_1181_ ;
 wire \alu/_1182_ ;
 wire \alu/_1183_ ;
 wire \alu/_1184_ ;
 wire \alu/_1185_ ;
 wire \alu/_1186_ ;
 wire \alu/_1187_ ;
 wire \alu/_1188_ ;
 wire \alu/_1189_ ;
 wire \alu/_1190_ ;
 wire \alu/_1191_ ;
 wire \alu/_1192_ ;
 wire \alu/_1193_ ;
 wire \alu/_1194_ ;
 wire \alu/_1195_ ;
 wire \alu/_1196_ ;
 wire \alu/_1197_ ;
 wire \alu/_1198_ ;
 wire \alu/_1199_ ;
 wire \alu/_1200_ ;
 wire \alu/_1201_ ;
 wire \alu/_1202_ ;
 wire \alu/_1203_ ;
 wire \alu/_1204_ ;
 wire \alu/_1205_ ;
 wire \alu/_1206_ ;
 wire \alu/_1207_ ;
 wire \alu/_1208_ ;
 wire \alu/_1209_ ;
 wire \alu/_1210_ ;
 wire \alu/_1211_ ;
 wire \alu/_1212_ ;
 wire \alu/_1213_ ;
 wire \alu/_1214_ ;
 wire \alu/_1215_ ;
 wire \alu/_1216_ ;
 wire \alu/_1217_ ;
 wire \alu/_1218_ ;
 wire \alu/_1219_ ;
 wire \alu/_1220_ ;
 wire \alu/_1221_ ;
 wire \alu/_1222_ ;
 wire \alu/_1223_ ;
 wire \alu/_1224_ ;
 wire \alu/_1225_ ;
 wire \alu/_1226_ ;
 wire \alu/_1227_ ;
 wire \alu/_1228_ ;
 wire \alu/_1229_ ;
 wire \alu/_1230_ ;
 wire \alu/_1231_ ;
 wire \alu/_1232_ ;
 wire \alu/_1233_ ;
 wire \alu/_1234_ ;
 wire \alu/_1235_ ;
 wire \alu/_1236_ ;
 wire \alu/_1237_ ;
 wire \alu/_1238_ ;
 wire \alu/_1239_ ;
 wire \alu/_1240_ ;
 wire \alu/_1241_ ;
 wire \alu/_1242_ ;
 wire \alu/_1243_ ;
 wire \alu/_1244_ ;
 wire \alu/_1245_ ;
 wire \alu/_1246_ ;
 wire \alu/_1247_ ;
 wire \alu/_1248_ ;
 wire \alu/_1249_ ;
 wire \alu/_1250_ ;
 wire \alu/_1251_ ;
 wire \alu/_1252_ ;
 wire \alu/_1253_ ;
 wire \alu/_1254_ ;
 wire \alu/_1255_ ;
 wire \alu/_1256_ ;
 wire \alu/_1257_ ;
 wire \alu/_1258_ ;
 wire \alu/_1259_ ;
 wire \alu/_1260_ ;
 wire \alu/_1261_ ;
 wire \alu/_1262_ ;
 wire \alu/_1263_ ;
 wire \alu/_1264_ ;
 wire \alu/_1265_ ;
 wire \alu/_1266_ ;
 wire \alu/_1267_ ;
 wire \alu/_1268_ ;
 wire \alu/_1269_ ;
 wire \alu/_1270_ ;
 wire \alu/_1271_ ;
 wire \alu/_1272_ ;
 wire \alu/_1273_ ;
 wire \alu/_1274_ ;
 wire \alu/_1275_ ;
 wire \alu/_1276_ ;
 wire \alu/_1277_ ;
 wire \alu/_1278_ ;
 wire \alu/_1279_ ;
 wire \alu/_1280_ ;
 wire \alu/_1281_ ;
 wire \alu/_1282_ ;
 wire \alu/_1283_ ;
 wire \alu/_1284_ ;
 wire \alu/_1285_ ;
 wire \alu/_1286_ ;
 wire \alu/_1287_ ;
 wire \alu/_1288_ ;
 wire \alu/_1289_ ;
 wire \alu/_1290_ ;
 wire \alu/_1291_ ;
 wire \alu/_1292_ ;
 wire \alu/_1293_ ;
 wire \alu/_1294_ ;
 wire \alu/_1295_ ;
 wire \alu/_1296_ ;
 wire \alu/_1297_ ;
 wire \alu/_1298_ ;
 wire \alu/_1299_ ;
 wire \alu/_1300_ ;
 wire \alu/_1301_ ;
 wire \alu/_1302_ ;
 wire \alu/_1303_ ;
 wire \alu/_1304_ ;
 wire \alu/_1305_ ;
 wire \alu/_1306_ ;
 wire \alu/_1307_ ;
 wire \alu/_1308_ ;
 wire \alu/_1309_ ;
 wire \alu/_1310_ ;
 wire \alu/_1311_ ;
 wire \alu/_1312_ ;
 wire \alu/_1313_ ;
 wire \alu/_1314_ ;
 wire \alu/_1315_ ;
 wire \alu/_1316_ ;
 wire \alu/_1317_ ;
 wire \alu/_1318_ ;
 wire \alu/_1319_ ;
 wire \alu/_1320_ ;
 wire \alu/_1321_ ;
 wire \alu/_1322_ ;
 wire \alu/_1323_ ;
 wire \alu/_1324_ ;
 wire \alu/_1325_ ;
 wire \alu/_1326_ ;
 wire \alu/_1327_ ;
 wire \alu/_1328_ ;
 wire \alu/_1329_ ;
 wire \alu/_1330_ ;
 wire \alu/_1331_ ;
 wire \alu/_1332_ ;
 wire \alu/_1333_ ;
 wire \alu/_1334_ ;
 wire \alu/_1335_ ;
 wire \alu/_1336_ ;
 wire \alu/_1337_ ;
 wire \alu/_1338_ ;
 wire \alu/_1339_ ;
 wire \alu/_1340_ ;
 wire \brancher/_0000_ ;
 wire \brancher/_0001_ ;
 wire \brancher/_0002_ ;
 wire \brancher/_0003_ ;
 wire \brancher/_0004_ ;
 wire \brancher/_0005_ ;
 wire \brancher/_0006_ ;
 wire \brancher/_0007_ ;
 wire \brancher/_0008_ ;
 wire \brancher/_0009_ ;
 wire \brancher/_0010_ ;
 wire \brancher/_0011_ ;
 wire \brancher/_0012_ ;
 wire \brancher/_0013_ ;
 wire \brancher/_0014_ ;
 wire \brancher/_0015_ ;
 wire \brancher/_0016_ ;
 wire \brancher/_0017_ ;
 wire \brancher/_0018_ ;
 wire \brancher/_0019_ ;
 wire \brancher/_0020_ ;
 wire \brancher/_0021_ ;
 wire \brancher/_0022_ ;
 wire \brancher/_0023_ ;
 wire \brancher/_0024_ ;
 wire \brancher/_0025_ ;
 wire \brancher/_0026_ ;
 wire \brancher/_0027_ ;
 wire \brancher/_0028_ ;
 wire \brancher/_0029_ ;
 wire \brancher/_0030_ ;
 wire \brancher/_0031_ ;
 wire \brancher/_0032_ ;
 wire \brancher/_0033_ ;
 wire \brancher/_0034_ ;
 wire \brancher/_0035_ ;
 wire \brancher/_0036_ ;
 wire \brancher/_0037_ ;
 wire \brancher/_0038_ ;
 wire \brancher/_0039_ ;
 wire \brancher/_0040_ ;
 wire \brancher/_0041_ ;
 wire \brancher/_0042_ ;
 wire \brancher/_0043_ ;
 wire \brancher/_0044_ ;
 wire \brancher/_0045_ ;
 wire \brancher/_0046_ ;
 wire \brancher/_0047_ ;
 wire \brancher/_0048_ ;
 wire \brancher/_0049_ ;
 wire \brancher/_0050_ ;
 wire \brancher/_0051_ ;
 wire \brancher/_0052_ ;
 wire \brancher/_0053_ ;
 wire \brancher/_0054_ ;
 wire \brancher/_0055_ ;
 wire \brancher/_0056_ ;
 wire \brancher/_0057_ ;
 wire \brancher/_0058_ ;
 wire \brancher/_0059_ ;
 wire \brancher/_0060_ ;
 wire \brancher/_0061_ ;
 wire \brancher/_0062_ ;
 wire \brancher/_0063_ ;
 wire \brancher/_0064_ ;
 wire \brancher/_0065_ ;
 wire \brancher/_0066_ ;
 wire \brancher/_0067_ ;
 wire \brancher/_0068_ ;
 wire \brancher/_0069_ ;
 wire \brancher/_0070_ ;
 wire \brancher/_0071_ ;
 wire \brancher/_0072_ ;
 wire \brancher/_0073_ ;
 wire \brancher/_0074_ ;
 wire \brancher/_0075_ ;
 wire \brancher/_0076_ ;
 wire \brancher/_0077_ ;
 wire \brancher/_0078_ ;
 wire \brancher/_0079_ ;
 wire \brancher/_0080_ ;
 wire \brancher/_0081_ ;
 wire \brancher/_0082_ ;
 wire \brancher/_0083_ ;
 wire \brancher/_0084_ ;
 wire \brancher/_0085_ ;
 wire \brancher/_0086_ ;
 wire \brancher/_0087_ ;
 wire \brancher/_0088_ ;
 wire \brancher/_0089_ ;
 wire \brancher/_0090_ ;
 wire \brancher/_0091_ ;
 wire \brancher/_0092_ ;
 wire \brancher/_0093_ ;
 wire \brancher/_0094_ ;
 wire \brancher/_0095_ ;
 wire \brancher/_0096_ ;
 wire \brancher/_0097_ ;
 wire \brancher/_0098_ ;
 wire \brancher/_0099_ ;
 wire \brancher/_0100_ ;
 wire \brancher/_0101_ ;
 wire \brancher/_0102_ ;
 wire \brancher/_0103_ ;
 wire \brancher/_0104_ ;
 wire \brancher/_0105_ ;
 wire \brancher/_0106_ ;
 wire \brancher/_0107_ ;
 wire \brancher/_0108_ ;
 wire \brancher/_0109_ ;
 wire \brancher/_0110_ ;
 wire \brancher/_0111_ ;
 wire \brancher/_0112_ ;
 wire \brancher/_0113_ ;
 wire \brancher/_0114_ ;
 wire \brancher/_0115_ ;
 wire \brancher/_0116_ ;
 wire \brancher/_0117_ ;
 wire \brancher/_0118_ ;
 wire \brancher/_0119_ ;
 wire \brancher/_0120_ ;
 wire \brancher/_0121_ ;
 wire \brancher/_0122_ ;
 wire \brancher/_0123_ ;
 wire \brancher/_0124_ ;
 wire \brancher/_0125_ ;
 wire \brancher/_0126_ ;
 wire \brancher/_0127_ ;
 wire \brancher/_0128_ ;
 wire \brancher/_0129_ ;
 wire \brancher/_0130_ ;
 wire \brancher/_0131_ ;
 wire \brancher/_0132_ ;
 wire \brancher/_0133_ ;
 wire \brancher/_0134_ ;
 wire \brancher/_0135_ ;
 wire \brancher/_0136_ ;
 wire \brancher/_0137_ ;
 wire \brancher/_0138_ ;
 wire \brancher/_0139_ ;
 wire \brancher/_0140_ ;
 wire \brancher/_0141_ ;
 wire \brancher/_0142_ ;
 wire \brancher/_0143_ ;
 wire \brancher/_0144_ ;
 wire \brancher/_0145_ ;
 wire \brancher/_0146_ ;
 wire \brancher/_0147_ ;
 wire \brancher/_0148_ ;
 wire \brancher/_0149_ ;
 wire \brancher/_0150_ ;
 wire \brancher/_0151_ ;
 wire \brancher/_0152_ ;
 wire \brancher/_0153_ ;
 wire \brancher/_0154_ ;
 wire \brancher/_0155_ ;
 wire \brancher/_0156_ ;
 wire \brancher/_0157_ ;
 wire \brancher/_0158_ ;
 wire \brancher/_0159_ ;
 wire \brancher/_0160_ ;
 wire \brancher/_0161_ ;
 wire \brancher/_0162_ ;
 wire \brancher/_0163_ ;
 wire \brancher/_0164_ ;
 wire \brancher/_0165_ ;
 wire \brancher/_0166_ ;
 wire \brancher/_0167_ ;
 wire \brancher/_0168_ ;
 wire \brancher/_0169_ ;
 wire \brancher/_0170_ ;
 wire \brancher/_0171_ ;
 wire \brancher/_0172_ ;
 wire \brancher/_0173_ ;
 wire \brancher/_0174_ ;
 wire \brancher/_0175_ ;
 wire \brancher/_0176_ ;
 wire \brancher/_0177_ ;
 wire \brancher/_0178_ ;
 wire \brancher/_0179_ ;
 wire \brancher/_0180_ ;
 wire \brancher/_0181_ ;
 wire \brancher/_0182_ ;
 wire \brancher/_0183_ ;
 wire \brancher/_0184_ ;
 wire \brancher/_0185_ ;
 wire \brancher/_0186_ ;
 wire \brancher/_0187_ ;
 wire \brancher/_0188_ ;
 wire \brancher/_0189_ ;
 wire \brancher/_0190_ ;
 wire \brancher/_0191_ ;
 wire \brancher/_0192_ ;
 wire \brancher/_0193_ ;
 wire \brancher/_0194_ ;
 wire \brancher/_0195_ ;
 wire \brancher/_0196_ ;
 wire \brancher/_0197_ ;
 wire \brancher/_0198_ ;
 wire \brancher/_0199_ ;
 wire \brancher/_0200_ ;
 wire \brancher/_0201_ ;
 wire \brancher/_0202_ ;
 wire \brancher/_0203_ ;
 wire \brancher/_0204_ ;
 wire \brancher/_0205_ ;
 wire \brancher/_0206_ ;
 wire \brancher/_0207_ ;
 wire \brancher/_0208_ ;
 wire \brancher/_0209_ ;
 wire \brancher/_0210_ ;
 wire \brancher/_0211_ ;
 wire \brancher/_0212_ ;
 wire \brancher/_0213_ ;
 wire \brancher/_0214_ ;
 wire \brancher/_0215_ ;
 wire \brancher/_0216_ ;
 wire \brancher/_0217_ ;
 wire \brancher/_0218_ ;
 wire \brancher/_0219_ ;
 wire \brancher/_0220_ ;
 wire \brancher/_0221_ ;
 wire \brancher/_0222_ ;
 wire \brancher/_0223_ ;
 wire \brancher/_0224_ ;
 wire \brancher/_0225_ ;
 wire \brancher/_0226_ ;
 wire \brancher/_0227_ ;
 wire \brancher/_0228_ ;
 wire \brancher/_0229_ ;
 wire \brancher/_0230_ ;
 wire \brancher/_0231_ ;
 wire \brancher/_0232_ ;
 wire \brancher/_0233_ ;
 wire \brancher/_0234_ ;
 wire \brancher/_0235_ ;
 wire \brancher/_0236_ ;
 wire \brancher/_0237_ ;
 wire \brancher/_0238_ ;
 wire \brancher/_0239_ ;
 wire \brancher/_0240_ ;
 wire \brancher/_0241_ ;
 wire \brancher/_0242_ ;
 wire \brancher/_0243_ ;
 wire \brancher/_0244_ ;
 wire \brancher/_0245_ ;
 wire \brancher/_0246_ ;
 wire \brancher/_0247_ ;
 wire \brancher/_0248_ ;
 wire \brancher/_0249_ ;
 wire \brancher/_0250_ ;
 wire \brancher/_0251_ ;
 wire \brancher/_0252_ ;
 wire \brancher/_0253_ ;
 wire \brancher/_0254_ ;
 wire \brancher/_0255_ ;
 wire \brancher/_0256_ ;
 wire \brancher/_0257_ ;
 wire \brancher/_0258_ ;
 wire \brancher/_0259_ ;
 wire \brancher/_0260_ ;
 wire \brancher/_0261_ ;
 wire \brancher/_0262_ ;
 wire \brancher/_0263_ ;
 wire \brancher/_0264_ ;
 wire \brancher/_0265_ ;
 wire \brancher/_0266_ ;
 wire \brancher/_0267_ ;
 wire \brancher/_0268_ ;
 wire \brancher/_0269_ ;
 wire \brancher/_0270_ ;
 wire \brancher/_0271_ ;
 wire \brancher/_0272_ ;
 wire \brancher/_0273_ ;
 wire \brancher/_0274_ ;
 wire \brancher/_0275_ ;
 wire \brancher/_0276_ ;
 wire \brancher/_0277_ ;
 wire \brancher/_0278_ ;
 wire \brancher/_0279_ ;
 wire \brancher/_0280_ ;
 wire \brancher/_0281_ ;
 wire \brancher/_0282_ ;
 wire \brancher/_0283_ ;
 wire \brancher/_0284_ ;
 wire \brancher/_0285_ ;
 wire \brancher/_0286_ ;
 wire \brancher/_0287_ ;
 wire \brancher/_0288_ ;
 wire \brancher/_0289_ ;
 wire \brancher/_0290_ ;
 wire \brancher/_0291_ ;
 wire \brancher/_0292_ ;
 wire \brancher/_0293_ ;
 wire \brancher/_0294_ ;
 wire \brancher/_0295_ ;
 wire \brancher/_0296_ ;
 wire \brancher/_0297_ ;
 wire \brancher/_0298_ ;
 wire \brancher/_0299_ ;
 wire \brancher/_0300_ ;
 wire \brancher/_0301_ ;
 wire \brancher/_0302_ ;
 wire \brancher/_0303_ ;
 wire \brancher/_0304_ ;
 wire \brancher/_0305_ ;
 wire \brancher/_0306_ ;
 wire \brancher/_0307_ ;
 wire \brancher/_0308_ ;
 wire \brancher/_0309_ ;
 wire \brancher/_0310_ ;
 wire \brancher/_0311_ ;
 wire \brancher/_0312_ ;
 wire \brancher/_0313_ ;
 wire \brancher/_0314_ ;
 wire \brancher/_0315_ ;
 wire \brancher/_0316_ ;
 wire \brancher/_0317_ ;
 wire \brancher/_0318_ ;
 wire \brancher/_0319_ ;
 wire \brancher/_0320_ ;
 wire \brancher/_0321_ ;
 wire \brancher/_0322_ ;
 wire \brancher/_0323_ ;
 wire \brancher/_0324_ ;
 wire \brancher/_0325_ ;
 wire \brancher/_0326_ ;
 wire \brancher/_0327_ ;
 wire \brancher/_0328_ ;
 wire \brancher/_0329_ ;
 wire \brancher/_0330_ ;
 wire \brancher/_0331_ ;
 wire \brancher/_0332_ ;
 wire \brancher/_0333_ ;
 wire \brancher/_0334_ ;
 wire \brancher/_0335_ ;
 wire \brancher/_0336_ ;
 wire \brancher/_0337_ ;
 wire \brancher/_0338_ ;
 wire \brancher/_0339_ ;
 wire \brancher/_0340_ ;
 wire \brancher/_0341_ ;
 wire \brancher/_0342_ ;
 wire \brancher/_0343_ ;
 wire \brancher/_0344_ ;
 wire \brancher/_0345_ ;
 wire \brancher/_0346_ ;
 wire \brancher/_0347_ ;
 wire \brancher/_0348_ ;
 wire \brancher/_0349_ ;
 wire \brancher/_0350_ ;
 wire \brancher/_0351_ ;
 wire \brancher/_0352_ ;
 wire \brancher/_0353_ ;
 wire \brancher/_0354_ ;
 wire \brancher/_0355_ ;
 wire \brancher/_0356_ ;
 wire \brancher/_0357_ ;
 wire \brancher/_0358_ ;
 wire \brancher/_0359_ ;
 wire \brancher/_0360_ ;
 wire \brancher/_0361_ ;
 wire \brancher/_0362_ ;
 wire \brancher/_0363_ ;
 wire \brancher/_0364_ ;
 wire \brancher/_0365_ ;
 wire \brancher/_0366_ ;
 wire \brancher/_0367_ ;
 wire \brancher/_0368_ ;
 wire \brancher/_0369_ ;
 wire \brancher/_0370_ ;
 wire \brancher/_0371_ ;
 wire \brancher/_0372_ ;
 wire \brancher/_0373_ ;
 wire \brancher/_0374_ ;
 wire \brancher/_0375_ ;
 wire \brancher/_0376_ ;
 wire \brancher/_0377_ ;
 wire \brancher/_0378_ ;
 wire \brancher/_0379_ ;
 wire \brancher/_0380_ ;
 wire \brancher/_0381_ ;
 wire \brancher/_0382_ ;
 wire \brancher/_0383_ ;
 wire \brancher/_0384_ ;
 wire \brancher/_0385_ ;
 wire \brancher/_0386_ ;
 wire \brancher/_0387_ ;
 wire \brancher/_0388_ ;
 wire \brancher/_0389_ ;
 wire \brancher/_0390_ ;
 wire \brancher/_0391_ ;
 wire \brancher/_0392_ ;
 wire \brancher/_0393_ ;
 wire \brancher/_0394_ ;
 wire \brancher/_0395_ ;
 wire \brancher/_0396_ ;
 wire \brancher/_0397_ ;
 wire \brancher/_0398_ ;
 wire \brancher/_0399_ ;
 wire \brancher/_0400_ ;
 wire \brancher/_0401_ ;
 wire \brancher/_0402_ ;
 wire \brancher/_0403_ ;
 wire \brancher/_0404_ ;
 wire \brancher/_0405_ ;
 wire \brancher/_0406_ ;
 wire \brancher/_0407_ ;
 wire \brancher/_0408_ ;
 wire \brancher/_0409_ ;
 wire \brancher/_0410_ ;
 wire \brancher/_0411_ ;
 wire \brancher/_0412_ ;
 wire \brancher/_0413_ ;
 wire \brancher/_0414_ ;
 wire \brancher/_0415_ ;
 wire \brancher/_0416_ ;
 wire \brancher/_0417_ ;
 wire \brancher/_0418_ ;
 wire \brancher/_0419_ ;
 wire \brancher/_0420_ ;
 wire \brancher/_0421_ ;
 wire \brancher/_0422_ ;
 wire \brancher/_0423_ ;
 wire \brancher/_0424_ ;
 wire \brancher/_0425_ ;
 wire \brancher/_0426_ ;
 wire \brancher/_0427_ ;
 wire \brancher/_0428_ ;
 wire \brancher/_0429_ ;
 wire \brancher/_0430_ ;
 wire \brancher/_0431_ ;
 wire \brancher/_0432_ ;
 wire \brancher/_0433_ ;
 wire \brancher/_0434_ ;
 wire \brancher/_0435_ ;
 wire \brancher/_0436_ ;
 wire \brancher/_0437_ ;
 wire \brancher/_0438_ ;
 wire \brancher/_0439_ ;
 wire \brancher/_0440_ ;
 wire \brancher/_0441_ ;
 wire \brancher/_0442_ ;
 wire \brancher/_0443_ ;
 wire \brancher/_0444_ ;
 wire \brancher/_0445_ ;
 wire \brancher/_0446_ ;
 wire \brancher/_0447_ ;
 wire \brancher/_0448_ ;
 wire \brancher/_0449_ ;
 wire \brancher/_0450_ ;
 wire \brancher/_0451_ ;
 wire \brancher/_0452_ ;
 wire \brancher/_0453_ ;
 wire \brancher/_0454_ ;
 wire \brancher/_0455_ ;
 wire \brancher/_0456_ ;
 wire \brancher/_0457_ ;
 wire \brancher/_0458_ ;
 wire \brancher/_0459_ ;
 wire \brancher/_0460_ ;
 wire \brancher/_0461_ ;
 wire \brancher/_0462_ ;
 wire \brancher/_0463_ ;
 wire \brancher/_0464_ ;
 wire \brancher/_0465_ ;
 wire \brancher/_0466_ ;
 wire \brancher/_0467_ ;
 wire \brancher/_0468_ ;
 wire \brancher/_0469_ ;
 wire \brancher/_0470_ ;
 wire \brancher/_0471_ ;
 wire \brancher/_0472_ ;
 wire \brancher/_0473_ ;
 wire \brancher/_0474_ ;
 wire \brancher/_0475_ ;
 wire \brancher/_0476_ ;
 wire \brancher/_0477_ ;
 wire \brancher/_0478_ ;
 wire \brancher/_0479_ ;
 wire \brancher/_0480_ ;
 wire \brancher/_0481_ ;
 wire \brancher/_0482_ ;
 wire \brancher/_0483_ ;
 wire \brancher/_0484_ ;
 wire \brancher/_0485_ ;
 wire \brancher/_0486_ ;
 wire \brancher/_0487_ ;
 wire \brancher/_0488_ ;
 wire \brancher/_0489_ ;
 wire \brancher/_0490_ ;
 wire \brancher/_0491_ ;
 wire \brancher/_0492_ ;
 wire \brancher/_0493_ ;
 wire \brancher/_0494_ ;
 wire \brancher/_0495_ ;
 wire \brancher/_0496_ ;
 wire \brancher/_0497_ ;
 wire \brancher/_0498_ ;
 wire \brancher/_0499_ ;
 wire \brancher/_0500_ ;
 wire \brancher/_0501_ ;
 wire \brancher/_0502_ ;
 wire \brancher/_0503_ ;
 wire \brancher/_0504_ ;
 wire \brancher/_0505_ ;
 wire \brancher/_0506_ ;
 wire \brancher/_0507_ ;
 wire \brancher/_0508_ ;
 wire \brancher/_0509_ ;
 wire \brancher/_0510_ ;
 wire \brancher/_0511_ ;
 wire \brancher/_0512_ ;
 wire \brancher/_0513_ ;
 wire \brancher/_0514_ ;
 wire \brancher/_0515_ ;
 wire \brancher/_0516_ ;
 wire \brancher/_0517_ ;
 wire \brancher/_0518_ ;
 wire \brancher/_0519_ ;
 wire \brancher/_0520_ ;
 wire \brancher/_0521_ ;
 wire \brancher/_0522_ ;
 wire \brancher/_0523_ ;
 wire \brancher/_0524_ ;
 wire \brancher/_0525_ ;
 wire \brancher/_0526_ ;
 wire \brancher/_0527_ ;
 wire \brancher/_0528_ ;
 wire \brancher/_0529_ ;
 wire \brancher/_0530_ ;
 wire \brancher/_0531_ ;
 wire \brancher/_0532_ ;
 wire \brancher/_0533_ ;
 wire \brancher/_0534_ ;
 wire \brancher/_0535_ ;
 wire \brancher/_0536_ ;
 wire \brancher/_0537_ ;
 wire \brancher/_0538_ ;
 wire \brancher/_0539_ ;
 wire \brancher/_0540_ ;
 wire \brancher/_0541_ ;
 wire \brancher/_0542_ ;
 wire \brancher/_0543_ ;
 wire \brancher/_0544_ ;
 wire \brancher/_0545_ ;
 wire \brancher/_0546_ ;
 wire \brancher/_0547_ ;
 wire \brancher/_0548_ ;
 wire \brancher/_0549_ ;
 wire \brancher/_0550_ ;
 wire \brancher/_0551_ ;
 wire \brancher/_0552_ ;
 wire \brancher/_0553_ ;
 wire \brancher/_0554_ ;
 wire \brancher/_0555_ ;
 wire \brancher/_0556_ ;
 wire \brancher/_0557_ ;
 wire \brancher/_0558_ ;
 wire \brancher/_0559_ ;
 wire \brancher/_0560_ ;
 wire \brancher/_0561_ ;
 wire \brancher/_0562_ ;
 wire \brancher/_0563_ ;
 wire \brancher/_0564_ ;
 wire \brancher/_0565_ ;
 wire \brancher/_0566_ ;
 wire \brancher/_0567_ ;
 wire \brancher/_0568_ ;
 wire \brancher/_0569_ ;
 wire \brancher/_0570_ ;
 wire \brancher/_0571_ ;
 wire \brancher/_0572_ ;
 wire \brancher/_0573_ ;
 wire \brancher/_0574_ ;
 wire \brancher/_0575_ ;
 wire \brancher/_0576_ ;
 wire \brancher/_0577_ ;
 wire \brancher/_0578_ ;
 wire \brancher/_0579_ ;
 wire \brancher/_0580_ ;
 wire \brancher/_0581_ ;
 wire \brancher/_0582_ ;
 wire \brancher/_0583_ ;
 wire \brancher/_0584_ ;
 wire \brancher/_0585_ ;
 wire \brancher/_0586_ ;
 wire \brancher/_0587_ ;
 wire \brancher/_0588_ ;
 wire \brancher/_0589_ ;
 wire \brancher/_0590_ ;
 wire \brancher/_0591_ ;
 wire \brancher/_0592_ ;
 wire \brancher/_0593_ ;
 wire \brancher/_0594_ ;
 wire \brancher/_0595_ ;
 wire \brancher/_0596_ ;
 wire \brancher/_0597_ ;
 wire \brancher/_0598_ ;
 wire \brancher/_0599_ ;
 wire \brancher/_0600_ ;
 wire \brancher/_0601_ ;
 wire \brancher/_0602_ ;
 wire \brancher/_0603_ ;
 wire \brancher/_0604_ ;
 wire \brancher/_0605_ ;
 wire \brancher/_0606_ ;
 wire \brancher/_0607_ ;
 wire \brancher/_0608_ ;
 wire \brancher/_0609_ ;
 wire \brancher/_0610_ ;
 wire \brancher/_0611_ ;
 wire \brancher/_0612_ ;
 wire \brancher/_0613_ ;
 wire \brancher/_0614_ ;
 wire \brancher/_0615_ ;
 wire \brancher/_0616_ ;
 wire \brancher/_0617_ ;
 wire \brancher/_0618_ ;
 wire \brancher/_0619_ ;
 wire \brancher/_0620_ ;
 wire \brancher/_0621_ ;
 wire \brancher/_0622_ ;
 wire \brancher/_0623_ ;
 wire \brancher/_0624_ ;
 wire \brancher/_0625_ ;
 wire \brancher/_0626_ ;
 wire \brancher/_0627_ ;
 wire \brancher/_0628_ ;
 wire \brancher/_0629_ ;
 wire \brancher/_0630_ ;
 wire \brancher/_0631_ ;
 wire \brancher/_0632_ ;
 wire \brancher/_0633_ ;
 wire \brancher/_0634_ ;
 wire \brancher/_0635_ ;
 wire \brancher/_0636_ ;
 wire \brancher/_0637_ ;
 wire \brancher/_0638_ ;
 wire \brancher/_0639_ ;
 wire \brancher/_0640_ ;
 wire \brancher/_0641_ ;
 wire \brancher/_0642_ ;
 wire \brancher/_0643_ ;
 wire \brancher/_0644_ ;
 wire \brancher/_0645_ ;
 wire \brancher/_0646_ ;
 wire \brancher/_0647_ ;
 wire \brancher/_0648_ ;
 wire \brancher/_0649_ ;
 wire \brancher/_0650_ ;
 wire \brancher/_0651_ ;
 wire \brancher/_0652_ ;
 wire \brancher/_0653_ ;
 wire \brancher/_0654_ ;
 wire \brancher/_0655_ ;
 wire \brancher/_0656_ ;
 wire \brancher/_0657_ ;
 wire \brancher/_0658_ ;
 wire \brancher/_0659_ ;
 wire \brancher/_0660_ ;
 wire \brancher/_0661_ ;
 wire \brancher/_0662_ ;
 wire \brancher/_0663_ ;
 wire \brancher/_0664_ ;
 wire \brancher/_0665_ ;
 wire \brancher/_0666_ ;
 wire \brancher/_0667_ ;
 wire \brancher/_0668_ ;
 wire \brancher/_0669_ ;
 wire \brancher/_0670_ ;
 wire \brancher/_0671_ ;
 wire \brancher/_0672_ ;
 wire \brancher/_0673_ ;
 wire \brancher/_0674_ ;
 wire \brancher/_0675_ ;
 wire \brancher/_0676_ ;
 wire \brancher/_0677_ ;
 wire \brancher/_0678_ ;
 wire \brancher/_0679_ ;
 wire \brancher/_0680_ ;
 wire \brancher/_0681_ ;
 wire \brancher/_0682_ ;
 wire \brancher/_0683_ ;
 wire \brancher/_0684_ ;
 wire \brancher/_0685_ ;
 wire \brancher/_0686_ ;
 wire \brancher/_0687_ ;
 wire \brancher/_0688_ ;
 wire \brancher/_0689_ ;
 wire \brancher/_0690_ ;
 wire \brancher/_0691_ ;
 wire \brancher/_0692_ ;
 wire \brancher/_0693_ ;
 wire \brancher/_0694_ ;
 wire \brancher/_0695_ ;
 wire \brancher/_0696_ ;
 wire \brancher/_0697_ ;
 wire \brancher/_0698_ ;
 wire \brancher/_0699_ ;
 wire \brancher/_0700_ ;
 wire \brancher/_0701_ ;
 wire \brancher/_0702_ ;
 wire \brancher/_0703_ ;
 wire \brancher/_0704_ ;
 wire \brancher/_0705_ ;
 wire \brancher/_0706_ ;
 wire \brancher/_0707_ ;
 wire \brancher/_0708_ ;
 wire \brancher/_0709_ ;
 wire \brancher/_0710_ ;
 wire \brancher/_0711_ ;
 wire \brancher/_0712_ ;
 wire \brancher/_0713_ ;
 wire \brancher/_0714_ ;
 wire \brancher/_0715_ ;
 wire \brancher/_0716_ ;
 wire \brancher/_0717_ ;
 wire \brancher/_0718_ ;
 wire \brancher/_0719_ ;
 wire \brancher/_0720_ ;
 wire \brancher/_0721_ ;
 wire \brancher/_0722_ ;
 wire \brancher/_0723_ ;
 wire \brancher/_0724_ ;
 wire \brancher/_0725_ ;
 wire \brancher/_0726_ ;
 wire \brancher/_0727_ ;
 wire \brancher/_0728_ ;
 wire \brancher/_0729_ ;
 wire \brancher/_0730_ ;
 wire \brancher/_0731_ ;
 wire \brancher/_0732_ ;
 wire \brancher/_0733_ ;
 wire \brancher/_0734_ ;
 wire \brancher/_0735_ ;
 wire \brancher/_0736_ ;
 wire \brancher/_0737_ ;
 wire \brancher/_0738_ ;
 wire \brancher/_0739_ ;
 wire \brancher/_0740_ ;
 wire \brancher/_0741_ ;
 wire \brancher/_0742_ ;
 wire \brancher/_0743_ ;
 wire \brancher/_0744_ ;
 wire \brancher/_0745_ ;
 wire \brancher/_0746_ ;
 wire \brancher/_0747_ ;
 wire \brancher/_0748_ ;
 wire \brancher/_0749_ ;
 wire \brancher/_0750_ ;
 wire \brancher/_0751_ ;
 wire \brancher/_0752_ ;
 wire \brancher/_0753_ ;
 wire \brancher/_0754_ ;
 wire \brancher/_0755_ ;
 wire \brancher/_0756_ ;
 wire \brancher/_0757_ ;
 wire \brancher/_0758_ ;
 wire \brancher/_0759_ ;
 wire \brancher/_0760_ ;
 wire \brancher/_0761_ ;
 wire \brancher/_0762_ ;
 wire \brancher/_0763_ ;
 wire \brancher/_0764_ ;
 wire \brancher/_0765_ ;
 wire \brancher/_0766_ ;
 wire \brancher/_0767_ ;
 wire \brancher/_0768_ ;
 wire \brancher/_0769_ ;
 wire \brancher/_0770_ ;
 wire \brancher/_0771_ ;
 wire \brancher/_0772_ ;
 wire \brancher/_0773_ ;
 wire \brancher/_0774_ ;
 wire \brancher/_0775_ ;
 wire \brancher/_0776_ ;
 wire \brancher/_0777_ ;
 wire \brancher/_0778_ ;
 wire \brancher/_0779_ ;
 wire \brancher/_0780_ ;
 wire \brancher/_0781_ ;
 wire \brancher/_0782_ ;
 wire \brancher/_0783_ ;
 wire \brancher/_0784_ ;
 wire \brancher/_0785_ ;
 wire \brancher/_0786_ ;
 wire \brancher/_0787_ ;
 wire \brancher/_0788_ ;
 wire \brancher/_0789_ ;
 wire \brancher/_0790_ ;
 wire \brancher/_0791_ ;
 wire \brancher/_0792_ ;
 wire \brancher/_0793_ ;
 wire \brancher/_0794_ ;
 wire \brancher/_0795_ ;
 wire \brancher/_0796_ ;
 wire \brancher/_0797_ ;
 wire \brancher/_0798_ ;
 wire \brancher/_0799_ ;
 wire \brancher/_0800_ ;
 wire \brancher/_0801_ ;
 wire \brancher/_0802_ ;
 wire \brancher/_0803_ ;
 wire \brancher/_0804_ ;
 wire \brancher/_0805_ ;
 wire \brancher/_0806_ ;
 wire \brancher/_0807_ ;
 wire \brancher/_0808_ ;
 wire \brancher/_0809_ ;
 wire \brancher/_0810_ ;
 wire \brancher/_0811_ ;
 wire \brancher/_0812_ ;
 wire \brancher/_0813_ ;
 wire \brancher/_0814_ ;
 wire \brancher/_0815_ ;
 wire \brancher/_0816_ ;
 wire \brancher/_0817_ ;
 wire \brancher/_0818_ ;
 wire \brancher/_0819_ ;
 wire \brancher/_0820_ ;
 wire \brancher/_0821_ ;
 wire \brancher/_0822_ ;
 wire \brancher/_0823_ ;
 wire \brancher/_0824_ ;
 wire \brancher/_0825_ ;
 wire \brancher/_0826_ ;
 wire \brancher/_0827_ ;
 wire \brancher/_0828_ ;
 wire \brancher/_0829_ ;
 wire \brancher/_0830_ ;
 wire \brancher/_0831_ ;
 wire \brancher/_0832_ ;
 wire \brancher/_0833_ ;
 wire \brancher/_0834_ ;
 wire \brancher/_0835_ ;
 wire \brancher/_0836_ ;
 wire \brancher/_0837_ ;
 wire \brancher/_0838_ ;
 wire \brancher/_0839_ ;
 wire \brancher/_0840_ ;
 wire \brancher/_0841_ ;
 wire \brancher/_0842_ ;
 wire \brancher/_0843_ ;
 wire \brancher/_0844_ ;
 wire \brancher/_0845_ ;
 wire \brancher/_0846_ ;
 wire \brancher/_0847_ ;
 wire \brancher/_0848_ ;
 wire \brancher/_0849_ ;
 wire \brancher/_0850_ ;
 wire \brancher/_0851_ ;
 wire \brancher/_0852_ ;
 wire \brancher/_0853_ ;
 wire \brancher/_0854_ ;
 wire \brancher/_0855_ ;
 wire \brancher/_0856_ ;
 wire \brancher/_0857_ ;
 wire \brancher/_0858_ ;
 wire \brancher/_0859_ ;
 wire \brancher/_0860_ ;
 wire \brancher/_0861_ ;
 wire \brancher/_0862_ ;
 wire \brancher/_0863_ ;
 wire \brancher/_0864_ ;
 wire \brancher/_0865_ ;
 wire \brancher/_0866_ ;
 wire \brancher/_0867_ ;
 wire \brancher/_0868_ ;
 wire \brancher/_0869_ ;
 wire \brancher/_0870_ ;
 wire \brancher/_0871_ ;
 wire \brancher/_0872_ ;
 wire \brancher/_0873_ ;
 wire \brancher/_0874_ ;
 wire \brancher/_0875_ ;
 wire \brancher/_0876_ ;
 wire \brancher/_0877_ ;
 wire \brancher/_0878_ ;
 wire \brancher/_0879_ ;
 wire \brancher/_0880_ ;
 wire \brancher/_0881_ ;
 wire \brancher/_0882_ ;
 wire \brancher/_0883_ ;
 wire \brancher/_0884_ ;
 wire \brancher/_0885_ ;
 wire \brancher/_0886_ ;
 wire \brancher/_0887_ ;
 wire \brancher/_0888_ ;
 wire \brancher/_0889_ ;
 wire \brancher/_0890_ ;
 wire \brancher/_0891_ ;
 wire \brancher/_0892_ ;
 wire \brancher/_0893_ ;
 wire \brancher/_0894_ ;
 wire \brancher/_0895_ ;
 wire \brancher/_0896_ ;
 wire \brancher/_0897_ ;
 wire \brancher/_0898_ ;
 wire \brancher/_0899_ ;
 wire \brancher/_0900_ ;
 wire \brancher/_0901_ ;
 wire \brancher/_0902_ ;
 wire \brancher/_0903_ ;
 wire \brancher/_0904_ ;
 wire \brancher/_0905_ ;
 wire \brancher/_0906_ ;
 wire \brancher/_0907_ ;
 wire \brancher/_0908_ ;
 wire \brancher/_0909_ ;
 wire \brancher/_0910_ ;
 wire \brancher/_0911_ ;
 wire \brancher/_0912_ ;
 wire \brancher/_0913_ ;
 wire \brancher/_0914_ ;
 wire \brancher/_0915_ ;
 wire \brancher/_0916_ ;
 wire \brancher/_0917_ ;
 wire \brancher/_0918_ ;
 wire \brancher/_0919_ ;
 wire \brancher/_0920_ ;
 wire \brancher/_0921_ ;
 wire \brancher/_0922_ ;
 wire \brancher/_0923_ ;
 wire \brancher/_0924_ ;
 wire \brancher/_0925_ ;
 wire \brancher/_0926_ ;
 wire \brancher/_0927_ ;
 wire \brancher/_0928_ ;
 wire \brancher/_0929_ ;
 wire \brancher/_0930_ ;
 wire \brancher/_0931_ ;
 wire \brancher/_0932_ ;
 wire \brancher/_0933_ ;
 wire \brancher/_0934_ ;
 wire \brancher/_0935_ ;
 wire \brancher/_0936_ ;
 wire \brancher/_0937_ ;
 wire \brancher/_0938_ ;
 wire \brancher/_0939_ ;
 wire \brancher/_0940_ ;
 wire \brancher/_0941_ ;
 wire \brancher/_0942_ ;
 wire \brancher/_0943_ ;
 wire \brancher/_0944_ ;
 wire \brancher/_0945_ ;
 wire \brancher/_0946_ ;
 wire \brancher/_0947_ ;
 wire \brancher/_0948_ ;
 wire \brancher/_0949_ ;
 wire \brancher/_0950_ ;
 wire \brancher/_0951_ ;
 wire \brancher/_0952_ ;
 wire \brancher/_0953_ ;
 wire \brancher/_0954_ ;
 wire \brancher/_0955_ ;
 wire \brancher/_0956_ ;
 wire \brancher/_0957_ ;
 wire \brancher/_0958_ ;
 wire \brancher/_0959_ ;
 wire \brancher/_0960_ ;
 wire \brancher/_0961_ ;
 wire \brancher/_0962_ ;
 wire \brancher/_0963_ ;
 wire \brancher/_0964_ ;
 wire \brancher/_0965_ ;
 wire \brancher/_0966_ ;
 wire \brancher/_0967_ ;
 wire \brancher/_0968_ ;
 wire \brancher/_0969_ ;
 wire \brancher/_0970_ ;
 wire \brancher/_0971_ ;
 wire \brancher/_0972_ ;
 wire \brancher/_0973_ ;
 wire \brancher/_0974_ ;
 wire \brancher/_0975_ ;
 wire \brancher/_0976_ ;
 wire \brancher/_0977_ ;
 wire \brancher/_0978_ ;
 wire \brancher/_0979_ ;
 wire \brancher/_0980_ ;
 wire \brancher/_0981_ ;
 wire \brancher/_0982_ ;
 wire \brancher/_0983_ ;
 wire \brancher/_0984_ ;
 wire \brancher/_0985_ ;
 wire \brancher/_0986_ ;
 wire \brancher/_0987_ ;
 wire \brancher/_0988_ ;
 wire \brancher/_0989_ ;
 wire \brancher/_0990_ ;
 wire \brancher/_0991_ ;
 wire \brancher/_0992_ ;
 wire \brancher/_0993_ ;
 wire \brancher/_0994_ ;
 wire \brancher/_0995_ ;
 wire \brancher/_0996_ ;
 wire \brancher/_0997_ ;
 wire \brancher/_0998_ ;
 wire \brancher/_0999_ ;
 wire \brancher/_1000_ ;
 wire \brancher/_1001_ ;
 wire \brancher/_1002_ ;
 wire \brancher/_1003_ ;
 wire \brancher/_1004_ ;
 wire \brancher/_1005_ ;
 wire \brancher/_1006_ ;
 wire \brancher/_1007_ ;
 wire \brancher/_1008_ ;
 wire \brancher/_1009_ ;
 wire \brancher/rAdder_b[10] ;
 wire \brancher/rAdder_b[11] ;
 wire \brancher/rAdder_b[12] ;
 wire \brancher/rAdder_b[13] ;
 wire \brancher/rAdder_b[1] ;
 wire \brancher/rAdder_b[2] ;
 wire \brancher/rAdder_b[3] ;
 wire \brancher/rAdder_b[4] ;
 wire \brancher/rAdder_b[5] ;
 wire \brancher/rAdder_b[6] ;
 wire \brancher/rAdder_b[7] ;
 wire \brancher/rAdder_b[8] ;
 wire \brancher/rAdder_b[9] ;
 wire \brancher/rAdder_jal[10] ;
 wire \brancher/rAdder_jal[11] ;
 wire \brancher/rAdder_jal[12] ;
 wire \brancher/rAdder_jal[13] ;
 wire \brancher/rAdder_jal[14] ;
 wire \brancher/rAdder_jal[15] ;
 wire \brancher/rAdder_jal[16] ;
 wire \brancher/rAdder_jal[17] ;
 wire \brancher/rAdder_jal[18] ;
 wire \brancher/rAdder_jal[19] ;
 wire \brancher/rAdder_jal[1] ;
 wire \brancher/rAdder_jal[20] ;
 wire \brancher/rAdder_jal[21] ;
 wire \brancher/rAdder_jal[2] ;
 wire \brancher/rAdder_jal[3] ;
 wire \brancher/rAdder_jal[4] ;
 wire \brancher/rAdder_jal[5] ;
 wire \brancher/rAdder_jal[6] ;
 wire \brancher/rAdder_jal[7] ;
 wire \brancher/rAdder_jal[8] ;
 wire \brancher/rAdder_jal[9] ;
 wire \brancher/rAlu_result[10] ;
 wire \brancher/rAlu_result[11] ;
 wire \brancher/rAlu_result[12] ;
 wire \brancher/rAlu_result[13] ;
 wire \brancher/rAlu_result[14] ;
 wire \brancher/rAlu_result[15] ;
 wire \brancher/rAlu_result[16] ;
 wire \brancher/rAlu_result[17] ;
 wire \brancher/rAlu_result[18] ;
 wire \brancher/rAlu_result[19] ;
 wire \brancher/rAlu_result[1] ;
 wire \brancher/rAlu_result[20] ;
 wire \brancher/rAlu_result[21] ;
 wire \brancher/rAlu_result[22] ;
 wire \brancher/rAlu_result[23] ;
 wire \brancher/rAlu_result[24] ;
 wire \brancher/rAlu_result[25] ;
 wire \brancher/rAlu_result[26] ;
 wire \brancher/rAlu_result[27] ;
 wire \brancher/rAlu_result[28] ;
 wire \brancher/rAlu_result[29] ;
 wire \brancher/rAlu_result[2] ;
 wire \brancher/rAlu_result[30] ;
 wire \brancher/rAlu_result[31] ;
 wire \brancher/rAlu_result[3] ;
 wire \brancher/rAlu_result[4] ;
 wire \brancher/rAlu_result[5] ;
 wire \brancher/rAlu_result[6] ;
 wire \brancher/rAlu_result[7] ;
 wire \brancher/rAlu_result[8] ;
 wire \brancher/rAlu_result[9] ;
 wire \brancher/rOp_b_type ;
 wire \brancher/rOp_jal ;
 wire \brancher/rOp_jalr ;
 wire \brancher/rPc_current_reg1[0] ;
 wire \brancher/rPc_current_reg1[10] ;
 wire \brancher/rPc_current_reg1[11] ;
 wire \brancher/rPc_current_reg1[12] ;
 wire \brancher/rPc_current_reg1[13] ;
 wire \brancher/rPc_current_reg1[14] ;
 wire \brancher/rPc_current_reg1[15] ;
 wire \brancher/rPc_current_reg1[16] ;
 wire \brancher/rPc_current_reg1[17] ;
 wire \brancher/rPc_current_reg1[18] ;
 wire \brancher/rPc_current_reg1[19] ;
 wire \brancher/rPc_current_reg1[1] ;
 wire \brancher/rPc_current_reg1[20] ;
 wire \brancher/rPc_current_reg1[21] ;
 wire \brancher/rPc_current_reg1[22] ;
 wire \brancher/rPc_current_reg1[23] ;
 wire \brancher/rPc_current_reg1[24] ;
 wire \brancher/rPc_current_reg1[25] ;
 wire \brancher/rPc_current_reg1[26] ;
 wire \brancher/rPc_current_reg1[27] ;
 wire \brancher/rPc_current_reg1[28] ;
 wire \brancher/rPc_current_reg1[29] ;
 wire \brancher/rPc_current_reg1[2] ;
 wire \brancher/rPc_current_reg1[30] ;
 wire \brancher/rPc_current_reg1[31] ;
 wire \brancher/rPc_current_reg1[3] ;
 wire \brancher/rPc_current_reg1[4] ;
 wire \brancher/rPc_current_reg1[5] ;
 wire \brancher/rPc_current_reg1[6] ;
 wire \brancher/rPc_current_reg1[7] ;
 wire \brancher/rPc_current_reg1[8] ;
 wire \brancher/rPc_current_reg1[9] ;
 wire \brancher/rPc_current_reg2[0] ;
 wire \brancher/rPc_current_reg2[10] ;
 wire \brancher/rPc_current_reg2[11] ;
 wire \brancher/rPc_current_reg2[12] ;
 wire \brancher/rPc_current_reg2[13] ;
 wire \brancher/rPc_current_reg2[14] ;
 wire \brancher/rPc_current_reg2[15] ;
 wire \brancher/rPc_current_reg2[16] ;
 wire \brancher/rPc_current_reg2[17] ;
 wire \brancher/rPc_current_reg2[18] ;
 wire \brancher/rPc_current_reg2[19] ;
 wire \brancher/rPc_current_reg2[1] ;
 wire \brancher/rPc_current_reg2[20] ;
 wire \brancher/rPc_current_reg2[21] ;
 wire \brancher/rPc_current_reg2[22] ;
 wire \brancher/rPc_current_reg2[23] ;
 wire \brancher/rPc_current_reg2[24] ;
 wire \brancher/rPc_current_reg2[25] ;
 wire \brancher/rPc_current_reg2[26] ;
 wire \brancher/rPc_current_reg2[27] ;
 wire \brancher/rPc_current_reg2[28] ;
 wire \brancher/rPc_current_reg2[29] ;
 wire \brancher/rPc_current_reg2[2] ;
 wire \brancher/rPc_current_reg2[30] ;
 wire \brancher/rPc_current_reg2[31] ;
 wire \brancher/rPc_current_reg2[3] ;
 wire \brancher/rPc_current_reg2[4] ;
 wire \brancher/rPc_current_reg2[5] ;
 wire \brancher/rPc_current_reg2[6] ;
 wire \brancher/rPc_current_reg2[7] ;
 wire \brancher/rPc_current_reg2[8] ;
 wire \brancher/rPc_current_reg2[9] ;
 wire \brancher/rPc_current_reg3[0] ;
 wire \brancher/rPc_current_reg3[10] ;
 wire \brancher/rPc_current_reg3[11] ;
 wire \brancher/rPc_current_reg3[12] ;
 wire \brancher/rPc_current_reg3[13] ;
 wire \brancher/rPc_current_reg3[14] ;
 wire \brancher/rPc_current_reg3[15] ;
 wire \brancher/rPc_current_reg3[16] ;
 wire \brancher/rPc_current_reg3[17] ;
 wire \brancher/rPc_current_reg3[18] ;
 wire \brancher/rPc_current_reg3[19] ;
 wire \brancher/rPc_current_reg3[1] ;
 wire \brancher/rPc_current_reg3[20] ;
 wire \brancher/rPc_current_reg3[21] ;
 wire \brancher/rPc_current_reg3[22] ;
 wire \brancher/rPc_current_reg3[23] ;
 wire \brancher/rPc_current_reg3[24] ;
 wire \brancher/rPc_current_reg3[25] ;
 wire \brancher/rPc_current_reg3[26] ;
 wire \brancher/rPc_current_reg3[27] ;
 wire \brancher/rPc_current_reg3[28] ;
 wire \brancher/rPc_current_reg3[29] ;
 wire \brancher/rPc_current_reg3[2] ;
 wire \brancher/rPc_current_reg3[30] ;
 wire \brancher/rPc_current_reg3[31] ;
 wire \brancher/rPc_current_reg3[3] ;
 wire \brancher/rPc_current_reg3[4] ;
 wire \brancher/rPc_current_reg3[5] ;
 wire \brancher/rPc_current_reg3[6] ;
 wire \brancher/rPc_current_reg3[7] ;
 wire \brancher/rPc_current_reg3[8] ;
 wire \brancher/rPc_current_reg3[9] ;
 wire \dec/_000_ ;
 wire \dec/_001_ ;
 wire \dec/_002_ ;
 wire \dec/_003_ ;
 wire \dec/_004_ ;
 wire \dec/_005_ ;
 wire \dec/_006_ ;
 wire \dec/_007_ ;
 wire \dec/_008_ ;
 wire \dec/_009_ ;
 wire \dec/_010_ ;
 wire \dec/_011_ ;
 wire \dec/_012_ ;
 wire \dec/_013_ ;
 wire \dec/_014_ ;
 wire \dec/_015_ ;
 wire \dec/_016_ ;
 wire \dec/_017_ ;
 wire \dec/_018_ ;
 wire \dec/_019_ ;
 wire \dec/_020_ ;
 wire \dec/_021_ ;
 wire \dec/_022_ ;
 wire \dec/_023_ ;
 wire \dec/_024_ ;
 wire \dec/_025_ ;
 wire \dec/_026_ ;
 wire \dec/_027_ ;
 wire \dec/_028_ ;
 wire \dec/_029_ ;
 wire \dec/_030_ ;
 wire \dec/_031_ ;
 wire \dec/_032_ ;
 wire \dec/_033_ ;
 wire \dec/_034_ ;
 wire \dec/_035_ ;
 wire \dec/_036_ ;
 wire \dec/_037_ ;
 wire \dec/_038_ ;
 wire \dec/_039_ ;
 wire \dec/_040_ ;
 wire \dec/_041_ ;
 wire \dec/_042_ ;
 wire \dec/_043_ ;
 wire \dec/_044_ ;
 wire \dec/_045_ ;
 wire \dec/_046_ ;
 wire \dec/_047_ ;
 wire \dec/_048_ ;
 wire \dec/_049_ ;
 wire \dec/_050_ ;
 wire \dec/_051_ ;
 wire \dec/_052_ ;
 wire \dec/_053_ ;
 wire \dec/_054_ ;
 wire \dec/_055_ ;
 wire \dec/_056_ ;
 wire \dec/_057_ ;
 wire \dec/_058_ ;
 wire \dec/_059_ ;
 wire \dec/_060_ ;
 wire \dec/_061_ ;
 wire \dec/_062_ ;
 wire \dec/_063_ ;
 wire \dec/_064_ ;
 wire \dec/_065_ ;
 wire \dec/_066_ ;
 wire \dec/_067_ ;
 wire \dec/_068_ ;
 wire \dec/_069_ ;
 wire \dec/_070_ ;
 wire \dec/_071_ ;
 wire \dec/_072_ ;
 wire \dec/_073_ ;
 wire \dec/_074_ ;
 wire \dec/_075_ ;
 wire \dec/_076_ ;
 wire \dec/_077_ ;
 wire \dec/_078_ ;
 wire \dec/_079_ ;
 wire \dec/_080_ ;
 wire \dec/_081_ ;
 wire \dec/_082_ ;
 wire \dec/_083_ ;
 wire \dec/_084_ ;
 wire \dec/_085_ ;
 wire \dec/_086_ ;
 wire \dec/_087_ ;
 wire \dec/_088_ ;
 wire \dec/_089_ ;
 wire \dec/_090_ ;
 wire \dec/_091_ ;
 wire \dec/_092_ ;
 wire \dec/_093_ ;
 wire \dec/_094_ ;
 wire \dec/_095_ ;
 wire \dec/_096_ ;
 wire \dec/_097_ ;
 wire \dec/_098_ ;
 wire \dec/_099_ ;
 wire \dec/_100_ ;
 wire \dec/_101_ ;
 wire \dec/_102_ ;
 wire \dec/_103_ ;
 wire \dec/_104_ ;
 wire \dec/_105_ ;
 wire \dec/_106_ ;
 wire \dec/_107_ ;
 wire \dec/_108_ ;
 wire \dec/_109_ ;
 wire \dec/_110_ ;
 wire \dec/_111_ ;
 wire \dec/_112_ ;
 wire \dec/_113_ ;
 wire \dec/_114_ ;
 wire \dec/_115_ ;
 wire \dec/_116_ ;
 wire \dec/_117_ ;
 wire \dec/_118_ ;
 wire \dec/_119_ ;
 wire \dec/_120_ ;
 wire \dec/_121_ ;
 wire \dec/_122_ ;
 wire \dec/_123_ ;
 wire \dec/_124_ ;
 wire \dec/_125_ ;
 wire \dec/_126_ ;
 wire \dec/_127_ ;
 wire \dec/_128_ ;
 wire \dec/_129_ ;
 wire \dec/_130_ ;
 wire \dec/_131_ ;
 wire \dec/_132_ ;
 wire \dec/_133_ ;
 wire \dec/_134_ ;
 wire \dec/_135_ ;
 wire \dec/_136_ ;
 wire \dec/_137_ ;
 wire \dec/_138_ ;
 wire \dec/_139_ ;
 wire \dec/_140_ ;
 wire \dec/_141_ ;
 wire \dec/_142_ ;
 wire \dec/_143_ ;
 wire \dec/_144_ ;
 wire \dec/_145_ ;
 wire \dec/_146_ ;
 wire \dec/_147_ ;
 wire \dec/_148_ ;
 wire \dec/_149_ ;
 wire \dec/_150_ ;
 wire \dec/_151_ ;
 wire \dec/_152_ ;
 wire \dec/_153_ ;
 wire \dec/_154_ ;
 wire \dec/_155_ ;
 wire \dec/_156_ ;
 wire \dec/_157_ ;
 wire \dec/_158_ ;
 wire \dec/_159_ ;
 wire \dec/_160_ ;
 wire \dec/_161_ ;
 wire \dec/_162_ ;
 wire \dec/_163_ ;
 wire \dec/_164_ ;
 wire \dec/_165_ ;
 wire \dec/_166_ ;
 wire \dec/_167_ ;
 wire \dec/_168_ ;
 wire \dec/_169_ ;
 wire \dec/_170_ ;
 wire \dec/_171_ ;
 wire \dec/_172_ ;
 wire \dec/_173_ ;
 wire \dec/_174_ ;
 wire \dec/_175_ ;
 wire \dec/_176_ ;
 wire \dec/_177_ ;
 wire \dec/_178_ ;
 wire \dec/_179_ ;
 wire \dec/_180_ ;
 wire \dec/_181_ ;
 wire \dec/_182_ ;
 wire \dec/_183_ ;
 wire \dec/_184_ ;
 wire \dec/_185_ ;
 wire \dec/_186_ ;
 wire \dec/_187_ ;
 wire \dec/_188_ ;
 wire \dec/_189_ ;
 wire \dec/_190_ ;
 wire \dec/_191_ ;
 wire \dec/_192_ ;
 wire \dec/_193_ ;
 wire \dec/_194_ ;
 wire \dec/_195_ ;
 wire \dec/_196_ ;
 wire \dec/_197_ ;
 wire \dec/_198_ ;
 wire \dec/_199_ ;
 wire \dec/_200_ ;
 wire \dec/_201_ ;
 wire \dec/_202_ ;
 wire \dec/_203_ ;
 wire \dec/_204_ ;
 wire \dec/_205_ ;
 wire \dec/_206_ ;
 wire \dec/_207_ ;
 wire \dec/_208_ ;
 wire \dec/_209_ ;
 wire \dec/_210_ ;
 wire \dec/_211_ ;
 wire \dec/_212_ ;
 wire \dec/_213_ ;
 wire \dec/_214_ ;
 wire \dec/_215_ ;
 wire \dec/_216_ ;
 wire \dec/_217_ ;
 wire \dec/_218_ ;
 wire \dec/_219_ ;
 wire \dec/_220_ ;
 wire \dec/_221_ ;
 wire \dec/_222_ ;
 wire \dec/_223_ ;
 wire \dec/_224_ ;
 wire \dec/_225_ ;
 wire \dec/_226_ ;
 wire \dec/_227_ ;
 wire \dec/_228_ ;
 wire \dec/_229_ ;
 wire \dec/_230_ ;
 wire \dec/_231_ ;
 wire \dec/_232_ ;
 wire \dec/_233_ ;
 wire \dec/_234_ ;
 wire \dec/_235_ ;
 wire \dec/_236_ ;
 wire \dec/_237_ ;
 wire \dec/_238_ ;
 wire \dec/_239_ ;
 wire \dec/_240_ ;
 wire \dec/_241_ ;
 wire \dec/_242_ ;
 wire \dec/_243_ ;
 wire \dec/_244_ ;
 wire \dec/_245_ ;
 wire \dec/_246_ ;
 wire \dec/_247_ ;
 wire \dec/_248_ ;
 wire \dec/_249_ ;
 wire \dec/_250_ ;
 wire \dec/_251_ ;
 wire \dec/_252_ ;
 wire \dec/_253_ ;
 wire \dec/_254_ ;
 wire \dec/_255_ ;
 wire \dec/_256_ ;
 wire \dec/_257_ ;
 wire \dec/_258_ ;
 wire \dec/_259_ ;
 wire \dec/_260_ ;
 wire \dec/_261_ ;
 wire \dec/_262_ ;
 wire \dec/_263_ ;
 wire \dec/_264_ ;
 wire \dec/_265_ ;
 wire \dec/_266_ ;
 wire \dec/_267_ ;
 wire \dec/_268_ ;
 wire \dec/_269_ ;
 wire \dec/_270_ ;
 wire \dec/_271_ ;
 wire \dec/_272_ ;
 wire \dec/_273_ ;
 wire \dec/_274_ ;
 wire \dec/_275_ ;
 wire \dec/_276_ ;
 wire \dec/_277_ ;
 wire \dec/_278_ ;
 wire \dec/_279_ ;
 wire \dec/_280_ ;
 wire \dec/_281_ ;
 wire \dec/_282_ ;
 wire \dec/_283_ ;
 wire \dec/_284_ ;
 wire \dec/_285_ ;
 wire \dec/_286_ ;
 wire \dec/_287_ ;
 wire \dec/_288_ ;
 wire \dec/_289_ ;
 wire \dec/_290_ ;
 wire \dec/_291_ ;
 wire \dec/_292_ ;
 wire \dec/_293_ ;
 wire \dec/_294_ ;
 wire \dec/_295_ ;
 wire \dec/_296_ ;
 wire \dec/_297_ ;
 wire \dec/_298_ ;
 wire \dec/_299_ ;
 wire \dec/_300_ ;
 wire \dec/rInstrustion1[0] ;
 wire \dec/rInstrustion1[10] ;
 wire \dec/rInstrustion1[11] ;
 wire \dec/rInstrustion1[12] ;
 wire \dec/rInstrustion1[13] ;
 wire \dec/rInstrustion1[14] ;
 wire \dec/rInstrustion1[15] ;
 wire \dec/rInstrustion1[16] ;
 wire \dec/rInstrustion1[17] ;
 wire \dec/rInstrustion1[18] ;
 wire \dec/rInstrustion1[19] ;
 wire \dec/rInstrustion1[1] ;
 wire \dec/rInstrustion1[20] ;
 wire \dec/rInstrustion1[21] ;
 wire \dec/rInstrustion1[22] ;
 wire \dec/rInstrustion1[23] ;
 wire \dec/rInstrustion1[24] ;
 wire \dec/rInstrustion1[25] ;
 wire \dec/rInstrustion1[26] ;
 wire \dec/rInstrustion1[27] ;
 wire \dec/rInstrustion1[28] ;
 wire \dec/rInstrustion1[29] ;
 wire \dec/rInstrustion1[2] ;
 wire \dec/rInstrustion1[30] ;
 wire \dec/rInstrustion1[31] ;
 wire \dec/rInstrustion1[3] ;
 wire \dec/rInstrustion1[4] ;
 wire \dec/rInstrustion1[5] ;
 wire \dec/rInstrustion1[6] ;
 wire \dec/rInstrustion1[7] ;
 wire \dec/rInstrustion1[8] ;
 wire \dec/rInstrustion1[9] ;
 wire \dec/rInstrustion2[0] ;
 wire \dec/rInstrustion2[10] ;
 wire \dec/rInstrustion2[11] ;
 wire \dec/rInstrustion2[12] ;
 wire \dec/rInstrustion2[13] ;
 wire \dec/rInstrustion2[14] ;
 wire \dec/rInstrustion2[15] ;
 wire \dec/rInstrustion2[16] ;
 wire \dec/rInstrustion2[17] ;
 wire \dec/rInstrustion2[18] ;
 wire \dec/rInstrustion2[19] ;
 wire \dec/rInstrustion2[1] ;
 wire \dec/rInstrustion2[20] ;
 wire \dec/rInstrustion2[21] ;
 wire \dec/rInstrustion2[22] ;
 wire \dec/rInstrustion2[23] ;
 wire \dec/rInstrustion2[24] ;
 wire \dec/rInstrustion2[25] ;
 wire \dec/rInstrustion2[26] ;
 wire \dec/rInstrustion2[27] ;
 wire \dec/rInstrustion2[28] ;
 wire \dec/rInstrustion2[29] ;
 wire \dec/rInstrustion2[2] ;
 wire \dec/rInstrustion2[30] ;
 wire \dec/rInstrustion2[31] ;
 wire \dec/rInstrustion2[3] ;
 wire \dec/rInstrustion2[4] ;
 wire \dec/rInstrustion2[5] ;
 wire \dec/rInstrustion2[6] ;
 wire \dec/rInstrustion2[7] ;
 wire \dec/rInstrustion2[8] ;
 wire \dec/rInstrustion2[9] ;
 wire \dec/rStall1 ;
 wire \dec/rStall2 ;
 wire \reg_module/_00000_ ;
 wire \reg_module/_00001_ ;
 wire \reg_module/_00002_ ;
 wire \reg_module/_00003_ ;
 wire \reg_module/_00004_ ;
 wire \reg_module/_00005_ ;
 wire \reg_module/_00006_ ;
 wire \reg_module/_00007_ ;
 wire \reg_module/_00008_ ;
 wire \reg_module/_00009_ ;
 wire \reg_module/_00010_ ;
 wire \reg_module/_00011_ ;
 wire \reg_module/_00012_ ;
 wire \reg_module/_00013_ ;
 wire \reg_module/_00014_ ;
 wire \reg_module/_00015_ ;
 wire \reg_module/_00016_ ;
 wire \reg_module/_00017_ ;
 wire \reg_module/_00018_ ;
 wire \reg_module/_00019_ ;
 wire \reg_module/_00020_ ;
 wire \reg_module/_00021_ ;
 wire \reg_module/_00022_ ;
 wire \reg_module/_00023_ ;
 wire \reg_module/_00024_ ;
 wire \reg_module/_00025_ ;
 wire \reg_module/_00026_ ;
 wire \reg_module/_00027_ ;
 wire \reg_module/_00028_ ;
 wire \reg_module/_00029_ ;
 wire \reg_module/_00030_ ;
 wire \reg_module/_00031_ ;
 wire \reg_module/_00032_ ;
 wire \reg_module/_00033_ ;
 wire \reg_module/_00034_ ;
 wire \reg_module/_00035_ ;
 wire \reg_module/_00036_ ;
 wire \reg_module/_00037_ ;
 wire \reg_module/_00038_ ;
 wire \reg_module/_00039_ ;
 wire \reg_module/_00040_ ;
 wire \reg_module/_00041_ ;
 wire \reg_module/_00042_ ;
 wire \reg_module/_00043_ ;
 wire \reg_module/_00044_ ;
 wire \reg_module/_00045_ ;
 wire \reg_module/_00046_ ;
 wire \reg_module/_00047_ ;
 wire \reg_module/_00048_ ;
 wire \reg_module/_00049_ ;
 wire \reg_module/_00050_ ;
 wire \reg_module/_00051_ ;
 wire \reg_module/_00052_ ;
 wire \reg_module/_00053_ ;
 wire \reg_module/_00054_ ;
 wire \reg_module/_00055_ ;
 wire \reg_module/_00056_ ;
 wire \reg_module/_00057_ ;
 wire \reg_module/_00058_ ;
 wire \reg_module/_00059_ ;
 wire \reg_module/_00060_ ;
 wire \reg_module/_00061_ ;
 wire \reg_module/_00062_ ;
 wire \reg_module/_00063_ ;
 wire \reg_module/_00064_ ;
 wire \reg_module/_00065_ ;
 wire \reg_module/_00066_ ;
 wire \reg_module/_00067_ ;
 wire \reg_module/_00068_ ;
 wire \reg_module/_00069_ ;
 wire \reg_module/_00070_ ;
 wire \reg_module/_00071_ ;
 wire \reg_module/_00072_ ;
 wire \reg_module/_00073_ ;
 wire \reg_module/_00074_ ;
 wire \reg_module/_00075_ ;
 wire \reg_module/_00076_ ;
 wire \reg_module/_00077_ ;
 wire \reg_module/_00078_ ;
 wire \reg_module/_00079_ ;
 wire \reg_module/_00080_ ;
 wire \reg_module/_00081_ ;
 wire \reg_module/_00082_ ;
 wire \reg_module/_00083_ ;
 wire \reg_module/_00084_ ;
 wire \reg_module/_00085_ ;
 wire \reg_module/_00086_ ;
 wire \reg_module/_00087_ ;
 wire \reg_module/_00088_ ;
 wire \reg_module/_00089_ ;
 wire \reg_module/_00090_ ;
 wire \reg_module/_00091_ ;
 wire \reg_module/_00092_ ;
 wire \reg_module/_00093_ ;
 wire \reg_module/_00094_ ;
 wire \reg_module/_00095_ ;
 wire \reg_module/_00096_ ;
 wire \reg_module/_00097_ ;
 wire \reg_module/_00098_ ;
 wire \reg_module/_00099_ ;
 wire \reg_module/_00100_ ;
 wire \reg_module/_00101_ ;
 wire \reg_module/_00102_ ;
 wire \reg_module/_00103_ ;
 wire \reg_module/_00104_ ;
 wire \reg_module/_00105_ ;
 wire \reg_module/_00106_ ;
 wire \reg_module/_00107_ ;
 wire \reg_module/_00108_ ;
 wire \reg_module/_00109_ ;
 wire \reg_module/_00110_ ;
 wire \reg_module/_00111_ ;
 wire \reg_module/_00112_ ;
 wire \reg_module/_00113_ ;
 wire \reg_module/_00114_ ;
 wire \reg_module/_00115_ ;
 wire \reg_module/_00116_ ;
 wire \reg_module/_00117_ ;
 wire \reg_module/_00118_ ;
 wire \reg_module/_00119_ ;
 wire \reg_module/_00120_ ;
 wire \reg_module/_00121_ ;
 wire \reg_module/_00122_ ;
 wire \reg_module/_00123_ ;
 wire \reg_module/_00124_ ;
 wire \reg_module/_00125_ ;
 wire \reg_module/_00126_ ;
 wire \reg_module/_00127_ ;
 wire \reg_module/_00128_ ;
 wire \reg_module/_00129_ ;
 wire \reg_module/_00130_ ;
 wire \reg_module/_00131_ ;
 wire \reg_module/_00132_ ;
 wire \reg_module/_00133_ ;
 wire \reg_module/_00134_ ;
 wire \reg_module/_00135_ ;
 wire \reg_module/_00136_ ;
 wire \reg_module/_00137_ ;
 wire \reg_module/_00138_ ;
 wire \reg_module/_00139_ ;
 wire \reg_module/_00140_ ;
 wire \reg_module/_00141_ ;
 wire \reg_module/_00142_ ;
 wire \reg_module/_00143_ ;
 wire \reg_module/_00144_ ;
 wire \reg_module/_00145_ ;
 wire \reg_module/_00146_ ;
 wire \reg_module/_00147_ ;
 wire \reg_module/_00148_ ;
 wire \reg_module/_00149_ ;
 wire \reg_module/_00150_ ;
 wire \reg_module/_00151_ ;
 wire \reg_module/_00152_ ;
 wire \reg_module/_00153_ ;
 wire \reg_module/_00154_ ;
 wire \reg_module/_00155_ ;
 wire \reg_module/_00156_ ;
 wire \reg_module/_00157_ ;
 wire \reg_module/_00158_ ;
 wire \reg_module/_00159_ ;
 wire \reg_module/_00160_ ;
 wire \reg_module/_00161_ ;
 wire \reg_module/_00162_ ;
 wire \reg_module/_00163_ ;
 wire \reg_module/_00164_ ;
 wire \reg_module/_00165_ ;
 wire \reg_module/_00166_ ;
 wire \reg_module/_00167_ ;
 wire \reg_module/_00168_ ;
 wire \reg_module/_00169_ ;
 wire \reg_module/_00170_ ;
 wire \reg_module/_00171_ ;
 wire \reg_module/_00172_ ;
 wire \reg_module/_00173_ ;
 wire \reg_module/_00174_ ;
 wire \reg_module/_00175_ ;
 wire \reg_module/_00176_ ;
 wire \reg_module/_00177_ ;
 wire \reg_module/_00178_ ;
 wire \reg_module/_00179_ ;
 wire \reg_module/_00180_ ;
 wire \reg_module/_00181_ ;
 wire \reg_module/_00182_ ;
 wire \reg_module/_00183_ ;
 wire \reg_module/_00184_ ;
 wire \reg_module/_00185_ ;
 wire \reg_module/_00186_ ;
 wire \reg_module/_00187_ ;
 wire \reg_module/_00188_ ;
 wire \reg_module/_00189_ ;
 wire \reg_module/_00190_ ;
 wire \reg_module/_00191_ ;
 wire \reg_module/_00192_ ;
 wire \reg_module/_00193_ ;
 wire \reg_module/_00194_ ;
 wire \reg_module/_00195_ ;
 wire \reg_module/_00196_ ;
 wire \reg_module/_00197_ ;
 wire \reg_module/_00198_ ;
 wire \reg_module/_00199_ ;
 wire \reg_module/_00200_ ;
 wire \reg_module/_00201_ ;
 wire \reg_module/_00202_ ;
 wire \reg_module/_00203_ ;
 wire \reg_module/_00204_ ;
 wire \reg_module/_00205_ ;
 wire \reg_module/_00206_ ;
 wire \reg_module/_00207_ ;
 wire \reg_module/_00208_ ;
 wire \reg_module/_00209_ ;
 wire \reg_module/_00210_ ;
 wire \reg_module/_00211_ ;
 wire \reg_module/_00212_ ;
 wire \reg_module/_00213_ ;
 wire \reg_module/_00214_ ;
 wire \reg_module/_00215_ ;
 wire \reg_module/_00216_ ;
 wire \reg_module/_00217_ ;
 wire \reg_module/_00218_ ;
 wire \reg_module/_00219_ ;
 wire \reg_module/_00220_ ;
 wire \reg_module/_00221_ ;
 wire \reg_module/_00222_ ;
 wire \reg_module/_00223_ ;
 wire \reg_module/_00224_ ;
 wire \reg_module/_00225_ ;
 wire \reg_module/_00226_ ;
 wire \reg_module/_00227_ ;
 wire \reg_module/_00228_ ;
 wire \reg_module/_00229_ ;
 wire \reg_module/_00230_ ;
 wire \reg_module/_00231_ ;
 wire \reg_module/_00232_ ;
 wire \reg_module/_00233_ ;
 wire \reg_module/_00234_ ;
 wire \reg_module/_00235_ ;
 wire \reg_module/_00236_ ;
 wire \reg_module/_00237_ ;
 wire \reg_module/_00238_ ;
 wire \reg_module/_00239_ ;
 wire \reg_module/_00240_ ;
 wire \reg_module/_00241_ ;
 wire \reg_module/_00242_ ;
 wire \reg_module/_00243_ ;
 wire \reg_module/_00244_ ;
 wire \reg_module/_00245_ ;
 wire \reg_module/_00246_ ;
 wire \reg_module/_00247_ ;
 wire \reg_module/_00248_ ;
 wire \reg_module/_00249_ ;
 wire \reg_module/_00250_ ;
 wire \reg_module/_00251_ ;
 wire \reg_module/_00252_ ;
 wire \reg_module/_00253_ ;
 wire \reg_module/_00254_ ;
 wire \reg_module/_00255_ ;
 wire \reg_module/_00256_ ;
 wire \reg_module/_00257_ ;
 wire \reg_module/_00258_ ;
 wire \reg_module/_00259_ ;
 wire \reg_module/_00260_ ;
 wire \reg_module/_00261_ ;
 wire \reg_module/_00262_ ;
 wire \reg_module/_00263_ ;
 wire \reg_module/_00264_ ;
 wire \reg_module/_00265_ ;
 wire \reg_module/_00266_ ;
 wire \reg_module/_00267_ ;
 wire \reg_module/_00268_ ;
 wire \reg_module/_00269_ ;
 wire \reg_module/_00270_ ;
 wire \reg_module/_00271_ ;
 wire \reg_module/_00272_ ;
 wire \reg_module/_00273_ ;
 wire \reg_module/_00274_ ;
 wire \reg_module/_00275_ ;
 wire \reg_module/_00276_ ;
 wire \reg_module/_00277_ ;
 wire \reg_module/_00278_ ;
 wire \reg_module/_00279_ ;
 wire \reg_module/_00280_ ;
 wire \reg_module/_00281_ ;
 wire \reg_module/_00282_ ;
 wire \reg_module/_00283_ ;
 wire \reg_module/_00284_ ;
 wire \reg_module/_00285_ ;
 wire \reg_module/_00286_ ;
 wire \reg_module/_00287_ ;
 wire \reg_module/_00288_ ;
 wire \reg_module/_00289_ ;
 wire \reg_module/_00290_ ;
 wire \reg_module/_00291_ ;
 wire \reg_module/_00292_ ;
 wire \reg_module/_00293_ ;
 wire \reg_module/_00294_ ;
 wire \reg_module/_00295_ ;
 wire \reg_module/_00296_ ;
 wire \reg_module/_00297_ ;
 wire \reg_module/_00298_ ;
 wire \reg_module/_00299_ ;
 wire \reg_module/_00300_ ;
 wire \reg_module/_00301_ ;
 wire \reg_module/_00302_ ;
 wire \reg_module/_00303_ ;
 wire \reg_module/_00304_ ;
 wire \reg_module/_00305_ ;
 wire \reg_module/_00306_ ;
 wire \reg_module/_00307_ ;
 wire \reg_module/_00308_ ;
 wire \reg_module/_00309_ ;
 wire \reg_module/_00310_ ;
 wire \reg_module/_00311_ ;
 wire \reg_module/_00312_ ;
 wire \reg_module/_00313_ ;
 wire \reg_module/_00314_ ;
 wire \reg_module/_00315_ ;
 wire \reg_module/_00316_ ;
 wire \reg_module/_00317_ ;
 wire \reg_module/_00318_ ;
 wire \reg_module/_00319_ ;
 wire \reg_module/_00320_ ;
 wire \reg_module/_00321_ ;
 wire \reg_module/_00322_ ;
 wire \reg_module/_00323_ ;
 wire \reg_module/_00324_ ;
 wire \reg_module/_00325_ ;
 wire \reg_module/_00326_ ;
 wire \reg_module/_00327_ ;
 wire \reg_module/_00328_ ;
 wire \reg_module/_00329_ ;
 wire \reg_module/_00330_ ;
 wire \reg_module/_00331_ ;
 wire \reg_module/_00332_ ;
 wire \reg_module/_00333_ ;
 wire \reg_module/_00334_ ;
 wire \reg_module/_00335_ ;
 wire \reg_module/_00336_ ;
 wire \reg_module/_00337_ ;
 wire \reg_module/_00338_ ;
 wire \reg_module/_00339_ ;
 wire \reg_module/_00340_ ;
 wire \reg_module/_00341_ ;
 wire \reg_module/_00342_ ;
 wire \reg_module/_00343_ ;
 wire \reg_module/_00344_ ;
 wire \reg_module/_00345_ ;
 wire \reg_module/_00346_ ;
 wire \reg_module/_00347_ ;
 wire \reg_module/_00348_ ;
 wire \reg_module/_00349_ ;
 wire \reg_module/_00350_ ;
 wire \reg_module/_00351_ ;
 wire \reg_module/_00352_ ;
 wire \reg_module/_00353_ ;
 wire \reg_module/_00354_ ;
 wire \reg_module/_00355_ ;
 wire \reg_module/_00356_ ;
 wire \reg_module/_00357_ ;
 wire \reg_module/_00358_ ;
 wire \reg_module/_00359_ ;
 wire \reg_module/_00360_ ;
 wire \reg_module/_00361_ ;
 wire \reg_module/_00362_ ;
 wire \reg_module/_00363_ ;
 wire \reg_module/_00364_ ;
 wire \reg_module/_00365_ ;
 wire \reg_module/_00366_ ;
 wire \reg_module/_00367_ ;
 wire \reg_module/_00368_ ;
 wire \reg_module/_00369_ ;
 wire \reg_module/_00370_ ;
 wire \reg_module/_00371_ ;
 wire \reg_module/_00372_ ;
 wire \reg_module/_00373_ ;
 wire \reg_module/_00374_ ;
 wire \reg_module/_00375_ ;
 wire \reg_module/_00376_ ;
 wire \reg_module/_00377_ ;
 wire \reg_module/_00378_ ;
 wire \reg_module/_00379_ ;
 wire \reg_module/_00380_ ;
 wire \reg_module/_00381_ ;
 wire \reg_module/_00382_ ;
 wire \reg_module/_00383_ ;
 wire \reg_module/_00384_ ;
 wire \reg_module/_00385_ ;
 wire \reg_module/_00386_ ;
 wire \reg_module/_00387_ ;
 wire \reg_module/_00388_ ;
 wire \reg_module/_00389_ ;
 wire \reg_module/_00390_ ;
 wire \reg_module/_00391_ ;
 wire \reg_module/_00392_ ;
 wire \reg_module/_00393_ ;
 wire \reg_module/_00394_ ;
 wire \reg_module/_00395_ ;
 wire \reg_module/_00396_ ;
 wire \reg_module/_00397_ ;
 wire \reg_module/_00398_ ;
 wire \reg_module/_00399_ ;
 wire \reg_module/_00400_ ;
 wire \reg_module/_00401_ ;
 wire \reg_module/_00402_ ;
 wire \reg_module/_00403_ ;
 wire \reg_module/_00404_ ;
 wire \reg_module/_00405_ ;
 wire \reg_module/_00406_ ;
 wire \reg_module/_00407_ ;
 wire \reg_module/_00408_ ;
 wire \reg_module/_00409_ ;
 wire \reg_module/_00410_ ;
 wire \reg_module/_00411_ ;
 wire \reg_module/_00412_ ;
 wire \reg_module/_00413_ ;
 wire \reg_module/_00414_ ;
 wire \reg_module/_00415_ ;
 wire \reg_module/_00416_ ;
 wire \reg_module/_00417_ ;
 wire \reg_module/_00418_ ;
 wire \reg_module/_00419_ ;
 wire \reg_module/_00420_ ;
 wire \reg_module/_00421_ ;
 wire \reg_module/_00422_ ;
 wire \reg_module/_00423_ ;
 wire \reg_module/_00424_ ;
 wire \reg_module/_00425_ ;
 wire \reg_module/_00426_ ;
 wire \reg_module/_00427_ ;
 wire \reg_module/_00428_ ;
 wire \reg_module/_00429_ ;
 wire \reg_module/_00430_ ;
 wire \reg_module/_00431_ ;
 wire \reg_module/_00432_ ;
 wire \reg_module/_00433_ ;
 wire \reg_module/_00434_ ;
 wire \reg_module/_00435_ ;
 wire \reg_module/_00436_ ;
 wire \reg_module/_00437_ ;
 wire \reg_module/_00438_ ;
 wire \reg_module/_00439_ ;
 wire \reg_module/_00440_ ;
 wire \reg_module/_00441_ ;
 wire \reg_module/_00442_ ;
 wire \reg_module/_00443_ ;
 wire \reg_module/_00444_ ;
 wire \reg_module/_00445_ ;
 wire \reg_module/_00446_ ;
 wire \reg_module/_00447_ ;
 wire \reg_module/_00448_ ;
 wire \reg_module/_00449_ ;
 wire \reg_module/_00450_ ;
 wire \reg_module/_00451_ ;
 wire \reg_module/_00452_ ;
 wire \reg_module/_00453_ ;
 wire \reg_module/_00454_ ;
 wire \reg_module/_00455_ ;
 wire \reg_module/_00456_ ;
 wire \reg_module/_00457_ ;
 wire \reg_module/_00458_ ;
 wire \reg_module/_00459_ ;
 wire \reg_module/_00460_ ;
 wire \reg_module/_00461_ ;
 wire \reg_module/_00462_ ;
 wire \reg_module/_00463_ ;
 wire \reg_module/_00464_ ;
 wire \reg_module/_00465_ ;
 wire \reg_module/_00466_ ;
 wire \reg_module/_00467_ ;
 wire \reg_module/_00468_ ;
 wire \reg_module/_00469_ ;
 wire \reg_module/_00470_ ;
 wire \reg_module/_00471_ ;
 wire \reg_module/_00472_ ;
 wire \reg_module/_00473_ ;
 wire \reg_module/_00474_ ;
 wire \reg_module/_00475_ ;
 wire \reg_module/_00476_ ;
 wire \reg_module/_00477_ ;
 wire \reg_module/_00478_ ;
 wire \reg_module/_00479_ ;
 wire \reg_module/_00480_ ;
 wire \reg_module/_00481_ ;
 wire \reg_module/_00482_ ;
 wire \reg_module/_00483_ ;
 wire \reg_module/_00484_ ;
 wire \reg_module/_00485_ ;
 wire \reg_module/_00486_ ;
 wire \reg_module/_00487_ ;
 wire \reg_module/_00488_ ;
 wire \reg_module/_00489_ ;
 wire \reg_module/_00490_ ;
 wire \reg_module/_00491_ ;
 wire \reg_module/_00492_ ;
 wire \reg_module/_00493_ ;
 wire \reg_module/_00494_ ;
 wire \reg_module/_00495_ ;
 wire \reg_module/_00496_ ;
 wire \reg_module/_00497_ ;
 wire \reg_module/_00498_ ;
 wire \reg_module/_00499_ ;
 wire \reg_module/_00500_ ;
 wire \reg_module/_00501_ ;
 wire \reg_module/_00502_ ;
 wire \reg_module/_00503_ ;
 wire \reg_module/_00504_ ;
 wire \reg_module/_00505_ ;
 wire \reg_module/_00506_ ;
 wire \reg_module/_00507_ ;
 wire \reg_module/_00508_ ;
 wire \reg_module/_00509_ ;
 wire \reg_module/_00510_ ;
 wire \reg_module/_00511_ ;
 wire \reg_module/_00512_ ;
 wire \reg_module/_00513_ ;
 wire \reg_module/_00514_ ;
 wire \reg_module/_00515_ ;
 wire \reg_module/_00516_ ;
 wire \reg_module/_00517_ ;
 wire \reg_module/_00518_ ;
 wire \reg_module/_00519_ ;
 wire \reg_module/_00520_ ;
 wire \reg_module/_00521_ ;
 wire \reg_module/_00522_ ;
 wire \reg_module/_00523_ ;
 wire \reg_module/_00524_ ;
 wire \reg_module/_00525_ ;
 wire \reg_module/_00526_ ;
 wire \reg_module/_00527_ ;
 wire \reg_module/_00528_ ;
 wire \reg_module/_00529_ ;
 wire \reg_module/_00530_ ;
 wire \reg_module/_00531_ ;
 wire \reg_module/_00532_ ;
 wire \reg_module/_00533_ ;
 wire \reg_module/_00534_ ;
 wire \reg_module/_00535_ ;
 wire \reg_module/_00536_ ;
 wire \reg_module/_00537_ ;
 wire \reg_module/_00538_ ;
 wire \reg_module/_00539_ ;
 wire \reg_module/_00540_ ;
 wire \reg_module/_00541_ ;
 wire \reg_module/_00542_ ;
 wire \reg_module/_00543_ ;
 wire \reg_module/_00544_ ;
 wire \reg_module/_00545_ ;
 wire \reg_module/_00546_ ;
 wire \reg_module/_00547_ ;
 wire \reg_module/_00548_ ;
 wire \reg_module/_00549_ ;
 wire \reg_module/_00550_ ;
 wire \reg_module/_00551_ ;
 wire \reg_module/_00552_ ;
 wire \reg_module/_00553_ ;
 wire \reg_module/_00554_ ;
 wire \reg_module/_00555_ ;
 wire \reg_module/_00556_ ;
 wire \reg_module/_00557_ ;
 wire \reg_module/_00558_ ;
 wire \reg_module/_00559_ ;
 wire \reg_module/_00560_ ;
 wire \reg_module/_00561_ ;
 wire \reg_module/_00562_ ;
 wire \reg_module/_00563_ ;
 wire \reg_module/_00564_ ;
 wire \reg_module/_00565_ ;
 wire \reg_module/_00566_ ;
 wire \reg_module/_00567_ ;
 wire \reg_module/_00568_ ;
 wire \reg_module/_00569_ ;
 wire \reg_module/_00570_ ;
 wire \reg_module/_00571_ ;
 wire \reg_module/_00572_ ;
 wire \reg_module/_00573_ ;
 wire \reg_module/_00574_ ;
 wire \reg_module/_00575_ ;
 wire \reg_module/_00576_ ;
 wire \reg_module/_00577_ ;
 wire \reg_module/_00578_ ;
 wire \reg_module/_00579_ ;
 wire \reg_module/_00580_ ;
 wire \reg_module/_00581_ ;
 wire \reg_module/_00582_ ;
 wire \reg_module/_00583_ ;
 wire \reg_module/_00584_ ;
 wire \reg_module/_00585_ ;
 wire \reg_module/_00586_ ;
 wire \reg_module/_00587_ ;
 wire \reg_module/_00588_ ;
 wire \reg_module/_00589_ ;
 wire \reg_module/_00590_ ;
 wire \reg_module/_00591_ ;
 wire \reg_module/_00592_ ;
 wire \reg_module/_00593_ ;
 wire \reg_module/_00594_ ;
 wire \reg_module/_00595_ ;
 wire \reg_module/_00596_ ;
 wire \reg_module/_00597_ ;
 wire \reg_module/_00598_ ;
 wire \reg_module/_00599_ ;
 wire \reg_module/_00600_ ;
 wire \reg_module/_00601_ ;
 wire \reg_module/_00602_ ;
 wire \reg_module/_00603_ ;
 wire \reg_module/_00604_ ;
 wire \reg_module/_00605_ ;
 wire \reg_module/_00606_ ;
 wire \reg_module/_00607_ ;
 wire \reg_module/_00608_ ;
 wire \reg_module/_00609_ ;
 wire \reg_module/_00610_ ;
 wire \reg_module/_00611_ ;
 wire \reg_module/_00612_ ;
 wire \reg_module/_00613_ ;
 wire \reg_module/_00614_ ;
 wire \reg_module/_00615_ ;
 wire \reg_module/_00616_ ;
 wire \reg_module/_00617_ ;
 wire \reg_module/_00618_ ;
 wire \reg_module/_00619_ ;
 wire \reg_module/_00620_ ;
 wire \reg_module/_00621_ ;
 wire \reg_module/_00622_ ;
 wire \reg_module/_00623_ ;
 wire \reg_module/_00624_ ;
 wire \reg_module/_00625_ ;
 wire \reg_module/_00626_ ;
 wire \reg_module/_00627_ ;
 wire \reg_module/_00628_ ;
 wire \reg_module/_00629_ ;
 wire \reg_module/_00630_ ;
 wire \reg_module/_00631_ ;
 wire \reg_module/_00632_ ;
 wire \reg_module/_00633_ ;
 wire \reg_module/_00634_ ;
 wire \reg_module/_00635_ ;
 wire \reg_module/_00636_ ;
 wire \reg_module/_00637_ ;
 wire \reg_module/_00638_ ;
 wire \reg_module/_00639_ ;
 wire \reg_module/_00640_ ;
 wire \reg_module/_00641_ ;
 wire \reg_module/_00642_ ;
 wire \reg_module/_00643_ ;
 wire \reg_module/_00644_ ;
 wire \reg_module/_00645_ ;
 wire \reg_module/_00646_ ;
 wire \reg_module/_00647_ ;
 wire \reg_module/_00648_ ;
 wire \reg_module/_00649_ ;
 wire \reg_module/_00650_ ;
 wire \reg_module/_00651_ ;
 wire \reg_module/_00652_ ;
 wire \reg_module/_00653_ ;
 wire \reg_module/_00654_ ;
 wire \reg_module/_00655_ ;
 wire \reg_module/_00656_ ;
 wire \reg_module/_00657_ ;
 wire \reg_module/_00658_ ;
 wire \reg_module/_00659_ ;
 wire \reg_module/_00660_ ;
 wire \reg_module/_00661_ ;
 wire \reg_module/_00662_ ;
 wire \reg_module/_00663_ ;
 wire \reg_module/_00664_ ;
 wire \reg_module/_00665_ ;
 wire \reg_module/_00666_ ;
 wire \reg_module/_00667_ ;
 wire \reg_module/_00668_ ;
 wire \reg_module/_00669_ ;
 wire \reg_module/_00670_ ;
 wire \reg_module/_00671_ ;
 wire \reg_module/_00672_ ;
 wire \reg_module/_00673_ ;
 wire \reg_module/_00674_ ;
 wire \reg_module/_00675_ ;
 wire \reg_module/_00676_ ;
 wire \reg_module/_00677_ ;
 wire \reg_module/_00678_ ;
 wire \reg_module/_00679_ ;
 wire \reg_module/_00680_ ;
 wire \reg_module/_00681_ ;
 wire \reg_module/_00682_ ;
 wire \reg_module/_00683_ ;
 wire \reg_module/_00684_ ;
 wire \reg_module/_00685_ ;
 wire \reg_module/_00686_ ;
 wire \reg_module/_00687_ ;
 wire \reg_module/_00688_ ;
 wire \reg_module/_00689_ ;
 wire \reg_module/_00690_ ;
 wire \reg_module/_00691_ ;
 wire \reg_module/_00692_ ;
 wire \reg_module/_00693_ ;
 wire \reg_module/_00694_ ;
 wire \reg_module/_00695_ ;
 wire \reg_module/_00696_ ;
 wire \reg_module/_00697_ ;
 wire \reg_module/_00698_ ;
 wire \reg_module/_00699_ ;
 wire \reg_module/_00700_ ;
 wire \reg_module/_00701_ ;
 wire \reg_module/_00702_ ;
 wire \reg_module/_00703_ ;
 wire \reg_module/_00704_ ;
 wire \reg_module/_00705_ ;
 wire \reg_module/_00706_ ;
 wire \reg_module/_00707_ ;
 wire \reg_module/_00708_ ;
 wire \reg_module/_00709_ ;
 wire \reg_module/_00710_ ;
 wire \reg_module/_00711_ ;
 wire \reg_module/_00712_ ;
 wire \reg_module/_00713_ ;
 wire \reg_module/_00714_ ;
 wire \reg_module/_00715_ ;
 wire \reg_module/_00716_ ;
 wire \reg_module/_00717_ ;
 wire \reg_module/_00718_ ;
 wire \reg_module/_00719_ ;
 wire \reg_module/_00720_ ;
 wire \reg_module/_00721_ ;
 wire \reg_module/_00722_ ;
 wire \reg_module/_00723_ ;
 wire \reg_module/_00724_ ;
 wire \reg_module/_00725_ ;
 wire \reg_module/_00726_ ;
 wire \reg_module/_00727_ ;
 wire \reg_module/_00728_ ;
 wire \reg_module/_00729_ ;
 wire \reg_module/_00730_ ;
 wire \reg_module/_00731_ ;
 wire \reg_module/_00732_ ;
 wire \reg_module/_00733_ ;
 wire \reg_module/_00734_ ;
 wire \reg_module/_00735_ ;
 wire \reg_module/_00736_ ;
 wire \reg_module/_00737_ ;
 wire \reg_module/_00738_ ;
 wire \reg_module/_00739_ ;
 wire \reg_module/_00740_ ;
 wire \reg_module/_00741_ ;
 wire \reg_module/_00742_ ;
 wire \reg_module/_00743_ ;
 wire \reg_module/_00744_ ;
 wire \reg_module/_00745_ ;
 wire \reg_module/_00746_ ;
 wire \reg_module/_00747_ ;
 wire \reg_module/_00748_ ;
 wire \reg_module/_00749_ ;
 wire \reg_module/_00750_ ;
 wire \reg_module/_00751_ ;
 wire \reg_module/_00752_ ;
 wire \reg_module/_00753_ ;
 wire \reg_module/_00754_ ;
 wire \reg_module/_00755_ ;
 wire \reg_module/_00756_ ;
 wire \reg_module/_00757_ ;
 wire \reg_module/_00758_ ;
 wire \reg_module/_00759_ ;
 wire \reg_module/_00760_ ;
 wire \reg_module/_00761_ ;
 wire \reg_module/_00762_ ;
 wire \reg_module/_00763_ ;
 wire \reg_module/_00764_ ;
 wire \reg_module/_00765_ ;
 wire \reg_module/_00766_ ;
 wire \reg_module/_00767_ ;
 wire \reg_module/_00768_ ;
 wire \reg_module/_00769_ ;
 wire \reg_module/_00770_ ;
 wire \reg_module/_00771_ ;
 wire \reg_module/_00772_ ;
 wire \reg_module/_00773_ ;
 wire \reg_module/_00774_ ;
 wire \reg_module/_00775_ ;
 wire \reg_module/_00776_ ;
 wire \reg_module/_00777_ ;
 wire \reg_module/_00778_ ;
 wire \reg_module/_00779_ ;
 wire \reg_module/_00780_ ;
 wire \reg_module/_00781_ ;
 wire \reg_module/_00782_ ;
 wire \reg_module/_00783_ ;
 wire \reg_module/_00784_ ;
 wire \reg_module/_00785_ ;
 wire \reg_module/_00786_ ;
 wire \reg_module/_00787_ ;
 wire \reg_module/_00788_ ;
 wire \reg_module/_00789_ ;
 wire \reg_module/_00790_ ;
 wire \reg_module/_00791_ ;
 wire \reg_module/_00792_ ;
 wire \reg_module/_00793_ ;
 wire \reg_module/_00794_ ;
 wire \reg_module/_00795_ ;
 wire \reg_module/_00796_ ;
 wire \reg_module/_00797_ ;
 wire \reg_module/_00798_ ;
 wire \reg_module/_00799_ ;
 wire \reg_module/_00800_ ;
 wire \reg_module/_00801_ ;
 wire \reg_module/_00802_ ;
 wire \reg_module/_00803_ ;
 wire \reg_module/_00804_ ;
 wire \reg_module/_00805_ ;
 wire \reg_module/_00806_ ;
 wire \reg_module/_00807_ ;
 wire \reg_module/_00808_ ;
 wire \reg_module/_00809_ ;
 wire \reg_module/_00810_ ;
 wire \reg_module/_00811_ ;
 wire \reg_module/_00812_ ;
 wire \reg_module/_00813_ ;
 wire \reg_module/_00814_ ;
 wire \reg_module/_00815_ ;
 wire \reg_module/_00816_ ;
 wire \reg_module/_00817_ ;
 wire \reg_module/_00818_ ;
 wire \reg_module/_00819_ ;
 wire \reg_module/_00820_ ;
 wire \reg_module/_00821_ ;
 wire \reg_module/_00822_ ;
 wire \reg_module/_00823_ ;
 wire \reg_module/_00824_ ;
 wire \reg_module/_00825_ ;
 wire \reg_module/_00826_ ;
 wire \reg_module/_00827_ ;
 wire \reg_module/_00828_ ;
 wire \reg_module/_00829_ ;
 wire \reg_module/_00830_ ;
 wire \reg_module/_00831_ ;
 wire \reg_module/_00832_ ;
 wire \reg_module/_00833_ ;
 wire \reg_module/_00834_ ;
 wire \reg_module/_00835_ ;
 wire \reg_module/_00836_ ;
 wire \reg_module/_00837_ ;
 wire \reg_module/_00838_ ;
 wire \reg_module/_00839_ ;
 wire \reg_module/_00840_ ;
 wire \reg_module/_00841_ ;
 wire \reg_module/_00842_ ;
 wire \reg_module/_00843_ ;
 wire \reg_module/_00844_ ;
 wire \reg_module/_00845_ ;
 wire \reg_module/_00846_ ;
 wire \reg_module/_00847_ ;
 wire \reg_module/_00848_ ;
 wire \reg_module/_00849_ ;
 wire \reg_module/_00850_ ;
 wire \reg_module/_00851_ ;
 wire \reg_module/_00852_ ;
 wire \reg_module/_00853_ ;
 wire \reg_module/_00854_ ;
 wire \reg_module/_00855_ ;
 wire \reg_module/_00856_ ;
 wire \reg_module/_00857_ ;
 wire \reg_module/_00858_ ;
 wire \reg_module/_00859_ ;
 wire \reg_module/_00860_ ;
 wire \reg_module/_00861_ ;
 wire \reg_module/_00862_ ;
 wire \reg_module/_00863_ ;
 wire \reg_module/_00864_ ;
 wire \reg_module/_00865_ ;
 wire \reg_module/_00866_ ;
 wire \reg_module/_00867_ ;
 wire \reg_module/_00868_ ;
 wire \reg_module/_00869_ ;
 wire \reg_module/_00870_ ;
 wire \reg_module/_00871_ ;
 wire \reg_module/_00872_ ;
 wire \reg_module/_00873_ ;
 wire \reg_module/_00874_ ;
 wire \reg_module/_00875_ ;
 wire \reg_module/_00876_ ;
 wire \reg_module/_00877_ ;
 wire \reg_module/_00878_ ;
 wire \reg_module/_00879_ ;
 wire \reg_module/_00880_ ;
 wire \reg_module/_00881_ ;
 wire \reg_module/_00882_ ;
 wire \reg_module/_00883_ ;
 wire \reg_module/_00884_ ;
 wire \reg_module/_00885_ ;
 wire \reg_module/_00886_ ;
 wire \reg_module/_00887_ ;
 wire \reg_module/_00888_ ;
 wire \reg_module/_00889_ ;
 wire \reg_module/_00890_ ;
 wire \reg_module/_00891_ ;
 wire \reg_module/_00892_ ;
 wire \reg_module/_00893_ ;
 wire \reg_module/_00894_ ;
 wire \reg_module/_00895_ ;
 wire \reg_module/_00896_ ;
 wire \reg_module/_00897_ ;
 wire \reg_module/_00898_ ;
 wire \reg_module/_00899_ ;
 wire \reg_module/_00900_ ;
 wire \reg_module/_00901_ ;
 wire \reg_module/_00902_ ;
 wire \reg_module/_00903_ ;
 wire \reg_module/_00904_ ;
 wire \reg_module/_00905_ ;
 wire \reg_module/_00906_ ;
 wire \reg_module/_00907_ ;
 wire \reg_module/_00908_ ;
 wire \reg_module/_00909_ ;
 wire \reg_module/_00910_ ;
 wire \reg_module/_00911_ ;
 wire \reg_module/_00912_ ;
 wire \reg_module/_00913_ ;
 wire \reg_module/_00914_ ;
 wire \reg_module/_00915_ ;
 wire \reg_module/_00916_ ;
 wire \reg_module/_00917_ ;
 wire \reg_module/_00918_ ;
 wire \reg_module/_00919_ ;
 wire \reg_module/_00920_ ;
 wire \reg_module/_00921_ ;
 wire \reg_module/_00922_ ;
 wire \reg_module/_00923_ ;
 wire \reg_module/_00924_ ;
 wire \reg_module/_00925_ ;
 wire \reg_module/_00926_ ;
 wire \reg_module/_00927_ ;
 wire \reg_module/_00928_ ;
 wire \reg_module/_00929_ ;
 wire \reg_module/_00930_ ;
 wire \reg_module/_00931_ ;
 wire \reg_module/_00932_ ;
 wire \reg_module/_00933_ ;
 wire \reg_module/_00934_ ;
 wire \reg_module/_00935_ ;
 wire \reg_module/_00936_ ;
 wire \reg_module/_00937_ ;
 wire \reg_module/_00938_ ;
 wire \reg_module/_00939_ ;
 wire \reg_module/_00940_ ;
 wire \reg_module/_00941_ ;
 wire \reg_module/_00942_ ;
 wire \reg_module/_00943_ ;
 wire \reg_module/_00944_ ;
 wire \reg_module/_00945_ ;
 wire \reg_module/_00946_ ;
 wire \reg_module/_00947_ ;
 wire \reg_module/_00948_ ;
 wire \reg_module/_00949_ ;
 wire \reg_module/_00950_ ;
 wire \reg_module/_00951_ ;
 wire \reg_module/_00952_ ;
 wire \reg_module/_00953_ ;
 wire \reg_module/_00954_ ;
 wire \reg_module/_00955_ ;
 wire \reg_module/_00956_ ;
 wire \reg_module/_00957_ ;
 wire \reg_module/_00958_ ;
 wire \reg_module/_00959_ ;
 wire \reg_module/_00960_ ;
 wire \reg_module/_00961_ ;
 wire \reg_module/_00962_ ;
 wire \reg_module/_00963_ ;
 wire \reg_module/_00964_ ;
 wire \reg_module/_00965_ ;
 wire \reg_module/_00966_ ;
 wire \reg_module/_00967_ ;
 wire \reg_module/_00968_ ;
 wire \reg_module/_00969_ ;
 wire \reg_module/_00970_ ;
 wire \reg_module/_00971_ ;
 wire \reg_module/_00972_ ;
 wire \reg_module/_00973_ ;
 wire \reg_module/_00974_ ;
 wire \reg_module/_00975_ ;
 wire \reg_module/_00976_ ;
 wire \reg_module/_00977_ ;
 wire \reg_module/_00978_ ;
 wire \reg_module/_00979_ ;
 wire \reg_module/_00980_ ;
 wire \reg_module/_00981_ ;
 wire \reg_module/_00982_ ;
 wire \reg_module/_00983_ ;
 wire \reg_module/_00984_ ;
 wire \reg_module/_00985_ ;
 wire \reg_module/_00986_ ;
 wire \reg_module/_00987_ ;
 wire \reg_module/_00988_ ;
 wire \reg_module/_00989_ ;
 wire \reg_module/_00990_ ;
 wire \reg_module/_00991_ ;
 wire \reg_module/_00992_ ;
 wire \reg_module/_00993_ ;
 wire \reg_module/_00994_ ;
 wire \reg_module/_00995_ ;
 wire \reg_module/_00996_ ;
 wire \reg_module/_00997_ ;
 wire \reg_module/_00998_ ;
 wire \reg_module/_00999_ ;
 wire \reg_module/_01000_ ;
 wire \reg_module/_01001_ ;
 wire \reg_module/_01002_ ;
 wire \reg_module/_01003_ ;
 wire \reg_module/_01004_ ;
 wire \reg_module/_01005_ ;
 wire \reg_module/_01006_ ;
 wire \reg_module/_01007_ ;
 wire \reg_module/_01008_ ;
 wire \reg_module/_01009_ ;
 wire \reg_module/_01010_ ;
 wire \reg_module/_01011_ ;
 wire \reg_module/_01012_ ;
 wire \reg_module/_01013_ ;
 wire \reg_module/_01014_ ;
 wire \reg_module/_01015_ ;
 wire \reg_module/_01016_ ;
 wire \reg_module/_01017_ ;
 wire \reg_module/_01018_ ;
 wire \reg_module/_01019_ ;
 wire \reg_module/_01020_ ;
 wire \reg_module/_01021_ ;
 wire \reg_module/_01022_ ;
 wire \reg_module/_01023_ ;
 wire \reg_module/_01024_ ;
 wire \reg_module/_01025_ ;
 wire \reg_module/_01026_ ;
 wire \reg_module/_01027_ ;
 wire \reg_module/_01028_ ;
 wire \reg_module/_01029_ ;
 wire \reg_module/_01030_ ;
 wire \reg_module/_01031_ ;
 wire \reg_module/_01032_ ;
 wire \reg_module/_01033_ ;
 wire \reg_module/_01034_ ;
 wire \reg_module/_01035_ ;
 wire \reg_module/_01036_ ;
 wire \reg_module/_01037_ ;
 wire \reg_module/_01038_ ;
 wire \reg_module/_01039_ ;
 wire \reg_module/_01040_ ;
 wire \reg_module/_01041_ ;
 wire \reg_module/_01042_ ;
 wire \reg_module/_01043_ ;
 wire \reg_module/_01044_ ;
 wire \reg_module/_01045_ ;
 wire \reg_module/_01046_ ;
 wire \reg_module/_01047_ ;
 wire \reg_module/_01048_ ;
 wire \reg_module/_01049_ ;
 wire \reg_module/_01050_ ;
 wire \reg_module/_01051_ ;
 wire \reg_module/_01052_ ;
 wire \reg_module/_01053_ ;
 wire \reg_module/_01054_ ;
 wire \reg_module/_01055_ ;
 wire \reg_module/_01056_ ;
 wire \reg_module/_01057_ ;
 wire \reg_module/_01058_ ;
 wire \reg_module/_01059_ ;
 wire \reg_module/_01060_ ;
 wire \reg_module/_01061_ ;
 wire \reg_module/_01062_ ;
 wire \reg_module/_01063_ ;
 wire \reg_module/_01064_ ;
 wire \reg_module/_01065_ ;
 wire \reg_module/_01066_ ;
 wire \reg_module/_01067_ ;
 wire \reg_module/_01068_ ;
 wire \reg_module/_01069_ ;
 wire \reg_module/_01070_ ;
 wire \reg_module/_01071_ ;
 wire \reg_module/_01072_ ;
 wire \reg_module/_01073_ ;
 wire \reg_module/_01074_ ;
 wire \reg_module/_01075_ ;
 wire \reg_module/_01076_ ;
 wire \reg_module/_01077_ ;
 wire \reg_module/_01078_ ;
 wire \reg_module/_01079_ ;
 wire \reg_module/_01080_ ;
 wire \reg_module/_01081_ ;
 wire \reg_module/_01082_ ;
 wire \reg_module/_01083_ ;
 wire \reg_module/_01084_ ;
 wire \reg_module/_01085_ ;
 wire \reg_module/_01086_ ;
 wire \reg_module/_01087_ ;
 wire \reg_module/_01088_ ;
 wire \reg_module/_01089_ ;
 wire \reg_module/_01090_ ;
 wire \reg_module/_01091_ ;
 wire \reg_module/_01092_ ;
 wire \reg_module/_01093_ ;
 wire \reg_module/_01094_ ;
 wire \reg_module/_01095_ ;
 wire \reg_module/_01096_ ;
 wire \reg_module/_01097_ ;
 wire \reg_module/_01098_ ;
 wire \reg_module/_01099_ ;
 wire \reg_module/_01100_ ;
 wire \reg_module/_01101_ ;
 wire \reg_module/_01102_ ;
 wire \reg_module/_01103_ ;
 wire \reg_module/_01104_ ;
 wire \reg_module/_01105_ ;
 wire \reg_module/_01106_ ;
 wire \reg_module/_01107_ ;
 wire \reg_module/_01108_ ;
 wire \reg_module/_01109_ ;
 wire \reg_module/_01110_ ;
 wire \reg_module/_01111_ ;
 wire \reg_module/_01112_ ;
 wire \reg_module/_01113_ ;
 wire \reg_module/_01114_ ;
 wire \reg_module/_01115_ ;
 wire \reg_module/_01116_ ;
 wire \reg_module/_01117_ ;
 wire \reg_module/_01118_ ;
 wire \reg_module/_01119_ ;
 wire \reg_module/_01120_ ;
 wire \reg_module/_01121_ ;
 wire \reg_module/_01122_ ;
 wire \reg_module/_01123_ ;
 wire \reg_module/_01124_ ;
 wire \reg_module/_01125_ ;
 wire \reg_module/_01126_ ;
 wire \reg_module/_01127_ ;
 wire \reg_module/_01128_ ;
 wire \reg_module/_01129_ ;
 wire \reg_module/_01130_ ;
 wire \reg_module/_01131_ ;
 wire \reg_module/_01132_ ;
 wire \reg_module/_01133_ ;
 wire \reg_module/_01134_ ;
 wire \reg_module/_01135_ ;
 wire \reg_module/_01136_ ;
 wire \reg_module/_01137_ ;
 wire \reg_module/_01138_ ;
 wire \reg_module/_01139_ ;
 wire \reg_module/_01140_ ;
 wire \reg_module/_01141_ ;
 wire \reg_module/_01142_ ;
 wire \reg_module/_01143_ ;
 wire \reg_module/_01144_ ;
 wire \reg_module/_01145_ ;
 wire \reg_module/_01146_ ;
 wire \reg_module/_01147_ ;
 wire \reg_module/_01148_ ;
 wire \reg_module/_01149_ ;
 wire \reg_module/_01150_ ;
 wire \reg_module/_01151_ ;
 wire \reg_module/_01152_ ;
 wire \reg_module/_01153_ ;
 wire \reg_module/_01154_ ;
 wire \reg_module/_01155_ ;
 wire \reg_module/_01156_ ;
 wire \reg_module/_01157_ ;
 wire \reg_module/_01158_ ;
 wire \reg_module/_01159_ ;
 wire \reg_module/_01160_ ;
 wire \reg_module/_01161_ ;
 wire \reg_module/_01162_ ;
 wire \reg_module/_01163_ ;
 wire \reg_module/_01164_ ;
 wire \reg_module/_01165_ ;
 wire \reg_module/_01166_ ;
 wire \reg_module/_01167_ ;
 wire \reg_module/_01168_ ;
 wire \reg_module/_01169_ ;
 wire \reg_module/_01170_ ;
 wire \reg_module/_01171_ ;
 wire \reg_module/_01172_ ;
 wire \reg_module/_01173_ ;
 wire \reg_module/_01174_ ;
 wire \reg_module/_01175_ ;
 wire \reg_module/_01176_ ;
 wire \reg_module/_01177_ ;
 wire \reg_module/_01178_ ;
 wire \reg_module/_01179_ ;
 wire \reg_module/_01180_ ;
 wire \reg_module/_01181_ ;
 wire \reg_module/_01182_ ;
 wire \reg_module/_01183_ ;
 wire \reg_module/_01184_ ;
 wire \reg_module/_01185_ ;
 wire \reg_module/_01186_ ;
 wire \reg_module/_01187_ ;
 wire \reg_module/_01188_ ;
 wire \reg_module/_01189_ ;
 wire \reg_module/_01190_ ;
 wire \reg_module/_01191_ ;
 wire \reg_module/_01192_ ;
 wire \reg_module/_01193_ ;
 wire \reg_module/_01194_ ;
 wire \reg_module/_01195_ ;
 wire \reg_module/_01196_ ;
 wire \reg_module/_01197_ ;
 wire \reg_module/_01198_ ;
 wire \reg_module/_01199_ ;
 wire \reg_module/_01200_ ;
 wire \reg_module/_01201_ ;
 wire \reg_module/_01202_ ;
 wire \reg_module/_01203_ ;
 wire \reg_module/_01204_ ;
 wire \reg_module/_01205_ ;
 wire \reg_module/_01206_ ;
 wire \reg_module/_01207_ ;
 wire \reg_module/_01208_ ;
 wire \reg_module/_01209_ ;
 wire \reg_module/_01210_ ;
 wire \reg_module/_01211_ ;
 wire \reg_module/_01212_ ;
 wire \reg_module/_01213_ ;
 wire \reg_module/_01214_ ;
 wire \reg_module/_01215_ ;
 wire \reg_module/_01216_ ;
 wire \reg_module/_01217_ ;
 wire \reg_module/_01218_ ;
 wire \reg_module/_01219_ ;
 wire \reg_module/_01220_ ;
 wire \reg_module/_01221_ ;
 wire \reg_module/_01222_ ;
 wire \reg_module/_01223_ ;
 wire \reg_module/_01224_ ;
 wire \reg_module/_01225_ ;
 wire \reg_module/_01226_ ;
 wire \reg_module/_01227_ ;
 wire \reg_module/_01228_ ;
 wire \reg_module/_01229_ ;
 wire \reg_module/_01230_ ;
 wire \reg_module/_01231_ ;
 wire \reg_module/_01232_ ;
 wire \reg_module/_01233_ ;
 wire \reg_module/_01234_ ;
 wire \reg_module/_01235_ ;
 wire \reg_module/_01236_ ;
 wire \reg_module/_01237_ ;
 wire \reg_module/_01238_ ;
 wire \reg_module/_01239_ ;
 wire \reg_module/_01240_ ;
 wire \reg_module/_01241_ ;
 wire \reg_module/_01242_ ;
 wire \reg_module/_01243_ ;
 wire \reg_module/_01244_ ;
 wire \reg_module/_01245_ ;
 wire \reg_module/_01246_ ;
 wire \reg_module/_01247_ ;
 wire \reg_module/_01248_ ;
 wire \reg_module/_01249_ ;
 wire \reg_module/_01250_ ;
 wire \reg_module/_01251_ ;
 wire \reg_module/_01252_ ;
 wire \reg_module/_01253_ ;
 wire \reg_module/_01254_ ;
 wire \reg_module/_01255_ ;
 wire \reg_module/_01256_ ;
 wire \reg_module/_01257_ ;
 wire \reg_module/_01258_ ;
 wire \reg_module/_01259_ ;
 wire \reg_module/_01260_ ;
 wire \reg_module/_01261_ ;
 wire \reg_module/_01262_ ;
 wire \reg_module/_01263_ ;
 wire \reg_module/_01264_ ;
 wire \reg_module/_01265_ ;
 wire \reg_module/_01266_ ;
 wire \reg_module/_01267_ ;
 wire \reg_module/_01268_ ;
 wire \reg_module/_01269_ ;
 wire \reg_module/_01270_ ;
 wire \reg_module/_01271_ ;
 wire \reg_module/_01272_ ;
 wire \reg_module/_01273_ ;
 wire \reg_module/_01274_ ;
 wire \reg_module/_01275_ ;
 wire \reg_module/_01276_ ;
 wire \reg_module/_01277_ ;
 wire \reg_module/_01278_ ;
 wire \reg_module/_01279_ ;
 wire \reg_module/_01280_ ;
 wire \reg_module/_01281_ ;
 wire \reg_module/_01282_ ;
 wire \reg_module/_01283_ ;
 wire \reg_module/_01284_ ;
 wire \reg_module/_01285_ ;
 wire \reg_module/_01286_ ;
 wire \reg_module/_01287_ ;
 wire \reg_module/_01288_ ;
 wire \reg_module/_01289_ ;
 wire \reg_module/_01290_ ;
 wire \reg_module/_01291_ ;
 wire \reg_module/_01292_ ;
 wire \reg_module/_01293_ ;
 wire \reg_module/_01294_ ;
 wire \reg_module/_01295_ ;
 wire \reg_module/_01296_ ;
 wire \reg_module/_01297_ ;
 wire \reg_module/_01298_ ;
 wire \reg_module/_01299_ ;
 wire \reg_module/_01300_ ;
 wire \reg_module/_01301_ ;
 wire \reg_module/_01302_ ;
 wire \reg_module/_01303_ ;
 wire \reg_module/_01304_ ;
 wire \reg_module/_01305_ ;
 wire \reg_module/_01306_ ;
 wire \reg_module/_01307_ ;
 wire \reg_module/_01308_ ;
 wire \reg_module/_01309_ ;
 wire \reg_module/_01310_ ;
 wire \reg_module/_01311_ ;
 wire \reg_module/_01312_ ;
 wire \reg_module/_01313_ ;
 wire \reg_module/_01314_ ;
 wire \reg_module/_01315_ ;
 wire \reg_module/_01316_ ;
 wire \reg_module/_01317_ ;
 wire \reg_module/_01318_ ;
 wire \reg_module/_01319_ ;
 wire \reg_module/_01320_ ;
 wire \reg_module/_01321_ ;
 wire \reg_module/_01322_ ;
 wire \reg_module/_01323_ ;
 wire \reg_module/_01324_ ;
 wire \reg_module/_01325_ ;
 wire \reg_module/_01326_ ;
 wire \reg_module/_01327_ ;
 wire \reg_module/_01328_ ;
 wire \reg_module/_01329_ ;
 wire \reg_module/_01330_ ;
 wire \reg_module/_01331_ ;
 wire \reg_module/_01332_ ;
 wire \reg_module/_01333_ ;
 wire \reg_module/_01334_ ;
 wire \reg_module/_01335_ ;
 wire \reg_module/_01336_ ;
 wire \reg_module/_01337_ ;
 wire \reg_module/_01338_ ;
 wire \reg_module/_01339_ ;
 wire \reg_module/_01340_ ;
 wire \reg_module/_01341_ ;
 wire \reg_module/_01342_ ;
 wire \reg_module/_01343_ ;
 wire \reg_module/_01344_ ;
 wire \reg_module/_01345_ ;
 wire \reg_module/_01346_ ;
 wire \reg_module/_01347_ ;
 wire \reg_module/_01348_ ;
 wire \reg_module/_01349_ ;
 wire \reg_module/_01350_ ;
 wire \reg_module/_01351_ ;
 wire \reg_module/_01352_ ;
 wire \reg_module/_01353_ ;
 wire \reg_module/_01354_ ;
 wire \reg_module/_01355_ ;
 wire \reg_module/_01356_ ;
 wire \reg_module/_01357_ ;
 wire \reg_module/_01358_ ;
 wire \reg_module/_01359_ ;
 wire \reg_module/_01360_ ;
 wire \reg_module/_01361_ ;
 wire \reg_module/_01362_ ;
 wire \reg_module/_01363_ ;
 wire \reg_module/_01364_ ;
 wire \reg_module/_01365_ ;
 wire \reg_module/_01366_ ;
 wire \reg_module/_01367_ ;
 wire \reg_module/_01368_ ;
 wire \reg_module/_01369_ ;
 wire \reg_module/_01370_ ;
 wire \reg_module/_01371_ ;
 wire \reg_module/_01372_ ;
 wire \reg_module/_01373_ ;
 wire \reg_module/_01374_ ;
 wire \reg_module/_01375_ ;
 wire \reg_module/_01376_ ;
 wire \reg_module/_01377_ ;
 wire \reg_module/_01378_ ;
 wire \reg_module/_01379_ ;
 wire \reg_module/_01380_ ;
 wire \reg_module/_01381_ ;
 wire \reg_module/_01382_ ;
 wire \reg_module/_01383_ ;
 wire \reg_module/_01384_ ;
 wire \reg_module/_01385_ ;
 wire \reg_module/_01386_ ;
 wire \reg_module/_01387_ ;
 wire \reg_module/_01388_ ;
 wire \reg_module/_01389_ ;
 wire \reg_module/_01390_ ;
 wire \reg_module/_01391_ ;
 wire \reg_module/_01392_ ;
 wire \reg_module/_01393_ ;
 wire \reg_module/_01394_ ;
 wire \reg_module/_01395_ ;
 wire \reg_module/_01396_ ;
 wire \reg_module/_01397_ ;
 wire \reg_module/_01398_ ;
 wire \reg_module/_01399_ ;
 wire \reg_module/_01400_ ;
 wire \reg_module/_01401_ ;
 wire \reg_module/_01402_ ;
 wire \reg_module/_01403_ ;
 wire \reg_module/_01404_ ;
 wire \reg_module/_01405_ ;
 wire \reg_module/_01406_ ;
 wire \reg_module/_01407_ ;
 wire \reg_module/_01408_ ;
 wire \reg_module/_01409_ ;
 wire \reg_module/_01410_ ;
 wire \reg_module/_01411_ ;
 wire \reg_module/_01412_ ;
 wire \reg_module/_01413_ ;
 wire \reg_module/_01414_ ;
 wire \reg_module/_01415_ ;
 wire \reg_module/_01416_ ;
 wire \reg_module/_01417_ ;
 wire \reg_module/_01418_ ;
 wire \reg_module/_01419_ ;
 wire \reg_module/_01420_ ;
 wire \reg_module/_01421_ ;
 wire \reg_module/_01422_ ;
 wire \reg_module/_01423_ ;
 wire \reg_module/_01424_ ;
 wire \reg_module/_01425_ ;
 wire \reg_module/_01426_ ;
 wire \reg_module/_01427_ ;
 wire \reg_module/_01428_ ;
 wire \reg_module/_01429_ ;
 wire \reg_module/_01430_ ;
 wire \reg_module/_01431_ ;
 wire \reg_module/_01432_ ;
 wire \reg_module/_01433_ ;
 wire \reg_module/_01434_ ;
 wire \reg_module/_01435_ ;
 wire \reg_module/_01436_ ;
 wire \reg_module/_01437_ ;
 wire \reg_module/_01438_ ;
 wire \reg_module/_01439_ ;
 wire \reg_module/_01440_ ;
 wire \reg_module/_01441_ ;
 wire \reg_module/_01442_ ;
 wire \reg_module/_01443_ ;
 wire \reg_module/_01444_ ;
 wire \reg_module/_01445_ ;
 wire \reg_module/_01446_ ;
 wire \reg_module/_01447_ ;
 wire \reg_module/_01448_ ;
 wire \reg_module/_01449_ ;
 wire \reg_module/_01450_ ;
 wire \reg_module/_01451_ ;
 wire \reg_module/_01452_ ;
 wire \reg_module/_01453_ ;
 wire \reg_module/_01454_ ;
 wire \reg_module/_01455_ ;
 wire \reg_module/_01456_ ;
 wire \reg_module/_01457_ ;
 wire \reg_module/_01458_ ;
 wire \reg_module/_01459_ ;
 wire \reg_module/_01460_ ;
 wire \reg_module/_01461_ ;
 wire \reg_module/_01462_ ;
 wire \reg_module/_01463_ ;
 wire \reg_module/_01464_ ;
 wire \reg_module/_01465_ ;
 wire \reg_module/_01466_ ;
 wire \reg_module/_01467_ ;
 wire \reg_module/_01468_ ;
 wire \reg_module/_01469_ ;
 wire \reg_module/_01470_ ;
 wire \reg_module/_01471_ ;
 wire \reg_module/_01472_ ;
 wire \reg_module/_01473_ ;
 wire \reg_module/_01474_ ;
 wire \reg_module/_01475_ ;
 wire \reg_module/_01476_ ;
 wire \reg_module/_01477_ ;
 wire \reg_module/_01478_ ;
 wire \reg_module/_01479_ ;
 wire \reg_module/_01480_ ;
 wire \reg_module/_01481_ ;
 wire \reg_module/_01482_ ;
 wire \reg_module/_01483_ ;
 wire \reg_module/_01484_ ;
 wire \reg_module/_01485_ ;
 wire \reg_module/_01486_ ;
 wire \reg_module/_01487_ ;
 wire \reg_module/_01488_ ;
 wire \reg_module/_01489_ ;
 wire \reg_module/_01490_ ;
 wire \reg_module/_01491_ ;
 wire \reg_module/_01492_ ;
 wire \reg_module/_01493_ ;
 wire \reg_module/_01494_ ;
 wire \reg_module/_01495_ ;
 wire \reg_module/_01496_ ;
 wire \reg_module/_01497_ ;
 wire \reg_module/_01498_ ;
 wire \reg_module/_01499_ ;
 wire \reg_module/_01500_ ;
 wire \reg_module/_01501_ ;
 wire \reg_module/_01502_ ;
 wire \reg_module/_01503_ ;
 wire \reg_module/_01504_ ;
 wire \reg_module/_01505_ ;
 wire \reg_module/_01506_ ;
 wire \reg_module/_01507_ ;
 wire \reg_module/_01508_ ;
 wire \reg_module/_01509_ ;
 wire \reg_module/_01510_ ;
 wire \reg_module/_01511_ ;
 wire \reg_module/_01512_ ;
 wire \reg_module/_01513_ ;
 wire \reg_module/_01514_ ;
 wire \reg_module/_01515_ ;
 wire \reg_module/_01516_ ;
 wire \reg_module/_01517_ ;
 wire \reg_module/_01518_ ;
 wire \reg_module/_01519_ ;
 wire \reg_module/_01520_ ;
 wire \reg_module/_01521_ ;
 wire \reg_module/_01522_ ;
 wire \reg_module/_01523_ ;
 wire \reg_module/_01524_ ;
 wire \reg_module/_01525_ ;
 wire \reg_module/_01526_ ;
 wire \reg_module/_01527_ ;
 wire \reg_module/_01528_ ;
 wire \reg_module/_01529_ ;
 wire \reg_module/_01530_ ;
 wire \reg_module/_01531_ ;
 wire \reg_module/_01532_ ;
 wire \reg_module/_01533_ ;
 wire \reg_module/_01534_ ;
 wire \reg_module/_01535_ ;
 wire \reg_module/_01536_ ;
 wire \reg_module/_01537_ ;
 wire \reg_module/_01538_ ;
 wire \reg_module/_01539_ ;
 wire \reg_module/_01540_ ;
 wire \reg_module/_01541_ ;
 wire \reg_module/_01542_ ;
 wire \reg_module/_01543_ ;
 wire \reg_module/_01544_ ;
 wire \reg_module/_01545_ ;
 wire \reg_module/_01546_ ;
 wire \reg_module/_01547_ ;
 wire \reg_module/_01548_ ;
 wire \reg_module/_01549_ ;
 wire \reg_module/_01550_ ;
 wire \reg_module/_01551_ ;
 wire \reg_module/_01552_ ;
 wire \reg_module/_01553_ ;
 wire \reg_module/_01554_ ;
 wire \reg_module/_01555_ ;
 wire \reg_module/_01556_ ;
 wire \reg_module/_01557_ ;
 wire \reg_module/_01558_ ;
 wire \reg_module/_01559_ ;
 wire \reg_module/_01560_ ;
 wire \reg_module/_01561_ ;
 wire \reg_module/_01562_ ;
 wire \reg_module/_01563_ ;
 wire \reg_module/_01564_ ;
 wire \reg_module/_01565_ ;
 wire \reg_module/_01566_ ;
 wire \reg_module/_01567_ ;
 wire \reg_module/_01568_ ;
 wire \reg_module/_01569_ ;
 wire \reg_module/_01570_ ;
 wire \reg_module/_01571_ ;
 wire \reg_module/_01572_ ;
 wire \reg_module/_01573_ ;
 wire \reg_module/_01574_ ;
 wire \reg_module/_01575_ ;
 wire \reg_module/_01576_ ;
 wire \reg_module/_01577_ ;
 wire \reg_module/_01578_ ;
 wire \reg_module/_01579_ ;
 wire \reg_module/_01580_ ;
 wire \reg_module/_01581_ ;
 wire \reg_module/_01582_ ;
 wire \reg_module/_01583_ ;
 wire \reg_module/_01584_ ;
 wire \reg_module/_01585_ ;
 wire \reg_module/_01586_ ;
 wire \reg_module/_01587_ ;
 wire \reg_module/_01588_ ;
 wire \reg_module/_01589_ ;
 wire \reg_module/_01590_ ;
 wire \reg_module/_01591_ ;
 wire \reg_module/_01592_ ;
 wire \reg_module/_01593_ ;
 wire \reg_module/_01594_ ;
 wire \reg_module/_01595_ ;
 wire \reg_module/_01596_ ;
 wire \reg_module/_01597_ ;
 wire \reg_module/_01598_ ;
 wire \reg_module/_01599_ ;
 wire \reg_module/_01600_ ;
 wire \reg_module/_01601_ ;
 wire \reg_module/_01602_ ;
 wire \reg_module/_01603_ ;
 wire \reg_module/_01604_ ;
 wire \reg_module/_01605_ ;
 wire \reg_module/_01606_ ;
 wire \reg_module/_01607_ ;
 wire \reg_module/_01608_ ;
 wire \reg_module/_01609_ ;
 wire \reg_module/_01610_ ;
 wire \reg_module/_01611_ ;
 wire \reg_module/_01612_ ;
 wire \reg_module/_01613_ ;
 wire \reg_module/_01614_ ;
 wire \reg_module/_01615_ ;
 wire \reg_module/_01616_ ;
 wire \reg_module/_01617_ ;
 wire \reg_module/_01618_ ;
 wire \reg_module/_01619_ ;
 wire \reg_module/_01620_ ;
 wire \reg_module/_01621_ ;
 wire \reg_module/_01622_ ;
 wire \reg_module/_01623_ ;
 wire \reg_module/_01624_ ;
 wire \reg_module/_01625_ ;
 wire \reg_module/_01626_ ;
 wire \reg_module/_01627_ ;
 wire \reg_module/_01628_ ;
 wire \reg_module/_01629_ ;
 wire \reg_module/_01630_ ;
 wire \reg_module/_01631_ ;
 wire \reg_module/_01632_ ;
 wire \reg_module/_01633_ ;
 wire \reg_module/_01634_ ;
 wire \reg_module/_01635_ ;
 wire \reg_module/_01636_ ;
 wire \reg_module/_01637_ ;
 wire \reg_module/_01638_ ;
 wire \reg_module/_01639_ ;
 wire \reg_module/_01640_ ;
 wire \reg_module/_01641_ ;
 wire \reg_module/_01642_ ;
 wire \reg_module/_01643_ ;
 wire \reg_module/_01644_ ;
 wire \reg_module/_01645_ ;
 wire \reg_module/_01646_ ;
 wire \reg_module/_01647_ ;
 wire \reg_module/_01648_ ;
 wire \reg_module/_01649_ ;
 wire \reg_module/_01650_ ;
 wire \reg_module/_01651_ ;
 wire \reg_module/_01652_ ;
 wire \reg_module/_01653_ ;
 wire \reg_module/_01654_ ;
 wire \reg_module/_01655_ ;
 wire \reg_module/_01656_ ;
 wire \reg_module/_01657_ ;
 wire \reg_module/_01658_ ;
 wire \reg_module/_01659_ ;
 wire \reg_module/_01660_ ;
 wire \reg_module/_01661_ ;
 wire \reg_module/_01662_ ;
 wire \reg_module/_01663_ ;
 wire \reg_module/_01664_ ;
 wire \reg_module/_01665_ ;
 wire \reg_module/_01666_ ;
 wire \reg_module/_01667_ ;
 wire \reg_module/_01668_ ;
 wire \reg_module/_01669_ ;
 wire \reg_module/_01670_ ;
 wire \reg_module/_01671_ ;
 wire \reg_module/_01672_ ;
 wire \reg_module/_01673_ ;
 wire \reg_module/_01674_ ;
 wire \reg_module/_01675_ ;
 wire \reg_module/_01676_ ;
 wire \reg_module/_01677_ ;
 wire \reg_module/_01678_ ;
 wire \reg_module/_01679_ ;
 wire \reg_module/_01680_ ;
 wire \reg_module/_01681_ ;
 wire \reg_module/_01682_ ;
 wire \reg_module/_01683_ ;
 wire \reg_module/_01684_ ;
 wire \reg_module/_01685_ ;
 wire \reg_module/_01686_ ;
 wire \reg_module/_01687_ ;
 wire \reg_module/_01688_ ;
 wire \reg_module/_01689_ ;
 wire \reg_module/_01690_ ;
 wire \reg_module/_01691_ ;
 wire \reg_module/_01692_ ;
 wire \reg_module/_01693_ ;
 wire \reg_module/_01694_ ;
 wire \reg_module/_01695_ ;
 wire \reg_module/_01696_ ;
 wire \reg_module/_01697_ ;
 wire \reg_module/_01698_ ;
 wire \reg_module/_01699_ ;
 wire \reg_module/_01700_ ;
 wire \reg_module/_01701_ ;
 wire \reg_module/_01702_ ;
 wire \reg_module/_01703_ ;
 wire \reg_module/_01704_ ;
 wire \reg_module/_01705_ ;
 wire \reg_module/_01706_ ;
 wire \reg_module/_01707_ ;
 wire \reg_module/_01708_ ;
 wire \reg_module/_01709_ ;
 wire \reg_module/_01710_ ;
 wire \reg_module/_01711_ ;
 wire \reg_module/_01712_ ;
 wire \reg_module/_01713_ ;
 wire \reg_module/_01714_ ;
 wire \reg_module/_01715_ ;
 wire \reg_module/_01716_ ;
 wire \reg_module/_01717_ ;
 wire \reg_module/_01718_ ;
 wire \reg_module/_01719_ ;
 wire \reg_module/_01720_ ;
 wire \reg_module/_01721_ ;
 wire \reg_module/_01722_ ;
 wire \reg_module/_01723_ ;
 wire \reg_module/_01724_ ;
 wire \reg_module/_01725_ ;
 wire \reg_module/_01726_ ;
 wire \reg_module/_01727_ ;
 wire \reg_module/_01728_ ;
 wire \reg_module/_01729_ ;
 wire \reg_module/_01730_ ;
 wire \reg_module/_01731_ ;
 wire \reg_module/_01732_ ;
 wire \reg_module/_01733_ ;
 wire \reg_module/_01734_ ;
 wire \reg_module/_01735_ ;
 wire \reg_module/_01736_ ;
 wire \reg_module/_01737_ ;
 wire \reg_module/_01738_ ;
 wire \reg_module/_01739_ ;
 wire \reg_module/_01740_ ;
 wire \reg_module/_01741_ ;
 wire \reg_module/_01742_ ;
 wire \reg_module/_01743_ ;
 wire \reg_module/_01744_ ;
 wire \reg_module/_01745_ ;
 wire \reg_module/_01746_ ;
 wire \reg_module/_01747_ ;
 wire \reg_module/_01748_ ;
 wire \reg_module/_01749_ ;
 wire \reg_module/_01750_ ;
 wire \reg_module/_01751_ ;
 wire \reg_module/_01752_ ;
 wire \reg_module/_01753_ ;
 wire \reg_module/_01754_ ;
 wire \reg_module/_01755_ ;
 wire \reg_module/_01756_ ;
 wire \reg_module/_01757_ ;
 wire \reg_module/_01758_ ;
 wire \reg_module/_01759_ ;
 wire \reg_module/_01760_ ;
 wire \reg_module/_01761_ ;
 wire \reg_module/_01762_ ;
 wire \reg_module/_01763_ ;
 wire \reg_module/_01764_ ;
 wire \reg_module/_01765_ ;
 wire \reg_module/_01766_ ;
 wire \reg_module/_01767_ ;
 wire \reg_module/_01768_ ;
 wire \reg_module/_01769_ ;
 wire \reg_module/_01770_ ;
 wire \reg_module/_01771_ ;
 wire \reg_module/_01772_ ;
 wire \reg_module/_01773_ ;
 wire \reg_module/_01774_ ;
 wire \reg_module/_01775_ ;
 wire \reg_module/_01776_ ;
 wire \reg_module/_01777_ ;
 wire \reg_module/_01778_ ;
 wire \reg_module/_01779_ ;
 wire \reg_module/_01780_ ;
 wire \reg_module/_01781_ ;
 wire \reg_module/_01782_ ;
 wire \reg_module/_01783_ ;
 wire \reg_module/_01784_ ;
 wire \reg_module/_01785_ ;
 wire \reg_module/_01786_ ;
 wire \reg_module/_01787_ ;
 wire \reg_module/_01788_ ;
 wire \reg_module/_01789_ ;
 wire \reg_module/_01790_ ;
 wire \reg_module/_01791_ ;
 wire \reg_module/_01792_ ;
 wire \reg_module/_01793_ ;
 wire \reg_module/_01794_ ;
 wire \reg_module/_01795_ ;
 wire \reg_module/_01796_ ;
 wire \reg_module/_01797_ ;
 wire \reg_module/_01798_ ;
 wire \reg_module/_01799_ ;
 wire \reg_module/_01800_ ;
 wire \reg_module/_01801_ ;
 wire \reg_module/_01802_ ;
 wire \reg_module/_01803_ ;
 wire \reg_module/_01804_ ;
 wire \reg_module/_01805_ ;
 wire \reg_module/_01806_ ;
 wire \reg_module/_01807_ ;
 wire \reg_module/_01808_ ;
 wire \reg_module/_01809_ ;
 wire \reg_module/_01810_ ;
 wire \reg_module/_01811_ ;
 wire \reg_module/_01812_ ;
 wire \reg_module/_01813_ ;
 wire \reg_module/_01814_ ;
 wire \reg_module/_01815_ ;
 wire \reg_module/_01816_ ;
 wire \reg_module/_01817_ ;
 wire \reg_module/_01818_ ;
 wire \reg_module/_01819_ ;
 wire \reg_module/_01820_ ;
 wire \reg_module/_01821_ ;
 wire \reg_module/_01822_ ;
 wire \reg_module/_01823_ ;
 wire \reg_module/_01824_ ;
 wire \reg_module/_01825_ ;
 wire \reg_module/_01826_ ;
 wire \reg_module/_01827_ ;
 wire \reg_module/_01828_ ;
 wire \reg_module/_01829_ ;
 wire \reg_module/_01830_ ;
 wire \reg_module/_01831_ ;
 wire \reg_module/_01832_ ;
 wire \reg_module/_01833_ ;
 wire \reg_module/_01834_ ;
 wire \reg_module/_01835_ ;
 wire \reg_module/_01836_ ;
 wire \reg_module/_01837_ ;
 wire \reg_module/_01838_ ;
 wire \reg_module/_01839_ ;
 wire \reg_module/_01840_ ;
 wire \reg_module/_01841_ ;
 wire \reg_module/_01842_ ;
 wire \reg_module/_01843_ ;
 wire \reg_module/_01844_ ;
 wire \reg_module/_01845_ ;
 wire \reg_module/_01846_ ;
 wire \reg_module/_01847_ ;
 wire \reg_module/_01848_ ;
 wire \reg_module/_01849_ ;
 wire \reg_module/_01850_ ;
 wire \reg_module/_01851_ ;
 wire \reg_module/_01852_ ;
 wire \reg_module/_01853_ ;
 wire \reg_module/_01854_ ;
 wire \reg_module/_01855_ ;
 wire \reg_module/_01856_ ;
 wire \reg_module/_01857_ ;
 wire \reg_module/_01858_ ;
 wire \reg_module/_01859_ ;
 wire \reg_module/_01860_ ;
 wire \reg_module/_01861_ ;
 wire \reg_module/_01862_ ;
 wire \reg_module/_01863_ ;
 wire \reg_module/_01864_ ;
 wire \reg_module/_01865_ ;
 wire \reg_module/_01866_ ;
 wire \reg_module/_01867_ ;
 wire \reg_module/_01868_ ;
 wire \reg_module/_01869_ ;
 wire \reg_module/_01870_ ;
 wire \reg_module/_01871_ ;
 wire \reg_module/_01872_ ;
 wire \reg_module/_01873_ ;
 wire \reg_module/_01874_ ;
 wire \reg_module/_01875_ ;
 wire \reg_module/_01876_ ;
 wire \reg_module/_01877_ ;
 wire \reg_module/_01878_ ;
 wire \reg_module/_01879_ ;
 wire \reg_module/_01880_ ;
 wire \reg_module/_01881_ ;
 wire \reg_module/_01882_ ;
 wire \reg_module/_01883_ ;
 wire \reg_module/_01884_ ;
 wire \reg_module/_01885_ ;
 wire \reg_module/_01886_ ;
 wire \reg_module/_01887_ ;
 wire \reg_module/_01888_ ;
 wire \reg_module/_01889_ ;
 wire \reg_module/_01890_ ;
 wire \reg_module/_01891_ ;
 wire \reg_module/_01892_ ;
 wire \reg_module/_01893_ ;
 wire \reg_module/_01894_ ;
 wire \reg_module/_01895_ ;
 wire \reg_module/_01896_ ;
 wire \reg_module/_01897_ ;
 wire \reg_module/_01898_ ;
 wire \reg_module/_01899_ ;
 wire \reg_module/_01900_ ;
 wire \reg_module/_01901_ ;
 wire \reg_module/_01902_ ;
 wire \reg_module/_01903_ ;
 wire \reg_module/_01904_ ;
 wire \reg_module/_01905_ ;
 wire \reg_module/_01906_ ;
 wire \reg_module/_01907_ ;
 wire \reg_module/_01908_ ;
 wire \reg_module/_01909_ ;
 wire \reg_module/_01910_ ;
 wire \reg_module/_01911_ ;
 wire \reg_module/_01912_ ;
 wire \reg_module/_01913_ ;
 wire \reg_module/_01914_ ;
 wire \reg_module/_01915_ ;
 wire \reg_module/_01916_ ;
 wire \reg_module/_01917_ ;
 wire \reg_module/_01918_ ;
 wire \reg_module/_01919_ ;
 wire \reg_module/_01920_ ;
 wire \reg_module/_01921_ ;
 wire \reg_module/_01922_ ;
 wire \reg_module/_01923_ ;
 wire \reg_module/_01924_ ;
 wire \reg_module/_01925_ ;
 wire \reg_module/_01926_ ;
 wire \reg_module/_01927_ ;
 wire \reg_module/_01928_ ;
 wire \reg_module/_01929_ ;
 wire \reg_module/_01930_ ;
 wire \reg_module/_01931_ ;
 wire \reg_module/_01932_ ;
 wire \reg_module/_01933_ ;
 wire \reg_module/_01934_ ;
 wire \reg_module/_01935_ ;
 wire \reg_module/_01936_ ;
 wire \reg_module/_01937_ ;
 wire \reg_module/_01938_ ;
 wire \reg_module/_01939_ ;
 wire \reg_module/_01940_ ;
 wire \reg_module/_01941_ ;
 wire \reg_module/_01942_ ;
 wire \reg_module/_01943_ ;
 wire \reg_module/_01944_ ;
 wire \reg_module/_01945_ ;
 wire \reg_module/_01946_ ;
 wire \reg_module/_01947_ ;
 wire \reg_module/_01948_ ;
 wire \reg_module/_01949_ ;
 wire \reg_module/_01950_ ;
 wire \reg_module/_01951_ ;
 wire \reg_module/_01952_ ;
 wire \reg_module/_01953_ ;
 wire \reg_module/_01954_ ;
 wire \reg_module/_01955_ ;
 wire \reg_module/_01956_ ;
 wire \reg_module/_01957_ ;
 wire \reg_module/_01958_ ;
 wire \reg_module/_01959_ ;
 wire \reg_module/_01960_ ;
 wire \reg_module/_01961_ ;
 wire \reg_module/_01962_ ;
 wire \reg_module/_01963_ ;
 wire \reg_module/_01964_ ;
 wire \reg_module/_01965_ ;
 wire \reg_module/_01966_ ;
 wire \reg_module/_01967_ ;
 wire \reg_module/_01968_ ;
 wire \reg_module/_01969_ ;
 wire \reg_module/_01970_ ;
 wire \reg_module/_01971_ ;
 wire \reg_module/_01972_ ;
 wire \reg_module/_01973_ ;
 wire \reg_module/_01974_ ;
 wire \reg_module/_01975_ ;
 wire \reg_module/_01976_ ;
 wire \reg_module/_01977_ ;
 wire \reg_module/_01978_ ;
 wire \reg_module/_01979_ ;
 wire \reg_module/_01980_ ;
 wire \reg_module/_01981_ ;
 wire \reg_module/_01982_ ;
 wire \reg_module/_01983_ ;
 wire \reg_module/_01984_ ;
 wire \reg_module/_01985_ ;
 wire \reg_module/_01986_ ;
 wire \reg_module/_01987_ ;
 wire \reg_module/_01988_ ;
 wire \reg_module/_01989_ ;
 wire \reg_module/_01990_ ;
 wire \reg_module/_01991_ ;
 wire \reg_module/_01992_ ;
 wire \reg_module/_01993_ ;
 wire \reg_module/_01994_ ;
 wire \reg_module/_01995_ ;
 wire \reg_module/_01996_ ;
 wire \reg_module/_01997_ ;
 wire \reg_module/_01998_ ;
 wire \reg_module/_01999_ ;
 wire \reg_module/_02000_ ;
 wire \reg_module/_02001_ ;
 wire \reg_module/_02002_ ;
 wire \reg_module/_02003_ ;
 wire \reg_module/_02004_ ;
 wire \reg_module/_02005_ ;
 wire \reg_module/_02006_ ;
 wire \reg_module/_02007_ ;
 wire \reg_module/_02008_ ;
 wire \reg_module/_02009_ ;
 wire \reg_module/_02010_ ;
 wire \reg_module/_02011_ ;
 wire \reg_module/_02012_ ;
 wire \reg_module/_02013_ ;
 wire \reg_module/_02014_ ;
 wire \reg_module/_02015_ ;
 wire \reg_module/_02016_ ;
 wire \reg_module/_02017_ ;
 wire \reg_module/_02018_ ;
 wire \reg_module/_02019_ ;
 wire \reg_module/_02020_ ;
 wire \reg_module/_02021_ ;
 wire \reg_module/_02022_ ;
 wire \reg_module/_02023_ ;
 wire \reg_module/_02024_ ;
 wire \reg_module/_02025_ ;
 wire \reg_module/_02026_ ;
 wire \reg_module/_02027_ ;
 wire \reg_module/_02028_ ;
 wire \reg_module/_02029_ ;
 wire \reg_module/_02030_ ;
 wire \reg_module/_02031_ ;
 wire \reg_module/_02032_ ;
 wire \reg_module/_02033_ ;
 wire \reg_module/_02034_ ;
 wire \reg_module/_02035_ ;
 wire \reg_module/_02036_ ;
 wire \reg_module/_02037_ ;
 wire \reg_module/_02038_ ;
 wire \reg_module/_02039_ ;
 wire \reg_module/_02040_ ;
 wire \reg_module/_02041_ ;
 wire \reg_module/_02042_ ;
 wire \reg_module/_02043_ ;
 wire \reg_module/_02044_ ;
 wire \reg_module/_02045_ ;
 wire \reg_module/_02046_ ;
 wire \reg_module/_02047_ ;
 wire \reg_module/_02048_ ;
 wire \reg_module/_02049_ ;
 wire \reg_module/_02050_ ;
 wire \reg_module/_02051_ ;
 wire \reg_module/_02052_ ;
 wire \reg_module/_02053_ ;
 wire \reg_module/_02054_ ;
 wire \reg_module/_02055_ ;
 wire \reg_module/_02056_ ;
 wire \reg_module/_02057_ ;
 wire \reg_module/_02058_ ;
 wire \reg_module/_02059_ ;
 wire \reg_module/_02060_ ;
 wire \reg_module/_02061_ ;
 wire \reg_module/_02062_ ;
 wire \reg_module/_02063_ ;
 wire \reg_module/_02064_ ;
 wire \reg_module/_02065_ ;
 wire \reg_module/_02066_ ;
 wire \reg_module/_02067_ ;
 wire \reg_module/_02068_ ;
 wire \reg_module/_02069_ ;
 wire \reg_module/_02070_ ;
 wire \reg_module/_02071_ ;
 wire \reg_module/_02072_ ;
 wire \reg_module/_02073_ ;
 wire \reg_module/_02074_ ;
 wire \reg_module/_02075_ ;
 wire \reg_module/_02076_ ;
 wire \reg_module/_02077_ ;
 wire \reg_module/_02078_ ;
 wire \reg_module/_02079_ ;
 wire \reg_module/_02080_ ;
 wire \reg_module/_02081_ ;
 wire \reg_module/_02082_ ;
 wire \reg_module/_02083_ ;
 wire \reg_module/_02084_ ;
 wire \reg_module/_02085_ ;
 wire \reg_module/_02086_ ;
 wire \reg_module/_02087_ ;
 wire \reg_module/_02088_ ;
 wire \reg_module/_02089_ ;
 wire \reg_module/_02090_ ;
 wire \reg_module/_02091_ ;
 wire \reg_module/_02092_ ;
 wire \reg_module/_02093_ ;
 wire \reg_module/_02094_ ;
 wire \reg_module/_02095_ ;
 wire \reg_module/_02096_ ;
 wire \reg_module/_02097_ ;
 wire \reg_module/_02098_ ;
 wire \reg_module/_02099_ ;
 wire \reg_module/_02100_ ;
 wire \reg_module/_02101_ ;
 wire \reg_module/_02102_ ;
 wire \reg_module/_02103_ ;
 wire \reg_module/_02104_ ;
 wire \reg_module/_02105_ ;
 wire \reg_module/_02106_ ;
 wire \reg_module/_02107_ ;
 wire \reg_module/_02108_ ;
 wire \reg_module/_02109_ ;
 wire \reg_module/_02110_ ;
 wire \reg_module/_02111_ ;
 wire \reg_module/_02112_ ;
 wire \reg_module/_02113_ ;
 wire \reg_module/_02114_ ;
 wire \reg_module/_02115_ ;
 wire \reg_module/_02116_ ;
 wire \reg_module/_02117_ ;
 wire \reg_module/_02118_ ;
 wire \reg_module/_02119_ ;
 wire \reg_module/_02120_ ;
 wire \reg_module/_02121_ ;
 wire \reg_module/_02122_ ;
 wire \reg_module/_02123_ ;
 wire \reg_module/_02124_ ;
 wire \reg_module/_02125_ ;
 wire \reg_module/_02126_ ;
 wire \reg_module/_02127_ ;
 wire \reg_module/_02128_ ;
 wire \reg_module/_02129_ ;
 wire \reg_module/_02130_ ;
 wire \reg_module/_02131_ ;
 wire \reg_module/_02132_ ;
 wire \reg_module/_02133_ ;
 wire \reg_module/_02134_ ;
 wire \reg_module/_02135_ ;
 wire \reg_module/_02136_ ;
 wire \reg_module/_02137_ ;
 wire \reg_module/_02138_ ;
 wire \reg_module/_02139_ ;
 wire \reg_module/_02140_ ;
 wire \reg_module/_02141_ ;
 wire \reg_module/_02142_ ;
 wire \reg_module/_02143_ ;
 wire \reg_module/_02144_ ;
 wire \reg_module/_02145_ ;
 wire \reg_module/_02146_ ;
 wire \reg_module/_02147_ ;
 wire \reg_module/_02148_ ;
 wire \reg_module/_02149_ ;
 wire \reg_module/_02150_ ;
 wire \reg_module/_02151_ ;
 wire \reg_module/_02152_ ;
 wire \reg_module/_02153_ ;
 wire \reg_module/_02154_ ;
 wire \reg_module/_02155_ ;
 wire \reg_module/_02156_ ;
 wire \reg_module/_02157_ ;
 wire \reg_module/_02158_ ;
 wire \reg_module/_02159_ ;
 wire \reg_module/_02160_ ;
 wire \reg_module/_02161_ ;
 wire \reg_module/_02162_ ;
 wire \reg_module/_02163_ ;
 wire \reg_module/_02164_ ;
 wire \reg_module/_02165_ ;
 wire \reg_module/_02166_ ;
 wire \reg_module/_02167_ ;
 wire \reg_module/_02168_ ;
 wire \reg_module/_02169_ ;
 wire \reg_module/_02170_ ;
 wire \reg_module/_02171_ ;
 wire \reg_module/_02172_ ;
 wire \reg_module/_02173_ ;
 wire \reg_module/_02174_ ;
 wire \reg_module/_02175_ ;
 wire \reg_module/_02176_ ;
 wire \reg_module/_02177_ ;
 wire \reg_module/_02178_ ;
 wire \reg_module/_02179_ ;
 wire \reg_module/_02180_ ;
 wire \reg_module/_02181_ ;
 wire \reg_module/_02182_ ;
 wire \reg_module/_02183_ ;
 wire \reg_module/_02184_ ;
 wire \reg_module/_02185_ ;
 wire \reg_module/_02186_ ;
 wire \reg_module/_02187_ ;
 wire \reg_module/_02188_ ;
 wire \reg_module/_02189_ ;
 wire \reg_module/_02190_ ;
 wire \reg_module/_02191_ ;
 wire \reg_module/_02192_ ;
 wire \reg_module/_02193_ ;
 wire \reg_module/_02194_ ;
 wire \reg_module/_02195_ ;
 wire \reg_module/_02196_ ;
 wire \reg_module/_02197_ ;
 wire \reg_module/_02198_ ;
 wire \reg_module/_02199_ ;
 wire \reg_module/_02200_ ;
 wire \reg_module/_02201_ ;
 wire \reg_module/_02202_ ;
 wire \reg_module/_02203_ ;
 wire \reg_module/_02204_ ;
 wire \reg_module/_02205_ ;
 wire \reg_module/_02206_ ;
 wire \reg_module/_02207_ ;
 wire \reg_module/_02208_ ;
 wire \reg_module/_02209_ ;
 wire \reg_module/_02210_ ;
 wire \reg_module/_02211_ ;
 wire \reg_module/_02212_ ;
 wire \reg_module/_02213_ ;
 wire \reg_module/_02214_ ;
 wire \reg_module/_02215_ ;
 wire \reg_module/_02216_ ;
 wire \reg_module/_02217_ ;
 wire \reg_module/_02218_ ;
 wire \reg_module/_02219_ ;
 wire \reg_module/_02220_ ;
 wire \reg_module/_02221_ ;
 wire \reg_module/_02222_ ;
 wire \reg_module/_02223_ ;
 wire \reg_module/_02224_ ;
 wire \reg_module/_02225_ ;
 wire \reg_module/_02226_ ;
 wire \reg_module/_02227_ ;
 wire \reg_module/_02228_ ;
 wire \reg_module/_02229_ ;
 wire \reg_module/_02230_ ;
 wire \reg_module/_02231_ ;
 wire \reg_module/_02232_ ;
 wire \reg_module/_02233_ ;
 wire \reg_module/_02234_ ;
 wire \reg_module/_02235_ ;
 wire \reg_module/_02236_ ;
 wire \reg_module/_02237_ ;
 wire \reg_module/_02238_ ;
 wire \reg_module/_02239_ ;
 wire \reg_module/_02240_ ;
 wire \reg_module/_02241_ ;
 wire \reg_module/_02242_ ;
 wire \reg_module/_02243_ ;
 wire \reg_module/_02244_ ;
 wire \reg_module/_02245_ ;
 wire \reg_module/_02246_ ;
 wire \reg_module/_02247_ ;
 wire \reg_module/_02248_ ;
 wire \reg_module/_02249_ ;
 wire \reg_module/_02250_ ;
 wire \reg_module/_02251_ ;
 wire \reg_module/_02252_ ;
 wire \reg_module/_02253_ ;
 wire \reg_module/_02254_ ;
 wire \reg_module/_02255_ ;
 wire \reg_module/_02256_ ;
 wire \reg_module/_02257_ ;
 wire \reg_module/_02258_ ;
 wire \reg_module/_02259_ ;
 wire \reg_module/_02260_ ;
 wire \reg_module/_02261_ ;
 wire \reg_module/_02262_ ;
 wire \reg_module/_02263_ ;
 wire \reg_module/_02264_ ;
 wire \reg_module/_02265_ ;
 wire \reg_module/_02266_ ;
 wire \reg_module/_02267_ ;
 wire \reg_module/_02268_ ;
 wire \reg_module/_02269_ ;
 wire \reg_module/_02270_ ;
 wire \reg_module/_02271_ ;
 wire \reg_module/_02272_ ;
 wire \reg_module/_02273_ ;
 wire \reg_module/_02274_ ;
 wire \reg_module/_02275_ ;
 wire \reg_module/_02276_ ;
 wire \reg_module/_02277_ ;
 wire \reg_module/_02278_ ;
 wire \reg_module/_02279_ ;
 wire \reg_module/_02280_ ;
 wire \reg_module/_02281_ ;
 wire \reg_module/_02282_ ;
 wire \reg_module/_02283_ ;
 wire \reg_module/_02284_ ;
 wire \reg_module/_02285_ ;
 wire \reg_module/_02286_ ;
 wire \reg_module/_02287_ ;
 wire \reg_module/_02288_ ;
 wire \reg_module/_02289_ ;
 wire \reg_module/_02290_ ;
 wire \reg_module/_02291_ ;
 wire \reg_module/_02292_ ;
 wire \reg_module/_02293_ ;
 wire \reg_module/_02294_ ;
 wire \reg_module/_02295_ ;
 wire \reg_module/_02296_ ;
 wire \reg_module/_02297_ ;
 wire \reg_module/_02298_ ;
 wire \reg_module/_02299_ ;
 wire \reg_module/_02300_ ;
 wire \reg_module/_02301_ ;
 wire \reg_module/_02302_ ;
 wire \reg_module/_02303_ ;
 wire \reg_module/_02304_ ;
 wire \reg_module/_02305_ ;
 wire \reg_module/_02306_ ;
 wire \reg_module/_02307_ ;
 wire \reg_module/_02308_ ;
 wire \reg_module/_02309_ ;
 wire \reg_module/_02310_ ;
 wire \reg_module/_02311_ ;
 wire \reg_module/_02312_ ;
 wire \reg_module/_02313_ ;
 wire \reg_module/_02314_ ;
 wire \reg_module/_02315_ ;
 wire \reg_module/_02316_ ;
 wire \reg_module/_02317_ ;
 wire \reg_module/_02318_ ;
 wire \reg_module/_02319_ ;
 wire \reg_module/_02320_ ;
 wire \reg_module/_02321_ ;
 wire \reg_module/_02322_ ;
 wire \reg_module/_02323_ ;
 wire \reg_module/_02324_ ;
 wire \reg_module/_02325_ ;
 wire \reg_module/_02326_ ;
 wire \reg_module/_02327_ ;
 wire \reg_module/_02328_ ;
 wire \reg_module/_02329_ ;
 wire \reg_module/_02330_ ;
 wire \reg_module/_02331_ ;
 wire \reg_module/_02332_ ;
 wire \reg_module/_02333_ ;
 wire \reg_module/_02334_ ;
 wire \reg_module/_02335_ ;
 wire \reg_module/_02336_ ;
 wire \reg_module/_02337_ ;
 wire \reg_module/_02338_ ;
 wire \reg_module/_02339_ ;
 wire \reg_module/_02340_ ;
 wire \reg_module/_02341_ ;
 wire \reg_module/_02342_ ;
 wire \reg_module/_02343_ ;
 wire \reg_module/_02344_ ;
 wire \reg_module/_02345_ ;
 wire \reg_module/_02346_ ;
 wire \reg_module/_02347_ ;
 wire \reg_module/_02348_ ;
 wire \reg_module/_02349_ ;
 wire \reg_module/_02350_ ;
 wire \reg_module/_02351_ ;
 wire \reg_module/_02352_ ;
 wire \reg_module/_02353_ ;
 wire \reg_module/_02354_ ;
 wire \reg_module/_02355_ ;
 wire \reg_module/_02356_ ;
 wire \reg_module/_02357_ ;
 wire \reg_module/_02358_ ;
 wire \reg_module/_02359_ ;
 wire \reg_module/_02360_ ;
 wire \reg_module/_02361_ ;
 wire \reg_module/_02362_ ;
 wire \reg_module/_02363_ ;
 wire \reg_module/_02364_ ;
 wire \reg_module/_02365_ ;
 wire \reg_module/_02366_ ;
 wire \reg_module/_02367_ ;
 wire \reg_module/_02368_ ;
 wire \reg_module/_02369_ ;
 wire \reg_module/_02370_ ;
 wire \reg_module/_02371_ ;
 wire \reg_module/_02372_ ;
 wire \reg_module/_02373_ ;
 wire \reg_module/_02374_ ;
 wire \reg_module/_02375_ ;
 wire \reg_module/_02376_ ;
 wire \reg_module/_02377_ ;
 wire \reg_module/_02378_ ;
 wire \reg_module/_02379_ ;
 wire \reg_module/_02380_ ;
 wire \reg_module/_02381_ ;
 wire \reg_module/_02382_ ;
 wire \reg_module/_02383_ ;
 wire \reg_module/_02384_ ;
 wire \reg_module/_02385_ ;
 wire \reg_module/_02386_ ;
 wire \reg_module/_02387_ ;
 wire \reg_module/_02388_ ;
 wire \reg_module/_02389_ ;
 wire \reg_module/_02390_ ;
 wire \reg_module/_02391_ ;
 wire \reg_module/_02392_ ;
 wire \reg_module/_02393_ ;
 wire \reg_module/_02394_ ;
 wire \reg_module/_02395_ ;
 wire \reg_module/_02396_ ;
 wire \reg_module/_02397_ ;
 wire \reg_module/_02398_ ;
 wire \reg_module/_02399_ ;
 wire \reg_module/_02400_ ;
 wire \reg_module/_02401_ ;
 wire \reg_module/_02402_ ;
 wire \reg_module/_02403_ ;
 wire \reg_module/_02404_ ;
 wire \reg_module/_02405_ ;
 wire \reg_module/_02406_ ;
 wire \reg_module/_02407_ ;
 wire \reg_module/_02408_ ;
 wire \reg_module/_02409_ ;
 wire \reg_module/_02410_ ;
 wire \reg_module/_02411_ ;
 wire \reg_module/_02412_ ;
 wire \reg_module/_02413_ ;
 wire \reg_module/_02414_ ;
 wire \reg_module/_02415_ ;
 wire \reg_module/_02416_ ;
 wire \reg_module/_02417_ ;
 wire \reg_module/_02418_ ;
 wire \reg_module/_02419_ ;
 wire \reg_module/_02420_ ;
 wire \reg_module/_02421_ ;
 wire \reg_module/_02422_ ;
 wire \reg_module/_02423_ ;
 wire \reg_module/_02424_ ;
 wire \reg_module/_02425_ ;
 wire \reg_module/_02426_ ;
 wire \reg_module/_02427_ ;
 wire \reg_module/_02428_ ;
 wire \reg_module/_02429_ ;
 wire \reg_module/_02430_ ;
 wire \reg_module/_02431_ ;
 wire \reg_module/_02432_ ;
 wire \reg_module/_02433_ ;
 wire \reg_module/_02434_ ;
 wire \reg_module/_02435_ ;
 wire \reg_module/_02436_ ;
 wire \reg_module/_02437_ ;
 wire \reg_module/_02438_ ;
 wire \reg_module/_02439_ ;
 wire \reg_module/_02440_ ;
 wire \reg_module/_02441_ ;
 wire \reg_module/_02442_ ;
 wire \reg_module/_02443_ ;
 wire \reg_module/_02444_ ;
 wire \reg_module/_02445_ ;
 wire \reg_module/_02446_ ;
 wire \reg_module/_02447_ ;
 wire \reg_module/_02448_ ;
 wire \reg_module/_02449_ ;
 wire \reg_module/_02450_ ;
 wire \reg_module/_02451_ ;
 wire \reg_module/_02452_ ;
 wire \reg_module/_02453_ ;
 wire \reg_module/_02454_ ;
 wire \reg_module/_02455_ ;
 wire \reg_module/_02456_ ;
 wire \reg_module/_02457_ ;
 wire \reg_module/_02458_ ;
 wire \reg_module/_02459_ ;
 wire \reg_module/_02460_ ;
 wire \reg_module/_02461_ ;
 wire \reg_module/_02462_ ;
 wire \reg_module/_02463_ ;
 wire \reg_module/_02464_ ;
 wire \reg_module/_02465_ ;
 wire \reg_module/_02466_ ;
 wire \reg_module/_02467_ ;
 wire \reg_module/_02468_ ;
 wire \reg_module/_02469_ ;
 wire \reg_module/_02470_ ;
 wire \reg_module/_02471_ ;
 wire \reg_module/_02472_ ;
 wire \reg_module/_02473_ ;
 wire \reg_module/_02474_ ;
 wire \reg_module/_02475_ ;
 wire \reg_module/_02476_ ;
 wire \reg_module/_02477_ ;
 wire \reg_module/_02478_ ;
 wire \reg_module/_02479_ ;
 wire \reg_module/_02480_ ;
 wire \reg_module/_02481_ ;
 wire \reg_module/_02482_ ;
 wire \reg_module/_02483_ ;
 wire \reg_module/_02484_ ;
 wire \reg_module/_02485_ ;
 wire \reg_module/_02486_ ;
 wire \reg_module/_02487_ ;
 wire \reg_module/_02488_ ;
 wire \reg_module/_02489_ ;
 wire \reg_module/_02490_ ;
 wire \reg_module/_02491_ ;
 wire \reg_module/_02492_ ;
 wire \reg_module/_02493_ ;
 wire \reg_module/_02494_ ;
 wire \reg_module/_02495_ ;
 wire \reg_module/_02496_ ;
 wire \reg_module/_02497_ ;
 wire \reg_module/_02498_ ;
 wire \reg_module/_02499_ ;
 wire \reg_module/_02500_ ;
 wire \reg_module/_02501_ ;
 wire \reg_module/_02502_ ;
 wire \reg_module/_02503_ ;
 wire \reg_module/_02504_ ;
 wire \reg_module/_02505_ ;
 wire \reg_module/_02506_ ;
 wire \reg_module/_02507_ ;
 wire \reg_module/_02508_ ;
 wire \reg_module/_02509_ ;
 wire \reg_module/_02510_ ;
 wire \reg_module/_02511_ ;
 wire \reg_module/_02512_ ;
 wire \reg_module/_02513_ ;
 wire \reg_module/_02514_ ;
 wire \reg_module/_02515_ ;
 wire \reg_module/_02516_ ;
 wire \reg_module/_02517_ ;
 wire \reg_module/_02518_ ;
 wire \reg_module/_02519_ ;
 wire \reg_module/_02520_ ;
 wire \reg_module/_02521_ ;
 wire \reg_module/_02522_ ;
 wire \reg_module/_02523_ ;
 wire \reg_module/_02524_ ;
 wire \reg_module/_02525_ ;
 wire \reg_module/_02526_ ;
 wire \reg_module/_02527_ ;
 wire \reg_module/_02528_ ;
 wire \reg_module/_02529_ ;
 wire \reg_module/_02530_ ;
 wire \reg_module/_02531_ ;
 wire \reg_module/_02532_ ;
 wire \reg_module/_02533_ ;
 wire \reg_module/_02534_ ;
 wire \reg_module/_02535_ ;
 wire \reg_module/_02536_ ;
 wire \reg_module/_02537_ ;
 wire \reg_module/_02538_ ;
 wire \reg_module/_02539_ ;
 wire \reg_module/_02540_ ;
 wire \reg_module/_02541_ ;
 wire \reg_module/_02542_ ;
 wire \reg_module/_02543_ ;
 wire \reg_module/_02544_ ;
 wire \reg_module/_02545_ ;
 wire \reg_module/_02546_ ;
 wire \reg_module/_02547_ ;
 wire \reg_module/_02548_ ;
 wire \reg_module/_02549_ ;
 wire \reg_module/_02550_ ;
 wire \reg_module/_02551_ ;
 wire \reg_module/_02552_ ;
 wire \reg_module/_02553_ ;
 wire \reg_module/_02554_ ;
 wire \reg_module/_02555_ ;
 wire \reg_module/_02556_ ;
 wire \reg_module/_02557_ ;
 wire \reg_module/_02558_ ;
 wire \reg_module/_02559_ ;
 wire \reg_module/_02560_ ;
 wire \reg_module/_02561_ ;
 wire \reg_module/_02562_ ;
 wire \reg_module/_02563_ ;
 wire \reg_module/_02564_ ;
 wire \reg_module/_02565_ ;
 wire \reg_module/_02566_ ;
 wire \reg_module/_02567_ ;
 wire \reg_module/_02568_ ;
 wire \reg_module/_02569_ ;
 wire \reg_module/_02570_ ;
 wire \reg_module/_02571_ ;
 wire \reg_module/_02572_ ;
 wire \reg_module/_02573_ ;
 wire \reg_module/_02574_ ;
 wire \reg_module/_02575_ ;
 wire \reg_module/_02576_ ;
 wire \reg_module/_02577_ ;
 wire \reg_module/_02578_ ;
 wire \reg_module/_02579_ ;
 wire \reg_module/_02580_ ;
 wire \reg_module/_02581_ ;
 wire \reg_module/_02582_ ;
 wire \reg_module/_02583_ ;
 wire \reg_module/_02584_ ;
 wire \reg_module/_02585_ ;
 wire \reg_module/_02586_ ;
 wire \reg_module/_02587_ ;
 wire \reg_module/_02588_ ;
 wire \reg_module/_02589_ ;
 wire \reg_module/_02590_ ;
 wire \reg_module/_02591_ ;
 wire \reg_module/_02592_ ;
 wire \reg_module/_02593_ ;
 wire \reg_module/_02594_ ;
 wire \reg_module/_02595_ ;
 wire \reg_module/_02596_ ;
 wire \reg_module/_02597_ ;
 wire \reg_module/_02598_ ;
 wire \reg_module/_02599_ ;
 wire \reg_module/_02600_ ;
 wire \reg_module/_02601_ ;
 wire \reg_module/_02602_ ;
 wire \reg_module/_02603_ ;
 wire \reg_module/_02604_ ;
 wire \reg_module/_02605_ ;
 wire \reg_module/_02606_ ;
 wire \reg_module/_02607_ ;
 wire \reg_module/_02608_ ;
 wire \reg_module/_02609_ ;
 wire \reg_module/_02610_ ;
 wire \reg_module/_02611_ ;
 wire \reg_module/_02612_ ;
 wire \reg_module/_02613_ ;
 wire \reg_module/_02614_ ;
 wire \reg_module/_02615_ ;
 wire \reg_module/_02616_ ;
 wire \reg_module/_02617_ ;
 wire \reg_module/_02618_ ;
 wire \reg_module/_02619_ ;
 wire \reg_module/_02620_ ;
 wire \reg_module/_02621_ ;
 wire \reg_module/_02622_ ;
 wire \reg_module/_02623_ ;
 wire \reg_module/_02624_ ;
 wire \reg_module/_02625_ ;
 wire \reg_module/_02626_ ;
 wire \reg_module/_02627_ ;
 wire \reg_module/_02628_ ;
 wire \reg_module/_02629_ ;
 wire \reg_module/_02630_ ;
 wire \reg_module/_02631_ ;
 wire \reg_module/_02632_ ;
 wire \reg_module/_02633_ ;
 wire \reg_module/_02634_ ;
 wire \reg_module/_02635_ ;
 wire \reg_module/_02636_ ;
 wire \reg_module/_02637_ ;
 wire \reg_module/_02638_ ;
 wire \reg_module/_02639_ ;
 wire \reg_module/_02640_ ;
 wire \reg_module/_02641_ ;
 wire \reg_module/_02642_ ;
 wire \reg_module/_02643_ ;
 wire \reg_module/_02644_ ;
 wire \reg_module/_02645_ ;
 wire \reg_module/_02646_ ;
 wire \reg_module/_02647_ ;
 wire \reg_module/_02648_ ;
 wire \reg_module/_02649_ ;
 wire \reg_module/_02650_ ;
 wire \reg_module/_02651_ ;
 wire \reg_module/_02652_ ;
 wire \reg_module/_02653_ ;
 wire \reg_module/_02654_ ;
 wire \reg_module/_02655_ ;
 wire \reg_module/_02656_ ;
 wire \reg_module/_02657_ ;
 wire \reg_module/_02658_ ;
 wire \reg_module/_02659_ ;
 wire \reg_module/_02660_ ;
 wire \reg_module/_02661_ ;
 wire \reg_module/_02662_ ;
 wire \reg_module/_02663_ ;
 wire \reg_module/_02664_ ;
 wire \reg_module/_02665_ ;
 wire \reg_module/_02666_ ;
 wire \reg_module/_02667_ ;
 wire \reg_module/_02668_ ;
 wire \reg_module/_02669_ ;
 wire \reg_module/_02670_ ;
 wire \reg_module/_02671_ ;
 wire \reg_module/_02672_ ;
 wire \reg_module/_02673_ ;
 wire \reg_module/_02674_ ;
 wire \reg_module/_02675_ ;
 wire \reg_module/_02676_ ;
 wire \reg_module/_02677_ ;
 wire \reg_module/_02678_ ;
 wire \reg_module/_02679_ ;
 wire \reg_module/_02680_ ;
 wire \reg_module/_02681_ ;
 wire \reg_module/_02682_ ;
 wire \reg_module/_02683_ ;
 wire \reg_module/_02684_ ;
 wire \reg_module/_02685_ ;
 wire \reg_module/_02686_ ;
 wire \reg_module/_02687_ ;
 wire \reg_module/_02688_ ;
 wire \reg_module/_02689_ ;
 wire \reg_module/_02690_ ;
 wire \reg_module/_02691_ ;
 wire \reg_module/_02692_ ;
 wire \reg_module/_02693_ ;
 wire \reg_module/_02694_ ;
 wire \reg_module/_02695_ ;
 wire \reg_module/_02696_ ;
 wire \reg_module/_02697_ ;
 wire \reg_module/_02698_ ;
 wire \reg_module/_02699_ ;
 wire \reg_module/_02700_ ;
 wire \reg_module/_02701_ ;
 wire \reg_module/_02702_ ;
 wire \reg_module/_02703_ ;
 wire \reg_module/_02704_ ;
 wire \reg_module/_02705_ ;
 wire \reg_module/_02706_ ;
 wire \reg_module/_02707_ ;
 wire \reg_module/_02708_ ;
 wire \reg_module/_02709_ ;
 wire \reg_module/_02710_ ;
 wire \reg_module/_02711_ ;
 wire \reg_module/_02712_ ;
 wire \reg_module/_02713_ ;
 wire \reg_module/_02714_ ;
 wire \reg_module/_02715_ ;
 wire \reg_module/_02716_ ;
 wire \reg_module/_02717_ ;
 wire \reg_module/_02718_ ;
 wire \reg_module/_02719_ ;
 wire \reg_module/_02720_ ;
 wire \reg_module/_02721_ ;
 wire \reg_module/_02722_ ;
 wire \reg_module/_02723_ ;
 wire \reg_module/_02724_ ;
 wire \reg_module/_02725_ ;
 wire \reg_module/_02726_ ;
 wire \reg_module/_02727_ ;
 wire \reg_module/_02728_ ;
 wire \reg_module/_02729_ ;
 wire \reg_module/_02730_ ;
 wire \reg_module/_02731_ ;
 wire \reg_module/_02732_ ;
 wire \reg_module/_02733_ ;
 wire \reg_module/_02734_ ;
 wire \reg_module/_02735_ ;
 wire \reg_module/_02736_ ;
 wire \reg_module/_02737_ ;
 wire \reg_module/_02738_ ;
 wire \reg_module/_02739_ ;
 wire \reg_module/_02740_ ;
 wire \reg_module/_02741_ ;
 wire \reg_module/_02742_ ;
 wire \reg_module/_02743_ ;
 wire \reg_module/_02744_ ;
 wire \reg_module/_02745_ ;
 wire \reg_module/_02746_ ;
 wire \reg_module/_02747_ ;
 wire \reg_module/_02748_ ;
 wire \reg_module/_02749_ ;
 wire \reg_module/_02750_ ;
 wire \reg_module/_02751_ ;
 wire \reg_module/_02752_ ;
 wire \reg_module/_02753_ ;
 wire \reg_module/_02754_ ;
 wire \reg_module/_02755_ ;
 wire \reg_module/_02756_ ;
 wire \reg_module/_02757_ ;
 wire \reg_module/_02758_ ;
 wire \reg_module/_02759_ ;
 wire \reg_module/_02760_ ;
 wire \reg_module/_02761_ ;
 wire \reg_module/_02762_ ;
 wire \reg_module/_02763_ ;
 wire \reg_module/_02764_ ;
 wire \reg_module/_02765_ ;
 wire \reg_module/_02766_ ;
 wire \reg_module/_02767_ ;
 wire \reg_module/_02768_ ;
 wire \reg_module/_02769_ ;
 wire \reg_module/_02770_ ;
 wire \reg_module/_02771_ ;
 wire \reg_module/_02772_ ;
 wire \reg_module/_02773_ ;
 wire \reg_module/_02774_ ;
 wire \reg_module/_02775_ ;
 wire \reg_module/_02776_ ;
 wire \reg_module/_02777_ ;
 wire \reg_module/_02778_ ;
 wire \reg_module/_02779_ ;
 wire \reg_module/_02780_ ;
 wire \reg_module/_02781_ ;
 wire \reg_module/_02782_ ;
 wire \reg_module/_02783_ ;
 wire \reg_module/_02784_ ;
 wire \reg_module/_02785_ ;
 wire \reg_module/_02786_ ;
 wire \reg_module/_02787_ ;
 wire \reg_module/_02788_ ;
 wire \reg_module/_02789_ ;
 wire \reg_module/_02790_ ;
 wire \reg_module/_02791_ ;
 wire \reg_module/_02792_ ;
 wire \reg_module/_02793_ ;
 wire \reg_module/_02794_ ;
 wire \reg_module/_02795_ ;
 wire \reg_module/_02796_ ;
 wire \reg_module/_02797_ ;
 wire \reg_module/_02798_ ;
 wire \reg_module/_02799_ ;
 wire \reg_module/_02800_ ;
 wire \reg_module/_02801_ ;
 wire \reg_module/_02802_ ;
 wire \reg_module/_02803_ ;
 wire \reg_module/_02804_ ;
 wire \reg_module/_02805_ ;
 wire \reg_module/_02806_ ;
 wire \reg_module/_02807_ ;
 wire \reg_module/_02808_ ;
 wire \reg_module/_02809_ ;
 wire \reg_module/_02810_ ;
 wire \reg_module/_02811_ ;
 wire \reg_module/_02812_ ;
 wire \reg_module/_02813_ ;
 wire \reg_module/_02814_ ;
 wire \reg_module/_02815_ ;
 wire \reg_module/_02816_ ;
 wire \reg_module/_02817_ ;
 wire \reg_module/_02818_ ;
 wire \reg_module/_02819_ ;
 wire \reg_module/_02820_ ;
 wire \reg_module/_02821_ ;
 wire \reg_module/_02822_ ;
 wire \reg_module/_02823_ ;
 wire \reg_module/_02824_ ;
 wire \reg_module/_02825_ ;
 wire \reg_module/_02826_ ;
 wire \reg_module/_02827_ ;
 wire \reg_module/_02828_ ;
 wire \reg_module/_02829_ ;
 wire \reg_module/_02830_ ;
 wire \reg_module/_02831_ ;
 wire \reg_module/_02832_ ;
 wire \reg_module/_02833_ ;
 wire \reg_module/_02834_ ;
 wire \reg_module/_02835_ ;
 wire \reg_module/_02836_ ;
 wire \reg_module/_02837_ ;
 wire \reg_module/_02838_ ;
 wire \reg_module/_02839_ ;
 wire \reg_module/_02840_ ;
 wire \reg_module/_02841_ ;
 wire \reg_module/_02842_ ;
 wire \reg_module/_02843_ ;
 wire \reg_module/_02844_ ;
 wire \reg_module/_02845_ ;
 wire \reg_module/_02846_ ;
 wire \reg_module/_02847_ ;
 wire \reg_module/_02848_ ;
 wire \reg_module/_02849_ ;
 wire \reg_module/_02850_ ;
 wire \reg_module/_02851_ ;
 wire \reg_module/_02852_ ;
 wire \reg_module/_02853_ ;
 wire \reg_module/_02854_ ;
 wire \reg_module/_02855_ ;
 wire \reg_module/_02856_ ;
 wire \reg_module/_02857_ ;
 wire \reg_module/_02858_ ;
 wire \reg_module/_02859_ ;
 wire \reg_module/_02860_ ;
 wire \reg_module/_02861_ ;
 wire \reg_module/_02862_ ;
 wire \reg_module/_02863_ ;
 wire \reg_module/_02864_ ;
 wire \reg_module/_02865_ ;
 wire \reg_module/_02866_ ;
 wire \reg_module/_02867_ ;
 wire \reg_module/_02868_ ;
 wire \reg_module/_02869_ ;
 wire \reg_module/_02870_ ;
 wire \reg_module/_02871_ ;
 wire \reg_module/_02872_ ;
 wire \reg_module/_02873_ ;
 wire \reg_module/_02874_ ;
 wire \reg_module/_02875_ ;
 wire \reg_module/_02876_ ;
 wire \reg_module/_02877_ ;
 wire \reg_module/_02878_ ;
 wire \reg_module/_02879_ ;
 wire \reg_module/_02880_ ;
 wire \reg_module/_02881_ ;
 wire \reg_module/_02882_ ;
 wire \reg_module/_02883_ ;
 wire \reg_module/_02884_ ;
 wire \reg_module/_02885_ ;
 wire \reg_module/_02886_ ;
 wire \reg_module/_02887_ ;
 wire \reg_module/_02888_ ;
 wire \reg_module/_02889_ ;
 wire \reg_module/_02890_ ;
 wire \reg_module/_02891_ ;
 wire \reg_module/_02892_ ;
 wire \reg_module/_02893_ ;
 wire \reg_module/_02894_ ;
 wire \reg_module/_02895_ ;
 wire \reg_module/_02896_ ;
 wire \reg_module/_02897_ ;
 wire \reg_module/_02898_ ;
 wire \reg_module/_02899_ ;
 wire \reg_module/_02900_ ;
 wire \reg_module/_02901_ ;
 wire \reg_module/_02902_ ;
 wire \reg_module/_02903_ ;
 wire \reg_module/_02904_ ;
 wire \reg_module/_02905_ ;
 wire \reg_module/_02906_ ;
 wire \reg_module/_02907_ ;
 wire \reg_module/_02908_ ;
 wire \reg_module/_02909_ ;
 wire \reg_module/_02910_ ;
 wire \reg_module/_02911_ ;
 wire \reg_module/_02912_ ;
 wire \reg_module/_02913_ ;
 wire \reg_module/_02914_ ;
 wire \reg_module/_02915_ ;
 wire \reg_module/_02916_ ;
 wire \reg_module/_02917_ ;
 wire \reg_module/_02918_ ;
 wire \reg_module/_02919_ ;
 wire \reg_module/_02920_ ;
 wire \reg_module/_02921_ ;
 wire \reg_module/_02922_ ;
 wire \reg_module/_02923_ ;
 wire \reg_module/_02924_ ;
 wire \reg_module/_02925_ ;
 wire \reg_module/_02926_ ;
 wire \reg_module/_02927_ ;
 wire \reg_module/_02928_ ;
 wire \reg_module/_02929_ ;
 wire \reg_module/_02930_ ;
 wire \reg_module/_02931_ ;
 wire \reg_module/_02932_ ;
 wire \reg_module/_02933_ ;
 wire \reg_module/_02934_ ;
 wire \reg_module/_02935_ ;
 wire \reg_module/_02936_ ;
 wire \reg_module/_02937_ ;
 wire \reg_module/_02938_ ;
 wire \reg_module/_02939_ ;
 wire \reg_module/_02940_ ;
 wire \reg_module/_02941_ ;
 wire \reg_module/_02942_ ;
 wire \reg_module/_02943_ ;
 wire \reg_module/_02944_ ;
 wire \reg_module/_02945_ ;
 wire \reg_module/_02946_ ;
 wire \reg_module/_02947_ ;
 wire \reg_module/_02948_ ;
 wire \reg_module/_02949_ ;
 wire \reg_module/_02950_ ;
 wire \reg_module/_02951_ ;
 wire \reg_module/_02952_ ;
 wire \reg_module/_02953_ ;
 wire \reg_module/_02954_ ;
 wire \reg_module/_02955_ ;
 wire \reg_module/_02956_ ;
 wire \reg_module/_02957_ ;
 wire \reg_module/_02958_ ;
 wire \reg_module/_02959_ ;
 wire \reg_module/_02960_ ;
 wire \reg_module/_02961_ ;
 wire \reg_module/_02962_ ;
 wire \reg_module/_02963_ ;
 wire \reg_module/_02964_ ;
 wire \reg_module/_02965_ ;
 wire \reg_module/_02966_ ;
 wire \reg_module/_02967_ ;
 wire \reg_module/_02968_ ;
 wire \reg_module/_02969_ ;
 wire \reg_module/_02970_ ;
 wire \reg_module/_02971_ ;
 wire \reg_module/_02972_ ;
 wire \reg_module/_02973_ ;
 wire \reg_module/_02974_ ;
 wire \reg_module/_02975_ ;
 wire \reg_module/_02976_ ;
 wire \reg_module/_02977_ ;
 wire \reg_module/_02978_ ;
 wire \reg_module/_02979_ ;
 wire \reg_module/_02980_ ;
 wire \reg_module/_02981_ ;
 wire \reg_module/_02982_ ;
 wire \reg_module/_02983_ ;
 wire \reg_module/_02984_ ;
 wire \reg_module/_02985_ ;
 wire \reg_module/_02986_ ;
 wire \reg_module/_02987_ ;
 wire \reg_module/_02988_ ;
 wire \reg_module/_02989_ ;
 wire \reg_module/_02990_ ;
 wire \reg_module/_02991_ ;
 wire \reg_module/_02992_ ;
 wire \reg_module/_02993_ ;
 wire \reg_module/_02994_ ;
 wire \reg_module/_02995_ ;
 wire \reg_module/_02996_ ;
 wire \reg_module/_02997_ ;
 wire \reg_module/_02998_ ;
 wire \reg_module/_02999_ ;
 wire \reg_module/_03000_ ;
 wire \reg_module/_03001_ ;
 wire \reg_module/_03002_ ;
 wire \reg_module/_03003_ ;
 wire \reg_module/_03004_ ;
 wire \reg_module/_03005_ ;
 wire \reg_module/_03006_ ;
 wire \reg_module/_03007_ ;
 wire \reg_module/_03008_ ;
 wire \reg_module/_03009_ ;
 wire \reg_module/_03010_ ;
 wire \reg_module/_03011_ ;
 wire \reg_module/_03012_ ;
 wire \reg_module/_03013_ ;
 wire \reg_module/_03014_ ;
 wire \reg_module/_03015_ ;
 wire \reg_module/_03016_ ;
 wire \reg_module/_03017_ ;
 wire \reg_module/_03018_ ;
 wire \reg_module/_03019_ ;
 wire \reg_module/_03020_ ;
 wire \reg_module/_03021_ ;
 wire \reg_module/_03022_ ;
 wire \reg_module/_03023_ ;
 wire \reg_module/_03024_ ;
 wire \reg_module/_03025_ ;
 wire \reg_module/_03026_ ;
 wire \reg_module/_03027_ ;
 wire \reg_module/_03028_ ;
 wire \reg_module/_03029_ ;
 wire \reg_module/_03030_ ;
 wire \reg_module/_03031_ ;
 wire \reg_module/_03032_ ;
 wire \reg_module/_03033_ ;
 wire \reg_module/_03034_ ;
 wire \reg_module/_03035_ ;
 wire \reg_module/_03036_ ;
 wire \reg_module/_03037_ ;
 wire \reg_module/_03038_ ;
 wire \reg_module/_03039_ ;
 wire \reg_module/_03040_ ;
 wire \reg_module/_03041_ ;
 wire \reg_module/_03042_ ;
 wire \reg_module/_03043_ ;
 wire \reg_module/_03044_ ;
 wire \reg_module/_03045_ ;
 wire \reg_module/_03046_ ;
 wire \reg_module/_03047_ ;
 wire \reg_module/_03048_ ;
 wire \reg_module/_03049_ ;
 wire \reg_module/_03050_ ;
 wire \reg_module/_03051_ ;
 wire \reg_module/_03052_ ;
 wire \reg_module/_03053_ ;
 wire \reg_module/_03054_ ;
 wire \reg_module/_03055_ ;
 wire \reg_module/_03056_ ;
 wire \reg_module/_03057_ ;
 wire \reg_module/_03058_ ;
 wire \reg_module/_03059_ ;
 wire \reg_module/_03060_ ;
 wire \reg_module/_03061_ ;
 wire \reg_module/_03062_ ;
 wire \reg_module/_03063_ ;
 wire \reg_module/_03064_ ;
 wire \reg_module/_03065_ ;
 wire \reg_module/_03066_ ;
 wire \reg_module/_03067_ ;
 wire \reg_module/_03068_ ;
 wire \reg_module/_03069_ ;
 wire \reg_module/_03070_ ;
 wire \reg_module/_03071_ ;
 wire \reg_module/_03072_ ;
 wire \reg_module/_03073_ ;
 wire \reg_module/_03074_ ;
 wire \reg_module/_03075_ ;
 wire \reg_module/_03076_ ;
 wire \reg_module/_03077_ ;
 wire \reg_module/_03078_ ;
 wire \reg_module/_03079_ ;
 wire \reg_module/_03080_ ;
 wire \reg_module/_03081_ ;
 wire \reg_module/_03082_ ;
 wire \reg_module/_03083_ ;
 wire \reg_module/_03084_ ;
 wire \reg_module/_03085_ ;
 wire \reg_module/_03086_ ;
 wire \reg_module/_03087_ ;
 wire \reg_module/_03088_ ;
 wire \reg_module/_03089_ ;
 wire \reg_module/_03090_ ;
 wire \reg_module/_03091_ ;
 wire \reg_module/_03092_ ;
 wire \reg_module/_03093_ ;
 wire \reg_module/_03094_ ;
 wire \reg_module/_03095_ ;
 wire \reg_module/_03096_ ;
 wire \reg_module/_03097_ ;
 wire \reg_module/_03098_ ;
 wire \reg_module/_03099_ ;
 wire \reg_module/_03100_ ;
 wire \reg_module/_03101_ ;
 wire \reg_module/_03102_ ;
 wire \reg_module/_03103_ ;
 wire \reg_module/_03104_ ;
 wire \reg_module/_03105_ ;
 wire \reg_module/_03106_ ;
 wire \reg_module/_03107_ ;
 wire \reg_module/_03108_ ;
 wire \reg_module/_03109_ ;
 wire \reg_module/_03110_ ;
 wire \reg_module/_03111_ ;
 wire \reg_module/_03112_ ;
 wire \reg_module/_03113_ ;
 wire \reg_module/_03114_ ;
 wire \reg_module/_03115_ ;
 wire \reg_module/_03116_ ;
 wire \reg_module/_03117_ ;
 wire \reg_module/_03118_ ;
 wire \reg_module/_03119_ ;
 wire \reg_module/_03120_ ;
 wire \reg_module/_03121_ ;
 wire \reg_module/_03122_ ;
 wire \reg_module/_03123_ ;
 wire \reg_module/_03124_ ;
 wire \reg_module/_03125_ ;
 wire \reg_module/_03126_ ;
 wire \reg_module/_03127_ ;
 wire \reg_module/_03128_ ;
 wire \reg_module/_03129_ ;
 wire \reg_module/_03130_ ;
 wire \reg_module/_03131_ ;
 wire \reg_module/_03132_ ;
 wire \reg_module/_03133_ ;
 wire \reg_module/_03134_ ;
 wire \reg_module/_03135_ ;
 wire \reg_module/_03136_ ;
 wire \reg_module/_03137_ ;
 wire \reg_module/_03138_ ;
 wire \reg_module/_03139_ ;
 wire \reg_module/_03140_ ;
 wire \reg_module/_03141_ ;
 wire \reg_module/_03142_ ;
 wire \reg_module/_03143_ ;
 wire \reg_module/_03144_ ;
 wire \reg_module/_03145_ ;
 wire \reg_module/_03146_ ;
 wire \reg_module/_03147_ ;
 wire \reg_module/_03148_ ;
 wire \reg_module/_03149_ ;
 wire \reg_module/_03150_ ;
 wire \reg_module/_03151_ ;
 wire \reg_module/_03152_ ;
 wire \reg_module/_03153_ ;
 wire \reg_module/_03154_ ;
 wire \reg_module/_03155_ ;
 wire \reg_module/_03156_ ;
 wire \reg_module/_03157_ ;
 wire \reg_module/_03158_ ;
 wire \reg_module/_03159_ ;
 wire \reg_module/_03160_ ;
 wire \reg_module/_03161_ ;
 wire \reg_module/_03162_ ;
 wire \reg_module/_03163_ ;
 wire \reg_module/_03164_ ;
 wire \reg_module/_03165_ ;
 wire \reg_module/_03166_ ;
 wire \reg_module/_03167_ ;
 wire \reg_module/_03168_ ;
 wire \reg_module/_03169_ ;
 wire \reg_module/_03170_ ;
 wire \reg_module/_03171_ ;
 wire \reg_module/_03172_ ;
 wire \reg_module/_03173_ ;
 wire \reg_module/_03174_ ;
 wire \reg_module/_03175_ ;
 wire \reg_module/_03176_ ;
 wire \reg_module/_03177_ ;
 wire \reg_module/_03178_ ;
 wire \reg_module/_03179_ ;
 wire \reg_module/_03180_ ;
 wire \reg_module/_03181_ ;
 wire \reg_module/_03182_ ;
 wire \reg_module/_03183_ ;
 wire \reg_module/_03184_ ;
 wire \reg_module/_03185_ ;
 wire \reg_module/_03186_ ;
 wire \reg_module/_03187_ ;
 wire \reg_module/_03188_ ;
 wire \reg_module/_03189_ ;
 wire \reg_module/_03190_ ;
 wire \reg_module/_03191_ ;
 wire \reg_module/_03192_ ;
 wire \reg_module/_03193_ ;
 wire \reg_module/_03194_ ;
 wire \reg_module/_03195_ ;
 wire \reg_module/_03196_ ;
 wire \reg_module/_03197_ ;
 wire \reg_module/_03198_ ;
 wire \reg_module/_03199_ ;
 wire \reg_module/_03200_ ;
 wire \reg_module/_03201_ ;
 wire \reg_module/_03202_ ;
 wire \reg_module/_03203_ ;
 wire \reg_module/_03204_ ;
 wire \reg_module/_03205_ ;
 wire \reg_module/_03206_ ;
 wire \reg_module/_03207_ ;
 wire \reg_module/_03208_ ;
 wire \reg_module/_03209_ ;
 wire \reg_module/_03210_ ;
 wire \reg_module/_03211_ ;
 wire \reg_module/_03212_ ;
 wire \reg_module/_03213_ ;
 wire \reg_module/_03214_ ;
 wire \reg_module/_03215_ ;
 wire \reg_module/_03216_ ;
 wire \reg_module/_03217_ ;
 wire \reg_module/_03218_ ;
 wire \reg_module/_03219_ ;
 wire \reg_module/_03220_ ;
 wire \reg_module/_03221_ ;
 wire \reg_module/_03222_ ;
 wire \reg_module/_03223_ ;
 wire \reg_module/_03224_ ;
 wire \reg_module/_03225_ ;
 wire \reg_module/_03226_ ;
 wire \reg_module/_03227_ ;
 wire \reg_module/_03228_ ;
 wire \reg_module/_03229_ ;
 wire \reg_module/_03230_ ;
 wire \reg_module/_03231_ ;
 wire \reg_module/_03232_ ;
 wire \reg_module/_03233_ ;
 wire \reg_module/_03234_ ;
 wire \reg_module/_03235_ ;
 wire \reg_module/_03236_ ;
 wire \reg_module/_03237_ ;
 wire \reg_module/_03238_ ;
 wire \reg_module/_03239_ ;
 wire \reg_module/_03240_ ;
 wire \reg_module/_03241_ ;
 wire \reg_module/_03242_ ;
 wire \reg_module/_03243_ ;
 wire \reg_module/_03244_ ;
 wire \reg_module/_03245_ ;
 wire \reg_module/_03246_ ;
 wire \reg_module/_03247_ ;
 wire \reg_module/_03248_ ;
 wire \reg_module/_03249_ ;
 wire \reg_module/_03250_ ;
 wire \reg_module/_03251_ ;
 wire \reg_module/_03252_ ;
 wire \reg_module/_03253_ ;
 wire \reg_module/_03254_ ;
 wire \reg_module/_03255_ ;
 wire \reg_module/_03256_ ;
 wire \reg_module/_03257_ ;
 wire \reg_module/_03258_ ;
 wire \reg_module/_03259_ ;
 wire \reg_module/_03260_ ;
 wire \reg_module/_03261_ ;
 wire \reg_module/_03262_ ;
 wire \reg_module/_03263_ ;
 wire \reg_module/_03264_ ;
 wire \reg_module/_03265_ ;
 wire \reg_module/_03266_ ;
 wire \reg_module/_03267_ ;
 wire \reg_module/_03268_ ;
 wire \reg_module/_03269_ ;
 wire \reg_module/_03270_ ;
 wire \reg_module/_03271_ ;
 wire \reg_module/_03272_ ;
 wire \reg_module/_03273_ ;
 wire \reg_module/_03274_ ;
 wire \reg_module/_03275_ ;
 wire \reg_module/_03276_ ;
 wire \reg_module/_03277_ ;
 wire \reg_module/_03278_ ;
 wire \reg_module/_03279_ ;
 wire \reg_module/_03280_ ;
 wire \reg_module/_03281_ ;
 wire \reg_module/_03282_ ;
 wire \reg_module/_03283_ ;
 wire \reg_module/_03284_ ;
 wire \reg_module/_03285_ ;
 wire \reg_module/_03286_ ;
 wire \reg_module/_03287_ ;
 wire \reg_module/_03288_ ;
 wire \reg_module/_03289_ ;
 wire \reg_module/_03290_ ;
 wire \reg_module/_03291_ ;
 wire \reg_module/_03292_ ;
 wire \reg_module/_03293_ ;
 wire \reg_module/_03294_ ;
 wire \reg_module/_03295_ ;
 wire \reg_module/_03296_ ;
 wire \reg_module/_03297_ ;
 wire \reg_module/_03298_ ;
 wire \reg_module/_03299_ ;
 wire \reg_module/_03300_ ;
 wire \reg_module/_03301_ ;
 wire \reg_module/_03302_ ;
 wire \reg_module/_03303_ ;
 wire \reg_module/_03304_ ;
 wire \reg_module/_03305_ ;
 wire \reg_module/_03306_ ;
 wire \reg_module/_03307_ ;
 wire \reg_module/_03308_ ;
 wire \reg_module/_03309_ ;
 wire \reg_module/_03310_ ;
 wire \reg_module/_03311_ ;
 wire \reg_module/_03312_ ;
 wire \reg_module/_03313_ ;
 wire \reg_module/_03314_ ;
 wire \reg_module/_03315_ ;
 wire \reg_module/_03316_ ;
 wire \reg_module/_03317_ ;
 wire \reg_module/_03318_ ;
 wire \reg_module/_03319_ ;
 wire \reg_module/_03320_ ;
 wire \reg_module/_03321_ ;
 wire \reg_module/_03322_ ;
 wire \reg_module/_03323_ ;
 wire \reg_module/_03324_ ;
 wire \reg_module/_03325_ ;
 wire \reg_module/_03326_ ;
 wire \reg_module/_03327_ ;
 wire \reg_module/_03328_ ;
 wire \reg_module/_03329_ ;
 wire \reg_module/_03330_ ;
 wire \reg_module/_03331_ ;
 wire \reg_module/_03332_ ;
 wire \reg_module/_03333_ ;
 wire \reg_module/_03334_ ;
 wire \reg_module/_03335_ ;
 wire \reg_module/_03336_ ;
 wire \reg_module/_03337_ ;
 wire \reg_module/_03338_ ;
 wire \reg_module/_03339_ ;
 wire \reg_module/_03340_ ;
 wire \reg_module/_03341_ ;
 wire \reg_module/_03342_ ;
 wire \reg_module/_03343_ ;
 wire \reg_module/_03344_ ;
 wire \reg_module/_03345_ ;
 wire \reg_module/_03346_ ;
 wire \reg_module/_03347_ ;
 wire \reg_module/_03348_ ;
 wire \reg_module/_03349_ ;
 wire \reg_module/_03350_ ;
 wire \reg_module/_03351_ ;
 wire \reg_module/_03352_ ;
 wire \reg_module/_03353_ ;
 wire \reg_module/_03354_ ;
 wire \reg_module/_03355_ ;
 wire \reg_module/_03356_ ;
 wire \reg_module/_03357_ ;
 wire \reg_module/_03358_ ;
 wire \reg_module/_03359_ ;
 wire \reg_module/_03360_ ;
 wire \reg_module/_03361_ ;
 wire \reg_module/_03362_ ;
 wire \reg_module/_03363_ ;
 wire \reg_module/_03364_ ;
 wire \reg_module/_03365_ ;
 wire \reg_module/_03366_ ;
 wire \reg_module/_03367_ ;
 wire \reg_module/_03368_ ;
 wire \reg_module/_03369_ ;
 wire \reg_module/_03370_ ;
 wire \reg_module/_03371_ ;
 wire \reg_module/_03372_ ;
 wire \reg_module/_03373_ ;
 wire \reg_module/_03374_ ;
 wire \reg_module/_03375_ ;
 wire \reg_module/_03376_ ;
 wire \reg_module/_03377_ ;
 wire \reg_module/_03378_ ;
 wire \reg_module/_03379_ ;
 wire \reg_module/_03380_ ;
 wire \reg_module/_03381_ ;
 wire \reg_module/_03382_ ;
 wire \reg_module/_03383_ ;
 wire \reg_module/_03384_ ;
 wire \reg_module/_03385_ ;
 wire \reg_module/_03386_ ;
 wire \reg_module/_03387_ ;
 wire \reg_module/_03388_ ;
 wire \reg_module/_03389_ ;
 wire \reg_module/_03390_ ;
 wire \reg_module/_03391_ ;
 wire \reg_module/_03392_ ;
 wire \reg_module/_03393_ ;
 wire \reg_module/_03394_ ;
 wire \reg_module/_03395_ ;
 wire \reg_module/_03396_ ;
 wire \reg_module/_03397_ ;
 wire \reg_module/_03398_ ;
 wire \reg_module/_03399_ ;
 wire \reg_module/_03400_ ;
 wire \reg_module/_03401_ ;
 wire \reg_module/_03402_ ;
 wire \reg_module/_03403_ ;
 wire \reg_module/_03404_ ;
 wire \reg_module/_03405_ ;
 wire \reg_module/_03406_ ;
 wire \reg_module/_03407_ ;
 wire \reg_module/_03408_ ;
 wire \reg_module/_03409_ ;
 wire \reg_module/_03410_ ;
 wire \reg_module/_03411_ ;
 wire \reg_module/_03412_ ;
 wire \reg_module/_03413_ ;
 wire \reg_module/_03414_ ;
 wire \reg_module/_03415_ ;
 wire \reg_module/_03416_ ;
 wire \reg_module/_03417_ ;
 wire \reg_module/_03418_ ;
 wire \reg_module/_03419_ ;
 wire \reg_module/_03420_ ;
 wire \reg_module/_03421_ ;
 wire \reg_module/_03422_ ;
 wire \reg_module/_03423_ ;
 wire \reg_module/_03424_ ;
 wire \reg_module/_03425_ ;
 wire \reg_module/_03426_ ;
 wire \reg_module/_03427_ ;
 wire \reg_module/_03428_ ;
 wire \reg_module/_03429_ ;
 wire \reg_module/_03430_ ;
 wire \reg_module/_03431_ ;
 wire \reg_module/_03432_ ;
 wire \reg_module/_03433_ ;
 wire \reg_module/_03434_ ;
 wire \reg_module/_03435_ ;
 wire \reg_module/_03436_ ;
 wire \reg_module/_03437_ ;
 wire \reg_module/_03438_ ;
 wire \reg_module/_03439_ ;
 wire \reg_module/_03440_ ;
 wire \reg_module/_03441_ ;
 wire \reg_module/_03442_ ;
 wire \reg_module/_03443_ ;
 wire \reg_module/_03444_ ;
 wire \reg_module/_03445_ ;
 wire \reg_module/_03446_ ;
 wire \reg_module/_03447_ ;
 wire \reg_module/_03448_ ;
 wire \reg_module/_03449_ ;
 wire \reg_module/_03450_ ;
 wire \reg_module/_03451_ ;
 wire \reg_module/_03452_ ;
 wire \reg_module/_03453_ ;
 wire \reg_module/_03454_ ;
 wire \reg_module/_03455_ ;
 wire \reg_module/_03456_ ;
 wire \reg_module/_03457_ ;
 wire \reg_module/_03458_ ;
 wire \reg_module/_03459_ ;
 wire \reg_module/_03460_ ;
 wire \reg_module/_03461_ ;
 wire \reg_module/_03462_ ;
 wire \reg_module/_03463_ ;
 wire \reg_module/_03464_ ;
 wire \reg_module/_03465_ ;
 wire \reg_module/_03466_ ;
 wire \reg_module/_03467_ ;
 wire \reg_module/_03468_ ;
 wire \reg_module/_03469_ ;
 wire \reg_module/_03470_ ;
 wire \reg_module/_03471_ ;
 wire \reg_module/_03472_ ;
 wire \reg_module/_03473_ ;
 wire \reg_module/_03474_ ;
 wire \reg_module/_03475_ ;
 wire \reg_module/_03476_ ;
 wire \reg_module/_03477_ ;
 wire \reg_module/_03478_ ;
 wire \reg_module/_03479_ ;
 wire \reg_module/_03480_ ;
 wire \reg_module/_03481_ ;
 wire \reg_module/_03482_ ;
 wire \reg_module/_03483_ ;
 wire \reg_module/_03484_ ;
 wire \reg_module/_03485_ ;
 wire \reg_module/_03486_ ;
 wire \reg_module/_03487_ ;
 wire \reg_module/_03488_ ;
 wire \reg_module/_03489_ ;
 wire \reg_module/_03490_ ;
 wire \reg_module/_03491_ ;
 wire \reg_module/_03492_ ;
 wire \reg_module/_03493_ ;
 wire \reg_module/_03494_ ;
 wire \reg_module/_03495_ ;
 wire \reg_module/_03496_ ;
 wire \reg_module/_03497_ ;
 wire \reg_module/_03498_ ;
 wire \reg_module/_03499_ ;
 wire \reg_module/_03500_ ;
 wire \reg_module/_03501_ ;
 wire \reg_module/_03502_ ;
 wire \reg_module/_03503_ ;
 wire \reg_module/_03504_ ;
 wire \reg_module/_03505_ ;
 wire \reg_module/_03506_ ;
 wire \reg_module/_03507_ ;
 wire \reg_module/_03508_ ;
 wire \reg_module/_03509_ ;
 wire \reg_module/_03510_ ;
 wire \reg_module/_03511_ ;
 wire \reg_module/_03512_ ;
 wire \reg_module/_03513_ ;
 wire \reg_module/_03514_ ;
 wire \reg_module/_03515_ ;
 wire \reg_module/_03516_ ;
 wire \reg_module/_03517_ ;
 wire \reg_module/_03518_ ;
 wire \reg_module/_03519_ ;
 wire \reg_module/_03520_ ;
 wire \reg_module/_03521_ ;
 wire \reg_module/_03522_ ;
 wire \reg_module/_03523_ ;
 wire \reg_module/_03524_ ;
 wire \reg_module/_03525_ ;
 wire \reg_module/_03526_ ;
 wire \reg_module/_03527_ ;
 wire \reg_module/_03528_ ;
 wire \reg_module/_03529_ ;
 wire \reg_module/_03530_ ;
 wire \reg_module/_03531_ ;
 wire \reg_module/_03532_ ;
 wire \reg_module/_03533_ ;
 wire \reg_module/_03534_ ;
 wire \reg_module/_03535_ ;
 wire \reg_module/_03536_ ;
 wire \reg_module/_03537_ ;
 wire \reg_module/_03538_ ;
 wire \reg_module/_03539_ ;
 wire \reg_module/_03540_ ;
 wire \reg_module/_03541_ ;
 wire \reg_module/_03542_ ;
 wire \reg_module/_03543_ ;
 wire \reg_module/_03544_ ;
 wire \reg_module/_03545_ ;
 wire \reg_module/_03546_ ;
 wire \reg_module/_03547_ ;
 wire \reg_module/_03548_ ;
 wire \reg_module/_03549_ ;
 wire \reg_module/_03550_ ;
 wire \reg_module/_03551_ ;
 wire \reg_module/_03552_ ;
 wire \reg_module/_03553_ ;
 wire \reg_module/_03554_ ;
 wire \reg_module/_03555_ ;
 wire \reg_module/_03556_ ;
 wire \reg_module/_03557_ ;
 wire \reg_module/_03558_ ;
 wire \reg_module/_03559_ ;
 wire \reg_module/_03560_ ;
 wire \reg_module/_03561_ ;
 wire \reg_module/_03562_ ;
 wire \reg_module/_03563_ ;
 wire \reg_module/_03564_ ;
 wire \reg_module/_03565_ ;
 wire \reg_module/_03566_ ;
 wire \reg_module/_03567_ ;
 wire \reg_module/_03568_ ;
 wire \reg_module/_03569_ ;
 wire \reg_module/_03570_ ;
 wire \reg_module/_03571_ ;
 wire \reg_module/_03572_ ;
 wire \reg_module/_03573_ ;
 wire \reg_module/_03574_ ;
 wire \reg_module/_03575_ ;
 wire \reg_module/_03576_ ;
 wire \reg_module/_03577_ ;
 wire \reg_module/_03578_ ;
 wire \reg_module/_03579_ ;
 wire \reg_module/_03580_ ;
 wire \reg_module/_03581_ ;
 wire \reg_module/_03582_ ;
 wire \reg_module/_03583_ ;
 wire \reg_module/_03584_ ;
 wire \reg_module/_03585_ ;
 wire \reg_module/_03586_ ;
 wire \reg_module/_03587_ ;
 wire \reg_module/_03588_ ;
 wire \reg_module/_03589_ ;
 wire \reg_module/_03590_ ;
 wire \reg_module/_03591_ ;
 wire \reg_module/_03592_ ;
 wire \reg_module/_03593_ ;
 wire \reg_module/_03594_ ;
 wire \reg_module/_03595_ ;
 wire \reg_module/_03596_ ;
 wire \reg_module/_03597_ ;
 wire \reg_module/_03598_ ;
 wire \reg_module/_03599_ ;
 wire \reg_module/_03600_ ;
 wire \reg_module/_03601_ ;
 wire \reg_module/_03602_ ;
 wire \reg_module/_03603_ ;
 wire \reg_module/_03604_ ;
 wire \reg_module/_03605_ ;
 wire \reg_module/_03606_ ;
 wire \reg_module/_03607_ ;
 wire \reg_module/_03608_ ;
 wire \reg_module/_03609_ ;
 wire \reg_module/_03610_ ;
 wire \reg_module/_03611_ ;
 wire \reg_module/_03612_ ;
 wire \reg_module/_03613_ ;
 wire \reg_module/_03614_ ;
 wire \reg_module/_03615_ ;
 wire \reg_module/_03616_ ;
 wire \reg_module/_03617_ ;
 wire \reg_module/_03618_ ;
 wire \reg_module/_03619_ ;
 wire \reg_module/_03620_ ;
 wire \reg_module/_03621_ ;
 wire \reg_module/_03622_ ;
 wire \reg_module/_03623_ ;
 wire \reg_module/_03624_ ;
 wire \reg_module/_03625_ ;
 wire \reg_module/_03626_ ;
 wire \reg_module/_03627_ ;
 wire \reg_module/_03628_ ;
 wire \reg_module/_03629_ ;
 wire \reg_module/_03630_ ;
 wire \reg_module/_03631_ ;
 wire \reg_module/_03632_ ;
 wire \reg_module/_03633_ ;
 wire \reg_module/_03634_ ;
 wire \reg_module/_03635_ ;
 wire \reg_module/_03636_ ;
 wire \reg_module/_03637_ ;
 wire \reg_module/_03638_ ;
 wire \reg_module/_03639_ ;
 wire \reg_module/_03640_ ;
 wire \reg_module/_03641_ ;
 wire \reg_module/_03642_ ;
 wire \reg_module/_03643_ ;
 wire \reg_module/_03644_ ;
 wire \reg_module/_03645_ ;
 wire \reg_module/_03646_ ;
 wire \reg_module/_03647_ ;
 wire \reg_module/_03648_ ;
 wire \reg_module/_03649_ ;
 wire \reg_module/_03650_ ;
 wire \reg_module/_03651_ ;
 wire \reg_module/_03652_ ;
 wire \reg_module/_03653_ ;
 wire \reg_module/_03654_ ;
 wire \reg_module/_03655_ ;
 wire \reg_module/_03656_ ;
 wire \reg_module/_03657_ ;
 wire \reg_module/_03658_ ;
 wire \reg_module/_03659_ ;
 wire \reg_module/_03660_ ;
 wire \reg_module/_03661_ ;
 wire \reg_module/_03662_ ;
 wire \reg_module/_03663_ ;
 wire \reg_module/_03664_ ;
 wire \reg_module/_03665_ ;
 wire \reg_module/_03666_ ;
 wire \reg_module/_03667_ ;
 wire \reg_module/_03668_ ;
 wire \reg_module/_03669_ ;
 wire \reg_module/_03670_ ;
 wire \reg_module/_03671_ ;
 wire \reg_module/_03672_ ;
 wire \reg_module/_03673_ ;
 wire \reg_module/_03674_ ;
 wire \reg_module/_03675_ ;
 wire \reg_module/_03676_ ;
 wire \reg_module/_03677_ ;
 wire \reg_module/_03678_ ;
 wire \reg_module/_03679_ ;
 wire \reg_module/_03680_ ;
 wire \reg_module/_03681_ ;
 wire \reg_module/_03682_ ;
 wire \reg_module/_03683_ ;
 wire \reg_module/_03684_ ;
 wire \reg_module/_03685_ ;
 wire \reg_module/_03686_ ;
 wire \reg_module/_03687_ ;
 wire \reg_module/_03688_ ;
 wire \reg_module/_03689_ ;
 wire \reg_module/_03690_ ;
 wire \reg_module/_03691_ ;
 wire \reg_module/_03692_ ;
 wire \reg_module/_03693_ ;
 wire \reg_module/_03694_ ;
 wire \reg_module/_03695_ ;
 wire \reg_module/_03696_ ;
 wire \reg_module/_03697_ ;
 wire \reg_module/_03698_ ;
 wire \reg_module/_03699_ ;
 wire \reg_module/_03700_ ;
 wire \reg_module/_03701_ ;
 wire \reg_module/_03702_ ;
 wire \reg_module/_03703_ ;
 wire \reg_module/_03704_ ;
 wire \reg_module/_03705_ ;
 wire \reg_module/_03706_ ;
 wire \reg_module/_03707_ ;
 wire \reg_module/_03708_ ;
 wire \reg_module/_03709_ ;
 wire \reg_module/_03710_ ;
 wire \reg_module/_03711_ ;
 wire \reg_module/_03712_ ;
 wire \reg_module/_03713_ ;
 wire \reg_module/_03714_ ;
 wire \reg_module/_03715_ ;
 wire \reg_module/_03716_ ;
 wire \reg_module/_03717_ ;
 wire \reg_module/_03718_ ;
 wire \reg_module/_03719_ ;
 wire \reg_module/_03720_ ;
 wire \reg_module/_03721_ ;
 wire \reg_module/_03722_ ;
 wire \reg_module/_03723_ ;
 wire \reg_module/_03724_ ;
 wire \reg_module/_03725_ ;
 wire \reg_module/_03726_ ;
 wire \reg_module/_03727_ ;
 wire \reg_module/_03728_ ;
 wire \reg_module/_03729_ ;
 wire \reg_module/_03730_ ;
 wire \reg_module/_03731_ ;
 wire \reg_module/_03732_ ;
 wire \reg_module/_03733_ ;
 wire \reg_module/_03734_ ;
 wire \reg_module/_03735_ ;
 wire \reg_module/_03736_ ;
 wire \reg_module/_03737_ ;
 wire \reg_module/_03738_ ;
 wire \reg_module/_03739_ ;
 wire \reg_module/_03740_ ;
 wire \reg_module/_03741_ ;
 wire \reg_module/_03742_ ;
 wire \reg_module/_03743_ ;
 wire \reg_module/_03744_ ;
 wire \reg_module/_03745_ ;
 wire \reg_module/_03746_ ;
 wire \reg_module/_03747_ ;
 wire \reg_module/_03748_ ;
 wire \reg_module/_03749_ ;
 wire \reg_module/_03750_ ;
 wire \reg_module/_03751_ ;
 wire \reg_module/_03752_ ;
 wire \reg_module/_03753_ ;
 wire \reg_module/_03754_ ;
 wire \reg_module/_03755_ ;
 wire \reg_module/_03756_ ;
 wire \reg_module/_03757_ ;
 wire \reg_module/_03758_ ;
 wire \reg_module/_03759_ ;
 wire \reg_module/_03760_ ;
 wire \reg_module/_03761_ ;
 wire \reg_module/_03762_ ;
 wire \reg_module/_03763_ ;
 wire \reg_module/_03764_ ;
 wire \reg_module/_03765_ ;
 wire \reg_module/_03766_ ;
 wire \reg_module/_03767_ ;
 wire \reg_module/_03768_ ;
 wire \reg_module/_03769_ ;
 wire \reg_module/_03770_ ;
 wire \reg_module/_03771_ ;
 wire \reg_module/_03772_ ;
 wire \reg_module/_03773_ ;
 wire \reg_module/_03774_ ;
 wire \reg_module/_03775_ ;
 wire \reg_module/_03776_ ;
 wire \reg_module/_03777_ ;
 wire \reg_module/_03778_ ;
 wire \reg_module/_03779_ ;
 wire \reg_module/_03780_ ;
 wire \reg_module/_03781_ ;
 wire \reg_module/_03782_ ;
 wire \reg_module/_03783_ ;
 wire \reg_module/_03784_ ;
 wire \reg_module/_03785_ ;
 wire \reg_module/_03786_ ;
 wire \reg_module/_03787_ ;
 wire \reg_module/_03788_ ;
 wire \reg_module/_03789_ ;
 wire \reg_module/_03790_ ;
 wire \reg_module/_03791_ ;
 wire \reg_module/_03792_ ;
 wire \reg_module/_03793_ ;
 wire \reg_module/_03794_ ;
 wire \reg_module/_03795_ ;
 wire \reg_module/_03796_ ;
 wire \reg_module/_03797_ ;
 wire \reg_module/_03798_ ;
 wire \reg_module/_03799_ ;
 wire \reg_module/_03800_ ;
 wire \reg_module/_03801_ ;
 wire \reg_module/_03802_ ;
 wire \reg_module/_03803_ ;
 wire \reg_module/_03804_ ;
 wire \reg_module/_03805_ ;
 wire \reg_module/_03806_ ;
 wire \reg_module/_03807_ ;
 wire \reg_module/_03808_ ;
 wire \reg_module/_03809_ ;
 wire \reg_module/_03810_ ;
 wire \reg_module/_03811_ ;
 wire \reg_module/_03812_ ;
 wire \reg_module/_03813_ ;
 wire \reg_module/_03814_ ;
 wire \reg_module/_03815_ ;
 wire \reg_module/_03816_ ;
 wire \reg_module/_03817_ ;
 wire \reg_module/_03818_ ;
 wire \reg_module/_03819_ ;
 wire \reg_module/_03820_ ;
 wire \reg_module/_03821_ ;
 wire \reg_module/_03822_ ;
 wire \reg_module/_03823_ ;
 wire \reg_module/_03824_ ;
 wire \reg_module/_03825_ ;
 wire \reg_module/_03826_ ;
 wire \reg_module/_03827_ ;
 wire \reg_module/_03828_ ;
 wire \reg_module/_03829_ ;
 wire \reg_module/_03830_ ;
 wire \reg_module/_03831_ ;
 wire \reg_module/_03832_ ;
 wire \reg_module/_03833_ ;
 wire \reg_module/_03834_ ;
 wire \reg_module/_03835_ ;
 wire \reg_module/_03836_ ;
 wire \reg_module/_03837_ ;
 wire \reg_module/_03838_ ;
 wire \reg_module/_03839_ ;
 wire \reg_module/_03840_ ;
 wire \reg_module/_03841_ ;
 wire \reg_module/_03842_ ;
 wire \reg_module/_03843_ ;
 wire \reg_module/_03844_ ;
 wire \reg_module/_03845_ ;
 wire \reg_module/_03846_ ;
 wire \reg_module/_03847_ ;
 wire \reg_module/_03848_ ;
 wire \reg_module/_03849_ ;
 wire \reg_module/_03850_ ;
 wire \reg_module/_03851_ ;
 wire \reg_module/_03852_ ;
 wire \reg_module/_03853_ ;
 wire \reg_module/_03854_ ;
 wire \reg_module/_03855_ ;
 wire \reg_module/_03856_ ;
 wire \reg_module/_03857_ ;
 wire \reg_module/_03858_ ;
 wire \reg_module/_03859_ ;
 wire \reg_module/_03860_ ;
 wire \reg_module/_03861_ ;
 wire \reg_module/_03862_ ;
 wire \reg_module/_03863_ ;
 wire \reg_module/_03864_ ;
 wire \reg_module/_03865_ ;
 wire \reg_module/_03866_ ;
 wire \reg_module/_03867_ ;
 wire \reg_module/_03868_ ;
 wire \reg_module/_03869_ ;
 wire \reg_module/_03870_ ;
 wire \reg_module/_03871_ ;
 wire \reg_module/_03872_ ;
 wire \reg_module/_03873_ ;
 wire \reg_module/_03874_ ;
 wire \reg_module/_03875_ ;
 wire \reg_module/_03876_ ;
 wire \reg_module/_03877_ ;
 wire \reg_module/_03878_ ;
 wire \reg_module/_03879_ ;
 wire \reg_module/_03880_ ;
 wire \reg_module/_03881_ ;
 wire \reg_module/_03882_ ;
 wire \reg_module/_03883_ ;
 wire \reg_module/_03884_ ;
 wire \reg_module/_03885_ ;
 wire \reg_module/_03886_ ;
 wire \reg_module/_03887_ ;
 wire \reg_module/_03888_ ;
 wire \reg_module/_03889_ ;
 wire \reg_module/_03890_ ;
 wire \reg_module/_03891_ ;
 wire \reg_module/_03892_ ;
 wire \reg_module/_03893_ ;
 wire \reg_module/_03894_ ;
 wire \reg_module/_03895_ ;
 wire \reg_module/_03896_ ;
 wire \reg_module/_03897_ ;
 wire \reg_module/_03898_ ;
 wire \reg_module/_03899_ ;
 wire \reg_module/_03900_ ;
 wire \reg_module/_03901_ ;
 wire \reg_module/_03902_ ;
 wire \reg_module/_03903_ ;
 wire \reg_module/_03904_ ;
 wire \reg_module/_03905_ ;
 wire \reg_module/_03906_ ;
 wire \reg_module/_03907_ ;
 wire \reg_module/_03908_ ;
 wire \reg_module/_03909_ ;
 wire \reg_module/_03910_ ;
 wire \reg_module/_03911_ ;
 wire \reg_module/_03912_ ;
 wire \reg_module/_03913_ ;
 wire \reg_module/_03914_ ;
 wire \reg_module/_03915_ ;
 wire \reg_module/_03916_ ;
 wire \reg_module/_03917_ ;
 wire \reg_module/_03918_ ;
 wire \reg_module/_03919_ ;
 wire \reg_module/_03920_ ;
 wire \reg_module/_03921_ ;
 wire \reg_module/_03922_ ;
 wire \reg_module/_03923_ ;
 wire \reg_module/_03924_ ;
 wire \reg_module/_03925_ ;
 wire \reg_module/_03926_ ;
 wire \reg_module/_03927_ ;
 wire \reg_module/_03928_ ;
 wire \reg_module/_03929_ ;
 wire \reg_module/_03930_ ;
 wire \reg_module/_03931_ ;
 wire \reg_module/_03932_ ;
 wire \reg_module/_03933_ ;
 wire \reg_module/_03934_ ;
 wire \reg_module/_03935_ ;
 wire \reg_module/_03936_ ;
 wire \reg_module/_03937_ ;
 wire \reg_module/_03938_ ;
 wire \reg_module/_03939_ ;
 wire \reg_module/_03940_ ;
 wire \reg_module/_03941_ ;
 wire \reg_module/_03942_ ;
 wire \reg_module/_03943_ ;
 wire \reg_module/_03944_ ;
 wire \reg_module/_03945_ ;
 wire \reg_module/_03946_ ;
 wire \reg_module/_03947_ ;
 wire \reg_module/_03948_ ;
 wire \reg_module/_03949_ ;
 wire \reg_module/_03950_ ;
 wire \reg_module/_03951_ ;
 wire \reg_module/_03952_ ;
 wire \reg_module/_03953_ ;
 wire \reg_module/_03954_ ;
 wire \reg_module/_03955_ ;
 wire \reg_module/_03956_ ;
 wire \reg_module/_03957_ ;
 wire \reg_module/_03958_ ;
 wire \reg_module/_03959_ ;
 wire \reg_module/_03960_ ;
 wire \reg_module/_03961_ ;
 wire \reg_module/_03962_ ;
 wire \reg_module/_03963_ ;
 wire \reg_module/_03964_ ;
 wire \reg_module/_03965_ ;
 wire \reg_module/_03966_ ;
 wire \reg_module/_03967_ ;
 wire \reg_module/_03968_ ;
 wire \reg_module/_03969_ ;
 wire \reg_module/_03970_ ;
 wire \reg_module/_03971_ ;
 wire \reg_module/_03972_ ;
 wire \reg_module/_03973_ ;
 wire \reg_module/_03974_ ;
 wire \reg_module/_03975_ ;
 wire \reg_module/_03976_ ;
 wire \reg_module/_03977_ ;
 wire \reg_module/_03978_ ;
 wire \reg_module/_03979_ ;
 wire \reg_module/_03980_ ;
 wire \reg_module/_03981_ ;
 wire \reg_module/_03982_ ;
 wire \reg_module/_03983_ ;
 wire \reg_module/_03984_ ;
 wire \reg_module/_03985_ ;
 wire \reg_module/_03986_ ;
 wire \reg_module/_03987_ ;
 wire \reg_module/_03988_ ;
 wire \reg_module/_03989_ ;
 wire \reg_module/_03990_ ;
 wire \reg_module/_03991_ ;
 wire \reg_module/_03992_ ;
 wire \reg_module/_03993_ ;
 wire \reg_module/_03994_ ;
 wire \reg_module/_03995_ ;
 wire \reg_module/_03996_ ;
 wire \reg_module/_03997_ ;
 wire \reg_module/_03998_ ;
 wire \reg_module/_03999_ ;
 wire \reg_module/_04000_ ;
 wire \reg_module/_04001_ ;
 wire \reg_module/_04002_ ;
 wire \reg_module/_04003_ ;
 wire \reg_module/_04004_ ;
 wire \reg_module/_04005_ ;
 wire \reg_module/_04006_ ;
 wire \reg_module/_04007_ ;
 wire \reg_module/_04008_ ;
 wire \reg_module/_04009_ ;
 wire \reg_module/_04010_ ;
 wire \reg_module/_04011_ ;
 wire \reg_module/_04012_ ;
 wire \reg_module/_04013_ ;
 wire \reg_module/_04014_ ;
 wire \reg_module/_04015_ ;
 wire \reg_module/_04016_ ;
 wire \reg_module/_04017_ ;
 wire \reg_module/_04018_ ;
 wire \reg_module/_04019_ ;
 wire \reg_module/_04020_ ;
 wire \reg_module/_04021_ ;
 wire \reg_module/_04022_ ;
 wire \reg_module/_04023_ ;
 wire \reg_module/_04024_ ;
 wire \reg_module/_04025_ ;
 wire \reg_module/_04026_ ;
 wire \reg_module/_04027_ ;
 wire \reg_module/_04028_ ;
 wire \reg_module/_04029_ ;
 wire \reg_module/_04030_ ;
 wire \reg_module/_04031_ ;
 wire \reg_module/_04032_ ;
 wire \reg_module/_04033_ ;
 wire \reg_module/_04034_ ;
 wire \reg_module/_04035_ ;
 wire \reg_module/_04036_ ;
 wire \reg_module/_04037_ ;
 wire \reg_module/_04038_ ;
 wire \reg_module/_04039_ ;
 wire \reg_module/_04040_ ;
 wire \reg_module/_04041_ ;
 wire \reg_module/_04042_ ;
 wire \reg_module/_04043_ ;
 wire \reg_module/_04044_ ;
 wire \reg_module/_04045_ ;
 wire \reg_module/_04046_ ;
 wire \reg_module/_04047_ ;
 wire \reg_module/_04048_ ;
 wire \reg_module/_04049_ ;
 wire \reg_module/_04050_ ;
 wire \reg_module/_04051_ ;
 wire \reg_module/_04052_ ;
 wire \reg_module/_04053_ ;
 wire \reg_module/_04054_ ;
 wire \reg_module/_04055_ ;
 wire \reg_module/_04056_ ;
 wire \reg_module/_04057_ ;
 wire \reg_module/_04058_ ;
 wire \reg_module/_04059_ ;
 wire \reg_module/_04060_ ;
 wire \reg_module/_04061_ ;
 wire \reg_module/_04062_ ;
 wire \reg_module/_04063_ ;
 wire \reg_module/_04064_ ;
 wire \reg_module/_04065_ ;
 wire \reg_module/_04066_ ;
 wire \reg_module/_04067_ ;
 wire \reg_module/_04068_ ;
 wire \reg_module/_04069_ ;
 wire \reg_module/_04070_ ;
 wire \reg_module/_04071_ ;
 wire \reg_module/_04072_ ;
 wire \reg_module/_04073_ ;
 wire \reg_module/_04074_ ;
 wire \reg_module/_04075_ ;
 wire \reg_module/_04076_ ;
 wire \reg_module/_04077_ ;
 wire \reg_module/_04078_ ;
 wire \reg_module/_04079_ ;
 wire \reg_module/_04080_ ;
 wire \reg_module/_04081_ ;
 wire \reg_module/_04082_ ;
 wire \reg_module/_04083_ ;
 wire \reg_module/_04084_ ;
 wire \reg_module/_04085_ ;
 wire \reg_module/_04086_ ;
 wire \reg_module/_04087_ ;
 wire \reg_module/_04088_ ;
 wire \reg_module/_04089_ ;
 wire \reg_module/_04090_ ;
 wire \reg_module/_04091_ ;
 wire \reg_module/_04092_ ;
 wire \reg_module/_04093_ ;
 wire \reg_module/_04094_ ;
 wire \reg_module/_04095_ ;
 wire \reg_module/_04096_ ;
 wire \reg_module/_04097_ ;
 wire \reg_module/_04098_ ;
 wire \reg_module/_04099_ ;
 wire \reg_module/_04100_ ;
 wire \reg_module/_04101_ ;
 wire \reg_module/_04102_ ;
 wire \reg_module/_04103_ ;
 wire \reg_module/_04104_ ;
 wire \reg_module/_04105_ ;
 wire \reg_module/_04106_ ;
 wire \reg_module/_04107_ ;
 wire \reg_module/_04108_ ;
 wire \reg_module/_04109_ ;
 wire \reg_module/_04110_ ;
 wire \reg_module/_04111_ ;
 wire \reg_module/_04112_ ;
 wire \reg_module/_04113_ ;
 wire \reg_module/_04114_ ;
 wire \reg_module/_04115_ ;
 wire \reg_module/_04116_ ;
 wire \reg_module/_04117_ ;
 wire \reg_module/_04118_ ;
 wire \reg_module/_04119_ ;
 wire \reg_module/_04120_ ;
 wire \reg_module/_04121_ ;
 wire \reg_module/_04122_ ;
 wire \reg_module/_04123_ ;
 wire \reg_module/_04124_ ;
 wire \reg_module/_04125_ ;
 wire \reg_module/_04126_ ;
 wire \reg_module/_04127_ ;
 wire \reg_module/_04128_ ;
 wire \reg_module/_04129_ ;
 wire \reg_module/_04130_ ;
 wire \reg_module/_04131_ ;
 wire \reg_module/_04132_ ;
 wire \reg_module/_04133_ ;
 wire \reg_module/_04134_ ;
 wire \reg_module/_04135_ ;
 wire \reg_module/_04136_ ;
 wire \reg_module/_04137_ ;
 wire \reg_module/_04138_ ;
 wire \reg_module/_04139_ ;
 wire \reg_module/_04140_ ;
 wire \reg_module/_04141_ ;
 wire \reg_module/_04142_ ;
 wire \reg_module/_04143_ ;
 wire \reg_module/_04144_ ;
 wire \reg_module/_04145_ ;
 wire \reg_module/_04146_ ;
 wire \reg_module/_04147_ ;
 wire \reg_module/_04148_ ;
 wire \reg_module/_04149_ ;
 wire \reg_module/_04150_ ;
 wire \reg_module/_04151_ ;
 wire \reg_module/_04152_ ;
 wire \reg_module/_04153_ ;
 wire \reg_module/_04154_ ;
 wire \reg_module/_04155_ ;
 wire \reg_module/_04156_ ;
 wire \reg_module/_04157_ ;
 wire \reg_module/_04158_ ;
 wire \reg_module/_04159_ ;
 wire \reg_module/_04160_ ;
 wire \reg_module/_04161_ ;
 wire \reg_module/_04162_ ;
 wire \reg_module/_04163_ ;
 wire \reg_module/_04164_ ;
 wire \reg_module/_04165_ ;
 wire \reg_module/_04166_ ;
 wire \reg_module/_04167_ ;
 wire \reg_module/_04168_ ;
 wire \reg_module/_04169_ ;
 wire \reg_module/_04170_ ;
 wire \reg_module/_04171_ ;
 wire \reg_module/_04172_ ;
 wire \reg_module/_04173_ ;
 wire \reg_module/_04174_ ;
 wire \reg_module/_04175_ ;
 wire \reg_module/_04176_ ;
 wire \reg_module/_04177_ ;
 wire \reg_module/_04178_ ;
 wire \reg_module/_04179_ ;
 wire \reg_module/_04180_ ;
 wire \reg_module/_04181_ ;
 wire \reg_module/_04182_ ;
 wire \reg_module/_04183_ ;
 wire \reg_module/_04184_ ;
 wire \reg_module/_04185_ ;
 wire \reg_module/_04186_ ;
 wire \reg_module/_04187_ ;
 wire \reg_module/_04188_ ;
 wire \reg_module/_04189_ ;
 wire \reg_module/_04190_ ;
 wire \reg_module/_04191_ ;
 wire \reg_module/_04192_ ;
 wire \reg_module/_04193_ ;
 wire \reg_module/_04194_ ;
 wire \reg_module/_04195_ ;
 wire \reg_module/_04196_ ;
 wire \reg_module/_04197_ ;
 wire \reg_module/_04198_ ;
 wire \reg_module/_04199_ ;
 wire \reg_module/_04200_ ;
 wire \reg_module/_04201_ ;
 wire \reg_module/_04202_ ;
 wire \reg_module/_04203_ ;
 wire \reg_module/_04204_ ;
 wire \reg_module/_04205_ ;
 wire \reg_module/_04206_ ;
 wire \reg_module/_04207_ ;
 wire \reg_module/_04208_ ;
 wire \reg_module/_04209_ ;
 wire \reg_module/_04210_ ;
 wire \reg_module/_04211_ ;
 wire \reg_module/_04212_ ;
 wire \reg_module/_04213_ ;
 wire \reg_module/_04214_ ;
 wire \reg_module/_04215_ ;
 wire \reg_module/_04216_ ;
 wire \reg_module/_04217_ ;
 wire \reg_module/_04218_ ;
 wire \reg_module/_04219_ ;
 wire \reg_module/_04220_ ;
 wire \reg_module/_04221_ ;
 wire \reg_module/_04222_ ;
 wire \reg_module/_04223_ ;
 wire \reg_module/_04224_ ;
 wire \reg_module/_04225_ ;
 wire \reg_module/_04226_ ;
 wire \reg_module/_04227_ ;
 wire \reg_module/_04228_ ;
 wire \reg_module/_04229_ ;
 wire \reg_module/_04230_ ;
 wire \reg_module/_04231_ ;
 wire \reg_module/_04232_ ;
 wire \reg_module/_04233_ ;
 wire \reg_module/_04234_ ;
 wire \reg_module/_04235_ ;
 wire \reg_module/_04236_ ;
 wire \reg_module/_04237_ ;
 wire \reg_module/_04238_ ;
 wire \reg_module/_04239_ ;
 wire \reg_module/_04240_ ;
 wire \reg_module/_04241_ ;
 wire \reg_module/_04242_ ;
 wire \reg_module/_04243_ ;
 wire \reg_module/_04244_ ;
 wire \reg_module/_04245_ ;
 wire \reg_module/_04246_ ;
 wire \reg_module/_04247_ ;
 wire \reg_module/_04248_ ;
 wire \reg_module/_04249_ ;
 wire \reg_module/_04250_ ;
 wire \reg_module/_04251_ ;
 wire \reg_module/_04252_ ;
 wire \reg_module/_04253_ ;
 wire \reg_module/_04254_ ;
 wire \reg_module/_04255_ ;
 wire \reg_module/_04256_ ;
 wire \reg_module/_04257_ ;
 wire \reg_module/_04258_ ;
 wire \reg_module/_04259_ ;
 wire \reg_module/_04260_ ;
 wire \reg_module/_04261_ ;
 wire \reg_module/_04262_ ;
 wire \reg_module/_04263_ ;
 wire \reg_module/_04264_ ;
 wire \reg_module/_04265_ ;
 wire \reg_module/_04266_ ;
 wire \reg_module/_04267_ ;
 wire \reg_module/_04268_ ;
 wire \reg_module/_04269_ ;
 wire \reg_module/_04270_ ;
 wire \reg_module/_04271_ ;
 wire \reg_module/_04272_ ;
 wire \reg_module/_04273_ ;
 wire \reg_module/_04274_ ;
 wire \reg_module/_04275_ ;
 wire \reg_module/_04276_ ;
 wire \reg_module/_04277_ ;
 wire \reg_module/_04278_ ;
 wire \reg_module/_04279_ ;
 wire \reg_module/_04280_ ;
 wire \reg_module/_04281_ ;
 wire \reg_module/_04282_ ;
 wire \reg_module/_04283_ ;
 wire \reg_module/_04284_ ;
 wire \reg_module/_04285_ ;
 wire \reg_module/_04286_ ;
 wire \reg_module/_04287_ ;
 wire \reg_module/_04288_ ;
 wire \reg_module/_04289_ ;
 wire \reg_module/_04290_ ;
 wire \reg_module/_04291_ ;
 wire \reg_module/_04292_ ;
 wire \reg_module/_04293_ ;
 wire \reg_module/_04294_ ;
 wire \reg_module/_04295_ ;
 wire \reg_module/_04296_ ;
 wire \reg_module/_04297_ ;
 wire \reg_module/_04298_ ;
 wire \reg_module/_04299_ ;
 wire \reg_module/_04300_ ;
 wire \reg_module/_04301_ ;
 wire \reg_module/_04302_ ;
 wire \reg_module/_04303_ ;
 wire \reg_module/_04304_ ;
 wire \reg_module/_04305_ ;
 wire \reg_module/_04306_ ;
 wire \reg_module/_04307_ ;
 wire \reg_module/_04308_ ;
 wire \reg_module/_04309_ ;
 wire \reg_module/_04310_ ;
 wire \reg_module/_04311_ ;
 wire \reg_module/_04312_ ;
 wire \reg_module/_04313_ ;
 wire \reg_module/_04314_ ;
 wire \reg_module/_04315_ ;
 wire \reg_module/_04316_ ;
 wire \reg_module/_04317_ ;
 wire \reg_module/_04318_ ;
 wire \reg_module/_04319_ ;
 wire \reg_module/_04320_ ;
 wire \reg_module/_04321_ ;
 wire \reg_module/_04322_ ;
 wire \reg_module/_04323_ ;
 wire \reg_module/_04324_ ;
 wire \reg_module/_04325_ ;
 wire \reg_module/_04326_ ;
 wire \reg_module/_04327_ ;
 wire \reg_module/_04328_ ;
 wire \reg_module/_04329_ ;
 wire \reg_module/_04330_ ;
 wire \reg_module/_04331_ ;
 wire \reg_module/_04332_ ;
 wire \reg_module/_04333_ ;
 wire \reg_module/_04334_ ;
 wire \reg_module/_04335_ ;
 wire \reg_module/_04336_ ;
 wire \reg_module/_04337_ ;
 wire \reg_module/_04338_ ;
 wire \reg_module/_04339_ ;
 wire \reg_module/_04340_ ;
 wire \reg_module/_04341_ ;
 wire \reg_module/_04342_ ;
 wire \reg_module/_04343_ ;
 wire \reg_module/_04344_ ;
 wire \reg_module/_04345_ ;
 wire \reg_module/_04346_ ;
 wire \reg_module/_04347_ ;
 wire \reg_module/_04348_ ;
 wire \reg_module/_04349_ ;
 wire \reg_module/_04350_ ;
 wire \reg_module/_04351_ ;
 wire \reg_module/_04352_ ;
 wire \reg_module/_04353_ ;
 wire \reg_module/_04354_ ;
 wire \reg_module/_04355_ ;
 wire \reg_module/_04356_ ;
 wire \reg_module/_04357_ ;
 wire \reg_module/_04358_ ;
 wire \reg_module/_04359_ ;
 wire \reg_module/_04360_ ;
 wire \reg_module/_04361_ ;
 wire \reg_module/_04362_ ;
 wire \reg_module/_04363_ ;
 wire \reg_module/_04364_ ;
 wire \reg_module/_04365_ ;
 wire \reg_module/_04366_ ;
 wire \reg_module/_04367_ ;
 wire \reg_module/_04368_ ;
 wire \reg_module/_04369_ ;
 wire \reg_module/_04370_ ;
 wire \reg_module/_04371_ ;
 wire \reg_module/_04372_ ;
 wire \reg_module/_04373_ ;
 wire \reg_module/_04374_ ;
 wire \reg_module/_04375_ ;
 wire \reg_module/_04376_ ;
 wire \reg_module/_04377_ ;
 wire \reg_module/_04378_ ;
 wire \reg_module/_04379_ ;
 wire \reg_module/_04380_ ;
 wire \reg_module/_04381_ ;
 wire \reg_module/_04382_ ;
 wire \reg_module/_04383_ ;
 wire \reg_module/_04384_ ;
 wire \reg_module/_04385_ ;
 wire \reg_module/_04386_ ;
 wire \reg_module/_04387_ ;
 wire \reg_module/_04388_ ;
 wire \reg_module/_04389_ ;
 wire \reg_module/_04390_ ;
 wire \reg_module/_04391_ ;
 wire \reg_module/_04392_ ;
 wire \reg_module/_04393_ ;
 wire \reg_module/_04394_ ;
 wire \reg_module/_04395_ ;
 wire \reg_module/_04396_ ;
 wire \reg_module/_04397_ ;
 wire \reg_module/_04398_ ;
 wire \reg_module/_04399_ ;
 wire \reg_module/_04400_ ;
 wire \reg_module/_04401_ ;
 wire \reg_module/_04402_ ;
 wire \reg_module/_04403_ ;
 wire \reg_module/_04404_ ;
 wire \reg_module/_04405_ ;
 wire \reg_module/_04406_ ;
 wire \reg_module/_04407_ ;
 wire \reg_module/_04408_ ;
 wire \reg_module/_04409_ ;
 wire \reg_module/_04410_ ;
 wire \reg_module/_04411_ ;
 wire \reg_module/_04412_ ;
 wire \reg_module/_04413_ ;
 wire \reg_module/_04414_ ;
 wire \reg_module/_04415_ ;
 wire \reg_module/_04416_ ;
 wire \reg_module/_04417_ ;
 wire \reg_module/_04418_ ;
 wire \reg_module/_04419_ ;
 wire \reg_module/_04420_ ;
 wire \reg_module/_04421_ ;
 wire \reg_module/_04422_ ;
 wire \reg_module/_04423_ ;
 wire \reg_module/_04424_ ;
 wire \reg_module/_04425_ ;
 wire \reg_module/_04426_ ;
 wire \reg_module/_04427_ ;
 wire \reg_module/_04428_ ;
 wire \reg_module/_04429_ ;
 wire \reg_module/_04430_ ;
 wire \reg_module/_04431_ ;
 wire \reg_module/_04432_ ;
 wire \reg_module/_04433_ ;
 wire \reg_module/_04434_ ;
 wire \reg_module/_04435_ ;
 wire \reg_module/_04436_ ;
 wire \reg_module/_04437_ ;
 wire \reg_module/_04438_ ;
 wire \reg_module/_04439_ ;
 wire \reg_module/_04440_ ;
 wire \reg_module/_04441_ ;
 wire \reg_module/_04442_ ;
 wire \reg_module/_04443_ ;
 wire \reg_module/_04444_ ;
 wire \reg_module/_04445_ ;
 wire \reg_module/_04446_ ;
 wire \reg_module/_04447_ ;
 wire \reg_module/_04448_ ;
 wire \reg_module/_04449_ ;
 wire \reg_module/_04450_ ;
 wire \reg_module/_04451_ ;
 wire \reg_module/_04452_ ;
 wire \reg_module/_04453_ ;
 wire \reg_module/_04454_ ;
 wire \reg_module/_04455_ ;
 wire \reg_module/_04456_ ;
 wire \reg_module/_04457_ ;
 wire \reg_module/_04458_ ;
 wire \reg_module/_04459_ ;
 wire \reg_module/_04460_ ;
 wire \reg_module/_04461_ ;
 wire \reg_module/_04462_ ;
 wire \reg_module/_04463_ ;
 wire \reg_module/_04464_ ;
 wire \reg_module/_04465_ ;
 wire \reg_module/_04466_ ;
 wire \reg_module/_04467_ ;
 wire \reg_module/_04468_ ;
 wire \reg_module/_04469_ ;
 wire \reg_module/_04470_ ;
 wire \reg_module/_04471_ ;
 wire \reg_module/_04472_ ;
 wire \reg_module/_04473_ ;
 wire \reg_module/_04474_ ;
 wire \reg_module/_04475_ ;
 wire \reg_module/_04476_ ;
 wire \reg_module/_04477_ ;
 wire \reg_module/_04478_ ;
 wire \reg_module/_04479_ ;
 wire \reg_module/_04480_ ;
 wire \reg_module/_04481_ ;
 wire \reg_module/_04482_ ;
 wire \reg_module/_04483_ ;
 wire \reg_module/_04484_ ;
 wire \reg_module/_04485_ ;
 wire \reg_module/_04486_ ;
 wire \reg_module/_04487_ ;
 wire \reg_module/_04488_ ;
 wire \reg_module/_04489_ ;
 wire \reg_module/_04490_ ;
 wire \reg_module/_04491_ ;
 wire \reg_module/_04492_ ;
 wire \reg_module/_04493_ ;
 wire \reg_module/_04494_ ;
 wire \reg_module/_04495_ ;
 wire \reg_module/_04496_ ;
 wire \reg_module/_04497_ ;
 wire \reg_module/_04498_ ;
 wire \reg_module/_04499_ ;
 wire \reg_module/_04500_ ;
 wire \reg_module/_04501_ ;
 wire \reg_module/_04502_ ;
 wire \reg_module/_04503_ ;
 wire \reg_module/_04504_ ;
 wire \reg_module/_04505_ ;
 wire \reg_module/_04506_ ;
 wire \reg_module/_04507_ ;
 wire \reg_module/_04508_ ;
 wire \reg_module/_04509_ ;
 wire \reg_module/_04510_ ;
 wire \reg_module/_04511_ ;
 wire \reg_module/_04512_ ;
 wire \reg_module/_04513_ ;
 wire \reg_module/_04514_ ;
 wire \reg_module/_04515_ ;
 wire \reg_module/_04516_ ;
 wire \reg_module/_04517_ ;
 wire \reg_module/_04518_ ;
 wire \reg_module/_04519_ ;
 wire \reg_module/_04520_ ;
 wire \reg_module/_04521_ ;
 wire \reg_module/_04522_ ;
 wire \reg_module/_04523_ ;
 wire \reg_module/_04524_ ;
 wire \reg_module/_04525_ ;
 wire \reg_module/_04526_ ;
 wire \reg_module/_04527_ ;
 wire \reg_module/_04528_ ;
 wire \reg_module/_04529_ ;
 wire \reg_module/_04530_ ;
 wire \reg_module/_04531_ ;
 wire \reg_module/_04532_ ;
 wire \reg_module/_04533_ ;
 wire \reg_module/_04534_ ;
 wire \reg_module/_04535_ ;
 wire \reg_module/_04536_ ;
 wire \reg_module/_04537_ ;
 wire \reg_module/_04538_ ;
 wire \reg_module/_04539_ ;
 wire \reg_module/_04540_ ;
 wire \reg_module/_04541_ ;
 wire \reg_module/_04542_ ;
 wire \reg_module/_04543_ ;
 wire \reg_module/_04544_ ;
 wire \reg_module/_04545_ ;
 wire \reg_module/_04546_ ;
 wire \reg_module/_04547_ ;
 wire \reg_module/_04548_ ;
 wire \reg_module/_04549_ ;
 wire \reg_module/_04550_ ;
 wire \reg_module/_04551_ ;
 wire \reg_module/_04552_ ;
 wire \reg_module/_04553_ ;
 wire \reg_module/_04554_ ;
 wire \reg_module/_04555_ ;
 wire \reg_module/_04556_ ;
 wire \reg_module/_04557_ ;
 wire \reg_module/_04558_ ;
 wire \reg_module/_04559_ ;
 wire \reg_module/_04560_ ;
 wire \reg_module/_04561_ ;
 wire \reg_module/_04562_ ;
 wire \reg_module/_04563_ ;
 wire \reg_module/_04564_ ;
 wire \reg_module/_04565_ ;
 wire \reg_module/_04566_ ;
 wire \reg_module/_04567_ ;
 wire \reg_module/_04568_ ;
 wire \reg_module/_04569_ ;
 wire \reg_module/_04570_ ;
 wire \reg_module/_04571_ ;
 wire \reg_module/_04572_ ;
 wire \reg_module/_04573_ ;
 wire \reg_module/_04574_ ;
 wire \reg_module/_04575_ ;
 wire \reg_module/_04576_ ;
 wire \reg_module/_04577_ ;
 wire \reg_module/_04578_ ;
 wire \reg_module/_04579_ ;
 wire \reg_module/_04580_ ;
 wire \reg_module/_04581_ ;
 wire \reg_module/_04582_ ;
 wire \reg_module/_04583_ ;
 wire \reg_module/_04584_ ;
 wire \reg_module/_04585_ ;
 wire \reg_module/_04586_ ;
 wire \reg_module/_04587_ ;
 wire \reg_module/_04588_ ;
 wire \reg_module/_04589_ ;
 wire \reg_module/_04590_ ;
 wire \reg_module/_04591_ ;
 wire \reg_module/_04592_ ;
 wire \reg_module/_04593_ ;
 wire \reg_module/_04594_ ;
 wire \reg_module/_04595_ ;
 wire \reg_module/_04596_ ;
 wire \reg_module/_04597_ ;
 wire \reg_module/_04598_ ;
 wire \reg_module/_04599_ ;
 wire \reg_module/_04600_ ;
 wire \reg_module/_04601_ ;
 wire \reg_module/_04602_ ;
 wire \reg_module/_04603_ ;
 wire \reg_module/_04604_ ;
 wire \reg_module/_04605_ ;
 wire \reg_module/_04606_ ;
 wire \reg_module/_04607_ ;
 wire \reg_module/_04608_ ;
 wire \reg_module/_04609_ ;
 wire \reg_module/_04610_ ;
 wire \reg_module/_04611_ ;
 wire \reg_module/_04612_ ;
 wire \reg_module/_04613_ ;
 wire \reg_module/_04614_ ;
 wire \reg_module/_04615_ ;
 wire \reg_module/_04616_ ;
 wire \reg_module/_04617_ ;
 wire \reg_module/_04618_ ;
 wire \reg_module/_04619_ ;
 wire \reg_module/_04620_ ;
 wire \reg_module/_04621_ ;
 wire \reg_module/_04622_ ;
 wire \reg_module/_04623_ ;
 wire \reg_module/_04624_ ;
 wire \reg_module/_04625_ ;
 wire \reg_module/_04626_ ;
 wire \reg_module/_04627_ ;
 wire \reg_module/_04628_ ;
 wire \reg_module/_04629_ ;
 wire \reg_module/_04630_ ;
 wire \reg_module/_04631_ ;
 wire \reg_module/_04632_ ;
 wire \reg_module/_04633_ ;
 wire \reg_module/_04634_ ;
 wire \reg_module/_04635_ ;
 wire \reg_module/_04636_ ;
 wire \reg_module/_04637_ ;
 wire \reg_module/_04638_ ;
 wire \reg_module/_04639_ ;
 wire \reg_module/_04640_ ;
 wire \reg_module/_04641_ ;
 wire \reg_module/_04642_ ;
 wire \reg_module/_04643_ ;
 wire \reg_module/_04644_ ;
 wire \reg_module/_04645_ ;
 wire \reg_module/_04646_ ;
 wire \reg_module/_04647_ ;
 wire \reg_module/_04648_ ;
 wire \reg_module/_04649_ ;
 wire \reg_module/_04650_ ;
 wire \reg_module/_04651_ ;
 wire \reg_module/_04652_ ;
 wire \reg_module/_04653_ ;
 wire \reg_module/_04654_ ;
 wire \reg_module/_04655_ ;
 wire \reg_module/_04656_ ;
 wire \reg_module/_04657_ ;
 wire \reg_module/_04658_ ;
 wire \reg_module/_04659_ ;
 wire \reg_module/_04660_ ;
 wire \reg_module/_04661_ ;
 wire \reg_module/_04662_ ;
 wire \reg_module/_04663_ ;
 wire \reg_module/_04664_ ;
 wire \reg_module/_04665_ ;
 wire \reg_module/_04666_ ;
 wire \reg_module/_04667_ ;
 wire \reg_module/_04668_ ;
 wire \reg_module/_04669_ ;
 wire \reg_module/_04670_ ;
 wire \reg_module/_04671_ ;
 wire \reg_module/_04672_ ;
 wire \reg_module/_04673_ ;
 wire \reg_module/_04674_ ;
 wire \reg_module/_04675_ ;
 wire \reg_module/_04676_ ;
 wire \reg_module/_04677_ ;
 wire \reg_module/_04678_ ;
 wire \reg_module/_04679_ ;
 wire \reg_module/_04680_ ;
 wire \reg_module/_04681_ ;
 wire \reg_module/_04682_ ;
 wire \reg_module/_04683_ ;
 wire \reg_module/_04684_ ;
 wire \reg_module/_04685_ ;
 wire \reg_module/_04686_ ;
 wire \reg_module/_04687_ ;
 wire \reg_module/_04688_ ;
 wire \reg_module/_04689_ ;
 wire \reg_module/_04690_ ;
 wire \reg_module/_04691_ ;
 wire \reg_module/_04692_ ;
 wire \reg_module/_04693_ ;
 wire \reg_module/_04694_ ;
 wire \reg_module/_04695_ ;
 wire \reg_module/_04696_ ;
 wire \reg_module/_04697_ ;
 wire \reg_module/_04698_ ;
 wire \reg_module/_04699_ ;
 wire \reg_module/_04700_ ;
 wire \reg_module/_04701_ ;
 wire \reg_module/_04702_ ;
 wire \reg_module/_04703_ ;
 wire \reg_module/_04704_ ;
 wire \reg_module/_04705_ ;
 wire \reg_module/_04706_ ;
 wire \reg_module/_04707_ ;
 wire \reg_module/_04708_ ;
 wire \reg_module/_04709_ ;
 wire \reg_module/_04710_ ;
 wire \reg_module/_04711_ ;
 wire \reg_module/_04712_ ;
 wire \reg_module/_04713_ ;
 wire \reg_module/_04714_ ;
 wire \reg_module/_04715_ ;
 wire \reg_module/_04716_ ;
 wire \reg_module/_04717_ ;
 wire \reg_module/_04718_ ;
 wire \reg_module/_04719_ ;
 wire \reg_module/_04720_ ;
 wire \reg_module/_04721_ ;
 wire \reg_module/_04722_ ;
 wire \reg_module/_04723_ ;
 wire \reg_module/_04724_ ;
 wire \reg_module/_04725_ ;
 wire \reg_module/_04726_ ;
 wire \reg_module/_04727_ ;
 wire \reg_module/_04728_ ;
 wire \reg_module/_04729_ ;
 wire \reg_module/_04730_ ;
 wire \reg_module/_04731_ ;
 wire \reg_module/_04732_ ;
 wire \reg_module/_04733_ ;
 wire \reg_module/_04734_ ;
 wire \reg_module/_04735_ ;
 wire \reg_module/_04736_ ;
 wire \reg_module/_04737_ ;
 wire \reg_module/_04738_ ;
 wire \reg_module/_04739_ ;
 wire \reg_module/_04740_ ;
 wire \reg_module/_04741_ ;
 wire \reg_module/_04742_ ;
 wire \reg_module/_04743_ ;
 wire \reg_module/_04744_ ;
 wire \reg_module/_04745_ ;
 wire \reg_module/_04746_ ;
 wire \reg_module/_04747_ ;
 wire \reg_module/_04748_ ;
 wire \reg_module/_04749_ ;
 wire \reg_module/_04750_ ;
 wire \reg_module/_04751_ ;
 wire \reg_module/_04752_ ;
 wire \reg_module/_04753_ ;
 wire \reg_module/_04754_ ;
 wire \reg_module/_04755_ ;
 wire \reg_module/_04756_ ;
 wire \reg_module/_04757_ ;
 wire \reg_module/_04758_ ;
 wire \reg_module/_04759_ ;
 wire \reg_module/_04760_ ;
 wire \reg_module/_04761_ ;
 wire \reg_module/_04762_ ;
 wire \reg_module/_04763_ ;
 wire \reg_module/_04764_ ;
 wire \reg_module/_04765_ ;
 wire \reg_module/_04766_ ;
 wire \reg_module/_04767_ ;
 wire \reg_module/_04768_ ;
 wire \reg_module/_04769_ ;
 wire \reg_module/_04770_ ;
 wire \reg_module/_04771_ ;
 wire \reg_module/_04772_ ;
 wire \reg_module/_04773_ ;
 wire \reg_module/_04774_ ;
 wire \reg_module/_04775_ ;
 wire \reg_module/_04776_ ;
 wire \reg_module/_04777_ ;
 wire \reg_module/_04778_ ;
 wire \reg_module/_04779_ ;
 wire \reg_module/_04780_ ;
 wire \reg_module/_04781_ ;
 wire \reg_module/_04782_ ;
 wire \reg_module/_04783_ ;
 wire \reg_module/_04784_ ;
 wire \reg_module/_04785_ ;
 wire \reg_module/_04786_ ;
 wire \reg_module/_04787_ ;
 wire \reg_module/_04788_ ;
 wire \reg_module/_04789_ ;
 wire \reg_module/_04790_ ;
 wire \reg_module/_04791_ ;
 wire \reg_module/_04792_ ;
 wire \reg_module/_04793_ ;
 wire \reg_module/_04794_ ;
 wire \reg_module/_04795_ ;
 wire \reg_module/_04796_ ;
 wire \reg_module/_04797_ ;
 wire \reg_module/_04798_ ;
 wire \reg_module/_04799_ ;
 wire \reg_module/_04800_ ;
 wire \reg_module/_04801_ ;
 wire \reg_module/_04802_ ;
 wire \reg_module/_04803_ ;
 wire \reg_module/_04804_ ;
 wire \reg_module/_04805_ ;
 wire \reg_module/_04806_ ;
 wire \reg_module/_04807_ ;
 wire \reg_module/_04808_ ;
 wire \reg_module/_04809_ ;
 wire \reg_module/_04810_ ;
 wire \reg_module/_04811_ ;
 wire \reg_module/_04812_ ;
 wire \reg_module/_04813_ ;
 wire \reg_module/_04814_ ;
 wire \reg_module/_04815_ ;
 wire \reg_module/_04816_ ;
 wire \reg_module/_04817_ ;
 wire \reg_module/_04818_ ;
 wire \reg_module/_04819_ ;
 wire \reg_module/_04820_ ;
 wire \reg_module/_04821_ ;
 wire \reg_module/_04822_ ;
 wire \reg_module/_04823_ ;
 wire \reg_module/_04824_ ;
 wire \reg_module/_04825_ ;
 wire \reg_module/_04826_ ;
 wire \reg_module/_04827_ ;
 wire \reg_module/_04828_ ;
 wire \reg_module/_04829_ ;
 wire \reg_module/_04830_ ;
 wire \reg_module/_04831_ ;
 wire \reg_module/_04832_ ;
 wire \reg_module/_04833_ ;
 wire \reg_module/_04834_ ;
 wire \reg_module/_04835_ ;
 wire \reg_module/_04836_ ;
 wire \reg_module/_04837_ ;
 wire \reg_module/_04838_ ;
 wire \reg_module/_04839_ ;
 wire \reg_module/_04840_ ;
 wire \reg_module/_04841_ ;
 wire \reg_module/_04842_ ;
 wire \reg_module/_04843_ ;
 wire \reg_module/_04844_ ;
 wire \reg_module/_04845_ ;
 wire \reg_module/_04846_ ;
 wire \reg_module/_04847_ ;
 wire \reg_module/_04848_ ;
 wire \reg_module/_04849_ ;
 wire \reg_module/_04850_ ;
 wire \reg_module/_04851_ ;
 wire \reg_module/_04852_ ;
 wire \reg_module/_04853_ ;
 wire \reg_module/_04854_ ;
 wire \reg_module/_04855_ ;
 wire \reg_module/_04856_ ;
 wire \reg_module/_04857_ ;
 wire \reg_module/_04858_ ;
 wire \reg_module/_04859_ ;
 wire \reg_module/_04860_ ;
 wire \reg_module/_04861_ ;
 wire \reg_module/_04862_ ;
 wire \reg_module/_04863_ ;
 wire \reg_module/_04864_ ;
 wire \reg_module/_04865_ ;
 wire \reg_module/_04866_ ;
 wire \reg_module/_04867_ ;
 wire \reg_module/_04868_ ;
 wire \reg_module/_04869_ ;
 wire \reg_module/_04870_ ;
 wire \reg_module/_04871_ ;
 wire \reg_module/_04872_ ;
 wire \reg_module/_04873_ ;
 wire \reg_module/_04874_ ;
 wire \reg_module/_04875_ ;
 wire \reg_module/_04876_ ;
 wire \reg_module/_04877_ ;
 wire \reg_module/_04878_ ;
 wire \reg_module/_04879_ ;
 wire \reg_module/_04880_ ;
 wire \reg_module/_04881_ ;
 wire \reg_module/_04882_ ;
 wire \reg_module/_04883_ ;
 wire \reg_module/_04884_ ;
 wire \reg_module/_04885_ ;
 wire \reg_module/_04886_ ;
 wire \reg_module/_04887_ ;
 wire \reg_module/_04888_ ;
 wire \reg_module/_04889_ ;
 wire \reg_module/_04890_ ;
 wire \reg_module/_04891_ ;
 wire \reg_module/_04892_ ;
 wire \reg_module/_04893_ ;
 wire \reg_module/_04894_ ;
 wire \reg_module/_04895_ ;
 wire \reg_module/_04896_ ;
 wire \reg_module/_04897_ ;
 wire \reg_module/_04898_ ;
 wire \reg_module/_04899_ ;
 wire \reg_module/_04900_ ;
 wire \reg_module/_04901_ ;
 wire \reg_module/_04902_ ;
 wire \reg_module/_04903_ ;
 wire \reg_module/_04904_ ;
 wire \reg_module/_04905_ ;
 wire \reg_module/_04906_ ;
 wire \reg_module/_04907_ ;
 wire \reg_module/_04908_ ;
 wire \reg_module/_04909_ ;
 wire \reg_module/_04910_ ;
 wire \reg_module/_04911_ ;
 wire \reg_module/_04912_ ;
 wire \reg_module/_04913_ ;
 wire \reg_module/_04914_ ;
 wire \reg_module/_04915_ ;
 wire \reg_module/_04916_ ;
 wire \reg_module/_04917_ ;
 wire \reg_module/_04918_ ;
 wire \reg_module/_04919_ ;
 wire \reg_module/_04920_ ;
 wire \reg_module/_04921_ ;
 wire \reg_module/_04922_ ;
 wire \reg_module/_04923_ ;
 wire \reg_module/_04924_ ;
 wire \reg_module/_04925_ ;
 wire \reg_module/_04926_ ;
 wire \reg_module/_04927_ ;
 wire \reg_module/_04928_ ;
 wire \reg_module/_04929_ ;
 wire \reg_module/_04930_ ;
 wire \reg_module/_04931_ ;
 wire \reg_module/_04932_ ;
 wire \reg_module/_04933_ ;
 wire \reg_module/_04934_ ;
 wire \reg_module/_04935_ ;
 wire \reg_module/_04936_ ;
 wire \reg_module/_04937_ ;
 wire \reg_module/_04938_ ;
 wire \reg_module/_04939_ ;
 wire \reg_module/_04940_ ;
 wire \reg_module/_04941_ ;
 wire \reg_module/_04942_ ;
 wire \reg_module/_04943_ ;
 wire \reg_module/_04944_ ;
 wire \reg_module/_04945_ ;
 wire \reg_module/_04946_ ;
 wire \reg_module/_04947_ ;
 wire \reg_module/_04948_ ;
 wire \reg_module/_04949_ ;
 wire \reg_module/_04950_ ;
 wire \reg_module/_04951_ ;
 wire \reg_module/_04952_ ;
 wire \reg_module/_04953_ ;
 wire \reg_module/_04954_ ;
 wire \reg_module/_04955_ ;
 wire \reg_module/_04956_ ;
 wire \reg_module/_04957_ ;
 wire \reg_module/_04958_ ;
 wire \reg_module/_04959_ ;
 wire \reg_module/_04960_ ;
 wire \reg_module/_04961_ ;
 wire \reg_module/_04962_ ;
 wire \reg_module/_04963_ ;
 wire \reg_module/_04964_ ;
 wire \reg_module/_04965_ ;
 wire \reg_module/_04966_ ;
 wire \reg_module/_04967_ ;
 wire \reg_module/_04968_ ;
 wire \reg_module/_04969_ ;
 wire \reg_module/_04970_ ;
 wire \reg_module/_04971_ ;
 wire \reg_module/_04972_ ;
 wire \reg_module/_04973_ ;
 wire \reg_module/_04974_ ;
 wire \reg_module/_04975_ ;
 wire \reg_module/_04976_ ;
 wire \reg_module/_04977_ ;
 wire \reg_module/_04978_ ;
 wire \reg_module/_04979_ ;
 wire \reg_module/_04980_ ;
 wire \reg_module/_04981_ ;
 wire \reg_module/_04982_ ;
 wire \reg_module/_04983_ ;
 wire \reg_module/_04984_ ;
 wire \reg_module/_04985_ ;
 wire \reg_module/_04986_ ;
 wire \reg_module/_04987_ ;
 wire \reg_module/_04988_ ;
 wire \reg_module/_04989_ ;
 wire \reg_module/_04990_ ;
 wire \reg_module/_04991_ ;
 wire \reg_module/_04992_ ;
 wire \reg_module/_04993_ ;
 wire \reg_module/_04994_ ;
 wire \reg_module/_04995_ ;
 wire \reg_module/_04996_ ;
 wire \reg_module/_04997_ ;
 wire \reg_module/_04998_ ;
 wire \reg_module/_04999_ ;
 wire \reg_module/_05000_ ;
 wire \reg_module/_05001_ ;
 wire \reg_module/_05002_ ;
 wire \reg_module/_05003_ ;
 wire \reg_module/_05004_ ;
 wire \reg_module/_05005_ ;
 wire \reg_module/_05006_ ;
 wire \reg_module/_05007_ ;
 wire \reg_module/_05008_ ;
 wire \reg_module/_05009_ ;
 wire \reg_module/_05010_ ;
 wire \reg_module/_05011_ ;
 wire \reg_module/_05012_ ;
 wire \reg_module/_05013_ ;
 wire \reg_module/_05014_ ;
 wire \reg_module/_05015_ ;
 wire \reg_module/_05016_ ;
 wire \reg_module/_05017_ ;
 wire \reg_module/_05018_ ;
 wire \reg_module/_05019_ ;
 wire \reg_module/_05020_ ;
 wire \reg_module/_05021_ ;
 wire \reg_module/_05022_ ;
 wire \reg_module/_05023_ ;
 wire \reg_module/_05024_ ;
 wire \reg_module/_05025_ ;
 wire \reg_module/_05026_ ;
 wire \reg_module/_05027_ ;
 wire \reg_module/_05028_ ;
 wire \reg_module/_05029_ ;
 wire \reg_module/_05030_ ;
 wire \reg_module/_05031_ ;
 wire \reg_module/_05032_ ;
 wire \reg_module/_05033_ ;
 wire \reg_module/_05034_ ;
 wire \reg_module/_05035_ ;
 wire \reg_module/_05036_ ;
 wire \reg_module/_05037_ ;
 wire \reg_module/_05038_ ;
 wire \reg_module/_05039_ ;
 wire \reg_module/_05040_ ;
 wire \reg_module/_05041_ ;
 wire \reg_module/_05042_ ;
 wire \reg_module/_05043_ ;
 wire \reg_module/_05044_ ;
 wire \reg_module/_05045_ ;
 wire \reg_module/_05046_ ;
 wire \reg_module/_05047_ ;
 wire \reg_module/_05048_ ;
 wire \reg_module/_05049_ ;
 wire \reg_module/_05050_ ;
 wire \reg_module/_05051_ ;
 wire \reg_module/_05052_ ;
 wire \reg_module/_05053_ ;
 wire \reg_module/_05054_ ;
 wire \reg_module/_05055_ ;
 wire \reg_module/_05056_ ;
 wire \reg_module/_05057_ ;
 wire \reg_module/_05058_ ;
 wire \reg_module/_05059_ ;
 wire \reg_module/_05060_ ;
 wire \reg_module/_05061_ ;
 wire \reg_module/_05062_ ;
 wire \reg_module/_05063_ ;
 wire \reg_module/_05064_ ;
 wire \reg_module/_05065_ ;
 wire \reg_module/_05066_ ;
 wire \reg_module/_05067_ ;
 wire \reg_module/_05068_ ;
 wire \reg_module/_05069_ ;
 wire \reg_module/_05070_ ;
 wire \reg_module/_05071_ ;
 wire \reg_module/_05072_ ;
 wire \reg_module/_05073_ ;
 wire \reg_module/_05074_ ;
 wire \reg_module/_05075_ ;
 wire \reg_module/_05076_ ;
 wire \reg_module/_05077_ ;
 wire \reg_module/_05078_ ;
 wire \reg_module/_05079_ ;
 wire \reg_module/_05080_ ;
 wire \reg_module/_05081_ ;
 wire \reg_module/_05082_ ;
 wire \reg_module/_05083_ ;
 wire \reg_module/_05084_ ;
 wire \reg_module/_05085_ ;
 wire \reg_module/_05086_ ;
 wire \reg_module/_05087_ ;
 wire \reg_module/_05088_ ;
 wire \reg_module/_05089_ ;
 wire \reg_module/_05090_ ;
 wire \reg_module/_05091_ ;
 wire \reg_module/_05092_ ;
 wire \reg_module/_05093_ ;
 wire \reg_module/_05094_ ;
 wire \reg_module/_05095_ ;
 wire \reg_module/_05096_ ;
 wire \reg_module/_05097_ ;
 wire \reg_module/_05098_ ;
 wire \reg_module/_05099_ ;
 wire \reg_module/_05100_ ;
 wire \reg_module/_05101_ ;
 wire \reg_module/_05102_ ;
 wire \reg_module/_05103_ ;
 wire \reg_module/_05104_ ;
 wire \reg_module/_05105_ ;
 wire \reg_module/_05106_ ;
 wire \reg_module/_05107_ ;
 wire \reg_module/_05108_ ;
 wire \reg_module/_05109_ ;
 wire \reg_module/_05110_ ;
 wire \reg_module/_05111_ ;
 wire \reg_module/_05112_ ;
 wire \reg_module/_05113_ ;
 wire \reg_module/_05114_ ;
 wire \reg_module/_05115_ ;
 wire \reg_module/_05116_ ;
 wire \reg_module/_05117_ ;
 wire \reg_module/_05118_ ;
 wire \reg_module/_05119_ ;
 wire \reg_module/_05120_ ;
 wire \reg_module/_05121_ ;
 wire \reg_module/_05122_ ;
 wire \reg_module/_05123_ ;
 wire \reg_module/_05124_ ;
 wire \reg_module/_05125_ ;
 wire \reg_module/_05126_ ;
 wire \reg_module/_05127_ ;
 wire \reg_module/_05128_ ;
 wire \reg_module/_05129_ ;
 wire \reg_module/_05130_ ;
 wire \reg_module/_05131_ ;
 wire \reg_module/_05132_ ;
 wire \reg_module/_05133_ ;
 wire \reg_module/_05134_ ;
 wire \reg_module/_05135_ ;
 wire \reg_module/_05136_ ;
 wire \reg_module/_05137_ ;
 wire \reg_module/_05138_ ;
 wire \reg_module/_05139_ ;
 wire \reg_module/_05140_ ;
 wire \reg_module/_05141_ ;
 wire \reg_module/_05142_ ;
 wire \reg_module/_05143_ ;
 wire \reg_module/_05144_ ;
 wire \reg_module/_05145_ ;
 wire \reg_module/_05146_ ;
 wire \reg_module/_05147_ ;
 wire \reg_module/_05148_ ;
 wire \reg_module/_05149_ ;
 wire \reg_module/_05150_ ;
 wire \reg_module/_05151_ ;
 wire \reg_module/_05152_ ;
 wire \reg_module/_05153_ ;
 wire \reg_module/_05154_ ;
 wire \reg_module/_05155_ ;
 wire \reg_module/_05156_ ;
 wire \reg_module/_05157_ ;
 wire \reg_module/_05158_ ;
 wire \reg_module/_05159_ ;
 wire \reg_module/_05160_ ;
 wire \reg_module/_05161_ ;
 wire \reg_module/_05162_ ;
 wire \reg_module/_05163_ ;
 wire \reg_module/_05164_ ;
 wire \reg_module/_05165_ ;
 wire \reg_module/_05166_ ;
 wire \reg_module/_05167_ ;
 wire \reg_module/_05168_ ;
 wire \reg_module/_05169_ ;
 wire \reg_module/_05170_ ;
 wire \reg_module/_05171_ ;
 wire \reg_module/_05172_ ;
 wire \reg_module/_05173_ ;
 wire \reg_module/_05174_ ;
 wire \reg_module/_05175_ ;
 wire \reg_module/_05176_ ;
 wire \reg_module/_05177_ ;
 wire \reg_module/_05178_ ;
 wire \reg_module/_05179_ ;
 wire \reg_module/_05180_ ;
 wire \reg_module/_05181_ ;
 wire \reg_module/_05182_ ;
 wire \reg_module/_05183_ ;
 wire \reg_module/_05184_ ;
 wire \reg_module/_05185_ ;
 wire \reg_module/_05186_ ;
 wire \reg_module/_05187_ ;
 wire \reg_module/_05188_ ;
 wire \reg_module/_05189_ ;
 wire \reg_module/_05190_ ;
 wire \reg_module/_05191_ ;
 wire \reg_module/_05192_ ;
 wire \reg_module/_05193_ ;
 wire \reg_module/_05194_ ;
 wire \reg_module/_05195_ ;
 wire \reg_module/_05196_ ;
 wire \reg_module/_05197_ ;
 wire \reg_module/_05198_ ;
 wire \reg_module/_05199_ ;
 wire \reg_module/_05200_ ;
 wire \reg_module/_05201_ ;
 wire \reg_module/_05202_ ;
 wire \reg_module/_05203_ ;
 wire \reg_module/_05204_ ;
 wire \reg_module/_05205_ ;
 wire \reg_module/_05206_ ;
 wire \reg_module/_05207_ ;
 wire \reg_module/_05208_ ;
 wire \reg_module/_05209_ ;
 wire \reg_module/_05210_ ;
 wire \reg_module/_05211_ ;
 wire \reg_module/_05212_ ;
 wire \reg_module/_05213_ ;
 wire \reg_module/_05214_ ;
 wire \reg_module/_05215_ ;
 wire \reg_module/_05216_ ;
 wire \reg_module/_05217_ ;
 wire \reg_module/_05218_ ;
 wire \reg_module/_05219_ ;
 wire \reg_module/_05220_ ;
 wire \reg_module/_05221_ ;
 wire \reg_module/_05222_ ;
 wire \reg_module/_05223_ ;
 wire \reg_module/_05224_ ;
 wire \reg_module/_05225_ ;
 wire \reg_module/_05226_ ;
 wire \reg_module/_05227_ ;
 wire \reg_module/_05228_ ;
 wire \reg_module/_05229_ ;
 wire \reg_module/_05230_ ;
 wire \reg_module/_05231_ ;
 wire \reg_module/_05232_ ;
 wire \reg_module/_05233_ ;
 wire \reg_module/_05234_ ;
 wire \reg_module/_05235_ ;
 wire \reg_module/_05236_ ;
 wire \reg_module/_05237_ ;
 wire \reg_module/_05238_ ;
 wire \reg_module/_05239_ ;
 wire \reg_module/_05240_ ;
 wire \reg_module/_05241_ ;
 wire \reg_module/_05242_ ;
 wire \reg_module/_05243_ ;
 wire \reg_module/_05244_ ;
 wire \reg_module/_05245_ ;
 wire \reg_module/_05246_ ;
 wire \reg_module/_05247_ ;
 wire \reg_module/_05248_ ;
 wire \reg_module/_05249_ ;
 wire \reg_module/_05250_ ;
 wire \reg_module/_05251_ ;
 wire \reg_module/_05252_ ;
 wire \reg_module/_05253_ ;
 wire \reg_module/_05254_ ;
 wire \reg_module/_05255_ ;
 wire \reg_module/_05256_ ;
 wire \reg_module/_05257_ ;
 wire \reg_module/_05258_ ;
 wire \reg_module/_05259_ ;
 wire \reg_module/_05260_ ;
 wire \reg_module/_05261_ ;
 wire \reg_module/_05262_ ;
 wire \reg_module/_05263_ ;
 wire \reg_module/_05264_ ;
 wire \reg_module/_05265_ ;
 wire \reg_module/_05266_ ;
 wire \reg_module/_05267_ ;
 wire \reg_module/_05268_ ;
 wire \reg_module/_05269_ ;
 wire \reg_module/_05270_ ;
 wire \reg_module/_05271_ ;
 wire \reg_module/_05272_ ;
 wire \reg_module/_05273_ ;
 wire \reg_module/_05274_ ;
 wire \reg_module/_05275_ ;
 wire \reg_module/_05276_ ;
 wire \reg_module/_05277_ ;
 wire \reg_module/_05278_ ;
 wire \reg_module/_05279_ ;
 wire \reg_module/_05280_ ;
 wire \reg_module/_05281_ ;
 wire \reg_module/_05282_ ;
 wire \reg_module/_05283_ ;
 wire \reg_module/_05284_ ;
 wire \reg_module/_05285_ ;
 wire \reg_module/_05286_ ;
 wire \reg_module/_05287_ ;
 wire \reg_module/_05288_ ;
 wire \reg_module/_05289_ ;
 wire \reg_module/_05290_ ;
 wire \reg_module/_05291_ ;
 wire \reg_module/_05292_ ;
 wire \reg_module/_05293_ ;
 wire \reg_module/_05294_ ;
 wire \reg_module/_05295_ ;
 wire \reg_module/_05296_ ;
 wire \reg_module/_05297_ ;
 wire \reg_module/_05298_ ;
 wire \reg_module/_05299_ ;
 wire \reg_module/_05300_ ;
 wire \reg_module/_05301_ ;
 wire \reg_module/_05302_ ;
 wire \reg_module/_05303_ ;
 wire \reg_module/_05304_ ;
 wire \reg_module/_05305_ ;
 wire \reg_module/_05306_ ;
 wire \reg_module/_05307_ ;
 wire \reg_module/_05308_ ;
 wire \reg_module/_05309_ ;
 wire \reg_module/_05310_ ;
 wire \reg_module/_05311_ ;
 wire \reg_module/_05312_ ;
 wire \reg_module/_05313_ ;
 wire \reg_module/_05314_ ;
 wire \reg_module/_05315_ ;
 wire \reg_module/_05316_ ;
 wire \reg_module/_05317_ ;
 wire \reg_module/_05318_ ;
 wire \reg_module/_05319_ ;
 wire \reg_module/_05320_ ;
 wire \reg_module/_05321_ ;
 wire \reg_module/_05322_ ;
 wire \reg_module/_05323_ ;
 wire \reg_module/_05324_ ;
 wire \reg_module/_05325_ ;
 wire \reg_module/_05326_ ;
 wire \reg_module/_05327_ ;
 wire \reg_module/_05328_ ;
 wire \reg_module/_05329_ ;
 wire \reg_module/_05330_ ;
 wire \reg_module/_05331_ ;
 wire \reg_module/_05332_ ;
 wire \reg_module/_05333_ ;
 wire \reg_module/_05334_ ;
 wire \reg_module/_05335_ ;
 wire \reg_module/_05336_ ;
 wire \reg_module/_05337_ ;
 wire \reg_module/_05338_ ;
 wire \reg_module/_05339_ ;
 wire \reg_module/_05340_ ;
 wire \reg_module/_05341_ ;
 wire \reg_module/_05342_ ;
 wire \reg_module/_05343_ ;
 wire \reg_module/_05344_ ;
 wire \reg_module/_05345_ ;
 wire \reg_module/_05346_ ;
 wire \reg_module/_05347_ ;
 wire \reg_module/_05348_ ;
 wire \reg_module/_05349_ ;
 wire \reg_module/_05350_ ;
 wire \reg_module/_05351_ ;
 wire \reg_module/_05352_ ;
 wire \reg_module/_05353_ ;
 wire \reg_module/_05354_ ;
 wire \reg_module/_05355_ ;
 wire \reg_module/_05356_ ;
 wire \reg_module/_05357_ ;
 wire \reg_module/_05358_ ;
 wire \reg_module/_05359_ ;
 wire \reg_module/_05360_ ;
 wire \reg_module/_05361_ ;
 wire \reg_module/_05362_ ;
 wire \reg_module/_05363_ ;
 wire \reg_module/_05364_ ;
 wire \reg_module/_05365_ ;
 wire \reg_module/_05366_ ;
 wire \reg_module/_05367_ ;
 wire \reg_module/_05368_ ;
 wire \reg_module/_05369_ ;
 wire \reg_module/_05370_ ;
 wire \reg_module/_05371_ ;
 wire \reg_module/_05372_ ;
 wire \reg_module/_05373_ ;
 wire \reg_module/_05374_ ;
 wire \reg_module/_05375_ ;
 wire \reg_module/_05376_ ;
 wire \reg_module/_05377_ ;
 wire \reg_module/_05378_ ;
 wire \reg_module/_05379_ ;
 wire \reg_module/_05380_ ;
 wire \reg_module/_05381_ ;
 wire \reg_module/_05382_ ;
 wire \reg_module/_05383_ ;
 wire \reg_module/_05384_ ;
 wire \reg_module/_05385_ ;
 wire \reg_module/_05386_ ;
 wire \reg_module/_05387_ ;
 wire \reg_module/_05388_ ;
 wire \reg_module/_05389_ ;
 wire \reg_module/_05390_ ;
 wire \reg_module/_05391_ ;
 wire \reg_module/_05392_ ;
 wire \reg_module/_05393_ ;
 wire \reg_module/_05394_ ;
 wire \reg_module/_05395_ ;
 wire \reg_module/_05396_ ;
 wire \reg_module/_05397_ ;
 wire \reg_module/_05398_ ;
 wire \reg_module/_05399_ ;
 wire \reg_module/_05400_ ;
 wire \reg_module/_05401_ ;
 wire \reg_module/_05402_ ;
 wire \reg_module/_05403_ ;
 wire \reg_module/_05404_ ;
 wire \reg_module/_05405_ ;
 wire \reg_module/_05406_ ;
 wire \reg_module/_05407_ ;
 wire \reg_module/_05408_ ;
 wire \reg_module/_05409_ ;
 wire \reg_module/_05410_ ;
 wire \reg_module/_05411_ ;
 wire \reg_module/_05412_ ;
 wire \reg_module/_05413_ ;
 wire \reg_module/_05414_ ;
 wire \reg_module/_05415_ ;
 wire \reg_module/_05416_ ;
 wire \reg_module/_05417_ ;
 wire \reg_module/_05418_ ;
 wire \reg_module/_05419_ ;
 wire \reg_module/_05420_ ;
 wire \reg_module/_05421_ ;
 wire \reg_module/_05422_ ;
 wire \reg_module/_05423_ ;
 wire \reg_module/_05424_ ;
 wire \reg_module/_05425_ ;
 wire \reg_module/_05426_ ;
 wire \reg_module/_05427_ ;
 wire \reg_module/_05428_ ;
 wire \reg_module/_05429_ ;
 wire \reg_module/_05430_ ;
 wire \reg_module/_05431_ ;
 wire \reg_module/_05432_ ;
 wire \reg_module/_05433_ ;
 wire \reg_module/_05434_ ;
 wire \reg_module/_05435_ ;
 wire \reg_module/_05436_ ;
 wire \reg_module/_05437_ ;
 wire \reg_module/_05438_ ;
 wire \reg_module/_05439_ ;
 wire \reg_module/_05440_ ;
 wire \reg_module/_05441_ ;
 wire \reg_module/_05442_ ;
 wire \reg_module/_05443_ ;
 wire \reg_module/_05444_ ;
 wire \reg_module/_05445_ ;
 wire \reg_module/_05446_ ;
 wire \reg_module/_05447_ ;
 wire \reg_module/_05448_ ;
 wire \reg_module/_05449_ ;
 wire \reg_module/_05450_ ;
 wire \reg_module/_05451_ ;
 wire \reg_module/_05452_ ;
 wire \reg_module/_05453_ ;
 wire \reg_module/_05454_ ;
 wire \reg_module/_05455_ ;
 wire \reg_module/_05456_ ;
 wire \reg_module/_05457_ ;
 wire \reg_module/_05458_ ;
 wire \reg_module/_05459_ ;
 wire \reg_module/_05460_ ;
 wire \reg_module/_05461_ ;
 wire \reg_module/_05462_ ;
 wire \reg_module/_05463_ ;
 wire \reg_module/_05464_ ;
 wire \reg_module/_05465_ ;
 wire \reg_module/_05466_ ;
 wire \reg_module/_05467_ ;
 wire \reg_module/_05468_ ;
 wire \reg_module/_05469_ ;
 wire \reg_module/_05470_ ;
 wire \reg_module/_05471_ ;
 wire \reg_module/_05472_ ;
 wire \reg_module/_05473_ ;
 wire \reg_module/_05474_ ;
 wire \reg_module/_05475_ ;
 wire \reg_module/_05476_ ;
 wire \reg_module/_05477_ ;
 wire \reg_module/_05478_ ;
 wire \reg_module/_05479_ ;
 wire \reg_module/_05480_ ;
 wire \reg_module/_05481_ ;
 wire \reg_module/_05482_ ;
 wire \reg_module/_05483_ ;
 wire \reg_module/_05484_ ;
 wire \reg_module/_05485_ ;
 wire \reg_module/_05486_ ;
 wire \reg_module/_05487_ ;
 wire \reg_module/_05488_ ;
 wire \reg_module/_05489_ ;
 wire \reg_module/_05490_ ;
 wire \reg_module/_05491_ ;
 wire \reg_module/_05492_ ;
 wire \reg_module/_05493_ ;
 wire \reg_module/_05494_ ;
 wire \reg_module/_05495_ ;
 wire \reg_module/_05496_ ;
 wire \reg_module/_05497_ ;
 wire \reg_module/_05498_ ;
 wire \reg_module/_05499_ ;
 wire \reg_module/_05500_ ;
 wire \reg_module/_05501_ ;
 wire \reg_module/_05502_ ;
 wire \reg_module/_05503_ ;
 wire \reg_module/_05504_ ;
 wire \reg_module/_05505_ ;
 wire \reg_module/_05506_ ;
 wire \reg_module/_05507_ ;
 wire \reg_module/_05508_ ;
 wire \reg_module/_05509_ ;
 wire \reg_module/_05510_ ;
 wire \reg_module/_05511_ ;
 wire \reg_module/_05512_ ;
 wire \reg_module/_05513_ ;
 wire \reg_module/_05514_ ;
 wire \reg_module/_05515_ ;
 wire \reg_module/_05516_ ;
 wire \reg_module/_05517_ ;
 wire \reg_module/_05518_ ;
 wire \reg_module/_05519_ ;
 wire \reg_module/_05520_ ;
 wire \reg_module/_05521_ ;
 wire \reg_module/_05522_ ;
 wire \reg_module/_05523_ ;
 wire \reg_module/_05524_ ;
 wire \reg_module/_05525_ ;
 wire \reg_module/_05526_ ;
 wire \reg_module/_05527_ ;
 wire \reg_module/_05528_ ;
 wire \reg_module/_05529_ ;
 wire \reg_module/_05530_ ;
 wire \reg_module/_05531_ ;
 wire \reg_module/_05532_ ;
 wire \reg_module/_05533_ ;
 wire \reg_module/_05534_ ;
 wire \reg_module/_05535_ ;
 wire \reg_module/_05536_ ;
 wire \reg_module/_05537_ ;
 wire \reg_module/_05538_ ;
 wire \reg_module/_05539_ ;
 wire \reg_module/_05540_ ;
 wire \reg_module/_05541_ ;
 wire \reg_module/_05542_ ;
 wire \reg_module/_05543_ ;
 wire \reg_module/_05544_ ;
 wire \reg_module/_05545_ ;
 wire \reg_module/_05546_ ;
 wire \reg_module/_05547_ ;
 wire \reg_module/_05548_ ;
 wire \reg_module/_05549_ ;
 wire \reg_module/_05550_ ;
 wire \reg_module/_05551_ ;
 wire \reg_module/_05552_ ;
 wire \reg_module/_05553_ ;
 wire \reg_module/_05554_ ;
 wire \reg_module/_05555_ ;
 wire \reg_module/_05556_ ;
 wire \reg_module/_05557_ ;
 wire \reg_module/_05558_ ;
 wire \reg_module/_05559_ ;
 wire \reg_module/_05560_ ;
 wire \reg_module/_05561_ ;
 wire \reg_module/_05562_ ;
 wire \reg_module/_05563_ ;
 wire \reg_module/_05564_ ;
 wire \reg_module/_05565_ ;
 wire \reg_module/_05566_ ;
 wire \reg_module/_05567_ ;
 wire \reg_module/_05568_ ;
 wire \reg_module/_05569_ ;
 wire \reg_module/_05570_ ;
 wire \reg_module/_05571_ ;
 wire \reg_module/_05572_ ;
 wire \reg_module/_05573_ ;
 wire \reg_module/_05574_ ;
 wire \reg_module/_05575_ ;
 wire \reg_module/_05576_ ;
 wire \reg_module/_05577_ ;
 wire \reg_module/_05578_ ;
 wire \reg_module/_05579_ ;
 wire \reg_module/_05580_ ;
 wire \reg_module/_05581_ ;
 wire \reg_module/_05582_ ;
 wire \reg_module/_05583_ ;
 wire \reg_module/_05584_ ;
 wire \reg_module/_05585_ ;
 wire \reg_module/_05586_ ;
 wire \reg_module/_05587_ ;
 wire \reg_module/_05588_ ;
 wire \reg_module/_05589_ ;
 wire \reg_module/_05590_ ;
 wire \reg_module/_05591_ ;
 wire \reg_module/_05592_ ;
 wire \reg_module/_05593_ ;
 wire \reg_module/_05594_ ;
 wire \reg_module/_05595_ ;
 wire \reg_module/_05596_ ;
 wire \reg_module/_05597_ ;
 wire \reg_module/_05598_ ;
 wire \reg_module/_05599_ ;
 wire \reg_module/_05600_ ;
 wire \reg_module/_05601_ ;
 wire \reg_module/_05602_ ;
 wire \reg_module/_05603_ ;
 wire \reg_module/_05604_ ;
 wire \reg_module/_05605_ ;
 wire \reg_module/_05606_ ;
 wire \reg_module/_05607_ ;
 wire \reg_module/_05608_ ;
 wire \reg_module/_05609_ ;
 wire \reg_module/_05610_ ;
 wire \reg_module/_05611_ ;
 wire \reg_module/_05612_ ;
 wire \reg_module/_05613_ ;
 wire \reg_module/_05614_ ;
 wire \reg_module/_05615_ ;
 wire \reg_module/_05616_ ;
 wire \reg_module/_05617_ ;
 wire \reg_module/_05618_ ;
 wire \reg_module/_05619_ ;
 wire \reg_module/_05620_ ;
 wire \reg_module/_05621_ ;
 wire \reg_module/_05622_ ;
 wire \reg_module/_05623_ ;
 wire \reg_module/_05624_ ;
 wire \reg_module/_05625_ ;
 wire \reg_module/_05626_ ;
 wire \reg_module/_05627_ ;
 wire \reg_module/_05628_ ;
 wire \reg_module/_05629_ ;
 wire \reg_module/_05630_ ;
 wire \reg_module/_05631_ ;
 wire \reg_module/_05632_ ;
 wire \reg_module/_05633_ ;
 wire \reg_module/_05634_ ;
 wire \reg_module/_05635_ ;
 wire \reg_module/_05636_ ;
 wire \reg_module/_05637_ ;
 wire \reg_module/_05638_ ;
 wire \reg_module/_05639_ ;
 wire \reg_module/_05640_ ;
 wire \reg_module/_05641_ ;
 wire \reg_module/_05642_ ;
 wire \reg_module/_05643_ ;
 wire \reg_module/_05644_ ;
 wire \reg_module/_05645_ ;
 wire \reg_module/_05646_ ;
 wire \reg_module/_05647_ ;
 wire \reg_module/_05648_ ;
 wire \reg_module/_05649_ ;
 wire \reg_module/_05650_ ;
 wire \reg_module/_05651_ ;
 wire \reg_module/_05652_ ;
 wire \reg_module/_05653_ ;
 wire \reg_module/_05654_ ;
 wire \reg_module/_05655_ ;
 wire \reg_module/_05656_ ;
 wire \reg_module/_05657_ ;
 wire \reg_module/_05658_ ;
 wire \reg_module/_05659_ ;
 wire \reg_module/_05660_ ;
 wire \reg_module/_05661_ ;
 wire \reg_module/_05662_ ;
 wire \reg_module/_05663_ ;
 wire \reg_module/_05664_ ;
 wire \reg_module/_05665_ ;
 wire \reg_module/_05666_ ;
 wire \reg_module/_05667_ ;
 wire \reg_module/_05668_ ;
 wire \reg_module/_05669_ ;
 wire \reg_module/_05670_ ;
 wire \reg_module/_05671_ ;
 wire \reg_module/_05672_ ;
 wire \reg_module/_05673_ ;
 wire \reg_module/_05674_ ;
 wire \reg_module/_05675_ ;
 wire \reg_module/_05676_ ;
 wire \reg_module/_05677_ ;
 wire \reg_module/_05678_ ;
 wire \reg_module/_05679_ ;
 wire \reg_module/_05680_ ;
 wire \reg_module/_05681_ ;
 wire \reg_module/_05682_ ;
 wire \reg_module/_05683_ ;
 wire \reg_module/_05684_ ;
 wire \reg_module/_05685_ ;
 wire \reg_module/_05686_ ;
 wire \reg_module/_05687_ ;
 wire \reg_module/_05688_ ;
 wire \reg_module/_05689_ ;
 wire \reg_module/_05690_ ;
 wire \reg_module/_05691_ ;
 wire \reg_module/_05692_ ;
 wire \reg_module/_05693_ ;
 wire \reg_module/_05694_ ;
 wire \reg_module/_05695_ ;
 wire \reg_module/_05696_ ;
 wire \reg_module/_05697_ ;
 wire \reg_module/_05698_ ;
 wire \reg_module/_05699_ ;
 wire \reg_module/_05700_ ;
 wire \reg_module/_05701_ ;
 wire \reg_module/_05702_ ;
 wire \reg_module/_05703_ ;
 wire \reg_module/_05704_ ;
 wire \reg_module/_05705_ ;
 wire \reg_module/_05706_ ;
 wire \reg_module/_05707_ ;
 wire \reg_module/_05708_ ;
 wire \reg_module/_05709_ ;
 wire \reg_module/_05710_ ;
 wire \reg_module/_05711_ ;
 wire \reg_module/_05712_ ;
 wire \reg_module/_05713_ ;
 wire \reg_module/_05714_ ;
 wire \reg_module/_05715_ ;
 wire \reg_module/_05716_ ;
 wire \reg_module/_05717_ ;
 wire \reg_module/_05718_ ;
 wire \reg_module/_05719_ ;
 wire \reg_module/_05720_ ;
 wire \reg_module/_05721_ ;
 wire \reg_module/_05722_ ;
 wire \reg_module/_05723_ ;
 wire \reg_module/_05724_ ;
 wire \reg_module/_05725_ ;
 wire \reg_module/_05726_ ;
 wire \reg_module/_05727_ ;
 wire \reg_module/_05728_ ;
 wire \reg_module/_05729_ ;
 wire \reg_module/_05730_ ;
 wire \reg_module/_05731_ ;
 wire \reg_module/_05732_ ;
 wire \reg_module/_05733_ ;
 wire \reg_module/_05734_ ;
 wire \reg_module/_05735_ ;
 wire \reg_module/_05736_ ;
 wire \reg_module/_05737_ ;
 wire \reg_module/_05738_ ;
 wire \reg_module/_05739_ ;
 wire \reg_module/_05740_ ;
 wire \reg_module/_05741_ ;
 wire \reg_module/_05742_ ;
 wire \reg_module/_05743_ ;
 wire \reg_module/_05744_ ;
 wire \reg_module/_05745_ ;
 wire \reg_module/_05746_ ;
 wire \reg_module/_05747_ ;
 wire \reg_module/_05748_ ;
 wire \reg_module/_05749_ ;
 wire \reg_module/_05750_ ;
 wire \reg_module/_05751_ ;
 wire \reg_module/_05752_ ;
 wire \reg_module/_05753_ ;
 wire \reg_module/_05754_ ;
 wire \reg_module/_05755_ ;
 wire \reg_module/_05756_ ;
 wire \reg_module/_05757_ ;
 wire \reg_module/_05758_ ;
 wire \reg_module/_05759_ ;
 wire \reg_module/_05760_ ;
 wire \reg_module/_05761_ ;
 wire \reg_module/_05762_ ;
 wire \reg_module/_05763_ ;
 wire \reg_module/_05764_ ;
 wire \reg_module/_05765_ ;
 wire \reg_module/_05766_ ;
 wire \reg_module/_05767_ ;
 wire \reg_module/_05768_ ;
 wire \reg_module/_05769_ ;
 wire \reg_module/_05770_ ;
 wire \reg_module/_05771_ ;
 wire \reg_module/_05772_ ;
 wire \reg_module/_05773_ ;
 wire \reg_module/_05774_ ;
 wire \reg_module/_05775_ ;
 wire \reg_module/_05776_ ;
 wire \reg_module/_05777_ ;
 wire \reg_module/_05778_ ;
 wire \reg_module/_05779_ ;
 wire \reg_module/_05780_ ;
 wire \reg_module/_05781_ ;
 wire \reg_module/_05782_ ;
 wire \reg_module/_05783_ ;
 wire \reg_module/_05784_ ;
 wire \reg_module/_05785_ ;
 wire \reg_module/_05786_ ;
 wire \reg_module/_05787_ ;
 wire \reg_module/_05788_ ;
 wire \reg_module/_05789_ ;
 wire \reg_module/_05790_ ;
 wire \reg_module/_05791_ ;
 wire \reg_module/_05792_ ;
 wire \reg_module/_05793_ ;
 wire \reg_module/_05794_ ;
 wire \reg_module/_05795_ ;
 wire \reg_module/_05796_ ;
 wire \reg_module/_05797_ ;
 wire \reg_module/_05798_ ;
 wire \reg_module/_05799_ ;
 wire \reg_module/_05800_ ;
 wire \reg_module/_05801_ ;
 wire \reg_module/_05802_ ;
 wire \reg_module/_05803_ ;
 wire \reg_module/_05804_ ;
 wire \reg_module/_05805_ ;
 wire \reg_module/_05806_ ;
 wire \reg_module/_05807_ ;
 wire \reg_module/_05808_ ;
 wire \reg_module/_05809_ ;
 wire \reg_module/_05810_ ;
 wire \reg_module/_05811_ ;
 wire \reg_module/_05812_ ;
 wire \reg_module/_05813_ ;
 wire \reg_module/_05814_ ;
 wire \reg_module/_05815_ ;
 wire \reg_module/_05816_ ;
 wire \reg_module/_05817_ ;
 wire \reg_module/_05818_ ;
 wire \reg_module/_05819_ ;
 wire \reg_module/_05820_ ;
 wire \reg_module/_05821_ ;
 wire \reg_module/_05822_ ;
 wire \reg_module/_05823_ ;
 wire \reg_module/_05824_ ;
 wire \reg_module/_05825_ ;
 wire \reg_module/_05826_ ;
 wire \reg_module/_05827_ ;
 wire \reg_module/_05828_ ;
 wire \reg_module/_05829_ ;
 wire \reg_module/_05830_ ;
 wire \reg_module/_05831_ ;
 wire \reg_module/_05832_ ;
 wire \reg_module/_05833_ ;
 wire \reg_module/_05834_ ;
 wire \reg_module/_05835_ ;
 wire \reg_module/_05836_ ;
 wire \reg_module/_05837_ ;
 wire \reg_module/_05838_ ;
 wire \reg_module/_05839_ ;
 wire \reg_module/_05840_ ;
 wire \reg_module/_05841_ ;
 wire \reg_module/_05842_ ;
 wire \reg_module/_05843_ ;
 wire \reg_module/_05844_ ;
 wire \reg_module/_05845_ ;
 wire \reg_module/_05846_ ;
 wire \reg_module/_05847_ ;
 wire \reg_module/_05848_ ;
 wire \reg_module/_05849_ ;
 wire \reg_module/_05850_ ;
 wire \reg_module/_05851_ ;
 wire \reg_module/_05852_ ;
 wire \reg_module/_05853_ ;
 wire \reg_module/_05854_ ;
 wire \reg_module/_05855_ ;
 wire \reg_module/_05856_ ;
 wire \reg_module/_05857_ ;
 wire \reg_module/_05858_ ;
 wire \reg_module/_05859_ ;
 wire \reg_module/_05860_ ;
 wire \reg_module/_05861_ ;
 wire \reg_module/_05862_ ;
 wire \reg_module/_05863_ ;
 wire \reg_module/_05864_ ;
 wire \reg_module/_05865_ ;
 wire \reg_module/_05866_ ;
 wire \reg_module/_05867_ ;
 wire \reg_module/_05868_ ;
 wire \reg_module/_05869_ ;
 wire \reg_module/_05870_ ;
 wire \reg_module/_05871_ ;
 wire \reg_module/_05872_ ;
 wire \reg_module/_05873_ ;
 wire \reg_module/_05874_ ;
 wire \reg_module/_05875_ ;
 wire \reg_module/_05876_ ;
 wire \reg_module/_05877_ ;
 wire \reg_module/_05878_ ;
 wire \reg_module/_05879_ ;
 wire \reg_module/_05880_ ;
 wire \reg_module/_05881_ ;
 wire \reg_module/_05882_ ;
 wire \reg_module/_05883_ ;
 wire \reg_module/_05884_ ;
 wire \reg_module/_05885_ ;
 wire \reg_module/_05886_ ;
 wire \reg_module/_05887_ ;
 wire \reg_module/_05888_ ;
 wire \reg_module/_05889_ ;
 wire \reg_module/_05890_ ;
 wire \reg_module/_05891_ ;
 wire \reg_module/_05892_ ;
 wire \reg_module/_05893_ ;
 wire \reg_module/_05894_ ;
 wire \reg_module/_05895_ ;
 wire \reg_module/_05896_ ;
 wire \reg_module/_05897_ ;
 wire \reg_module/_05898_ ;
 wire \reg_module/_05899_ ;
 wire \reg_module/_05900_ ;
 wire \reg_module/_05901_ ;
 wire \reg_module/_05902_ ;
 wire \reg_module/_05903_ ;
 wire \reg_module/_05904_ ;
 wire \reg_module/_05905_ ;
 wire \reg_module/_05906_ ;
 wire \reg_module/_05907_ ;
 wire \reg_module/_05908_ ;
 wire \reg_module/_05909_ ;
 wire \reg_module/_05910_ ;
 wire \reg_module/_05911_ ;
 wire \reg_module/_05912_ ;
 wire \reg_module/_05913_ ;
 wire \reg_module/_05914_ ;
 wire \reg_module/_05915_ ;
 wire \reg_module/_05916_ ;
 wire \reg_module/_05917_ ;
 wire \reg_module/_05918_ ;
 wire \reg_module/_05919_ ;
 wire \reg_module/_05920_ ;
 wire \reg_module/_05921_ ;
 wire \reg_module/_05922_ ;
 wire \reg_module/_05923_ ;
 wire \reg_module/_05924_ ;
 wire \reg_module/_05925_ ;
 wire \reg_module/_05926_ ;
 wire \reg_module/_05927_ ;
 wire \reg_module/_05928_ ;
 wire \reg_module/_05929_ ;
 wire \reg_module/_05930_ ;
 wire \reg_module/_05931_ ;
 wire \reg_module/_05932_ ;
 wire \reg_module/_05933_ ;
 wire \reg_module/_05934_ ;
 wire \reg_module/_05935_ ;
 wire \reg_module/_05936_ ;
 wire \reg_module/_05937_ ;
 wire \reg_module/_05938_ ;
 wire \reg_module/_05939_ ;
 wire \reg_module/_05940_ ;
 wire \reg_module/_05941_ ;
 wire \reg_module/_05942_ ;
 wire \reg_module/_05943_ ;
 wire \reg_module/_05944_ ;
 wire \reg_module/_05945_ ;
 wire \reg_module/_05946_ ;
 wire \reg_module/_05947_ ;
 wire \reg_module/_05948_ ;
 wire \reg_module/_05949_ ;
 wire \reg_module/_05950_ ;
 wire \reg_module/_05951_ ;
 wire \reg_module/_05952_ ;
 wire \reg_module/_05953_ ;
 wire \reg_module/_05954_ ;
 wire \reg_module/_05955_ ;
 wire \reg_module/_05956_ ;
 wire \reg_module/_05957_ ;
 wire \reg_module/_05958_ ;
 wire \reg_module/_05959_ ;
 wire \reg_module/_05960_ ;
 wire \reg_module/_05961_ ;
 wire \reg_module/_05962_ ;
 wire \reg_module/_05963_ ;
 wire \reg_module/_05964_ ;
 wire \reg_module/_05965_ ;
 wire \reg_module/_05966_ ;
 wire \reg_module/_05967_ ;
 wire \reg_module/_05968_ ;
 wire \reg_module/_05969_ ;
 wire \reg_module/_05970_ ;
 wire \reg_module/_05971_ ;
 wire \reg_module/_05972_ ;
 wire \reg_module/_05973_ ;
 wire \reg_module/_05974_ ;
 wire \reg_module/_05975_ ;
 wire \reg_module/_05976_ ;
 wire \reg_module/_05977_ ;
 wire \reg_module/_05978_ ;
 wire \reg_module/_05979_ ;
 wire \reg_module/_05980_ ;
 wire \reg_module/_05981_ ;
 wire \reg_module/_05982_ ;
 wire \reg_module/_05983_ ;
 wire \reg_module/_05984_ ;
 wire \reg_module/_05985_ ;
 wire \reg_module/_05986_ ;
 wire \reg_module/_05987_ ;
 wire \reg_module/_05988_ ;
 wire \reg_module/_05989_ ;
 wire \reg_module/_05990_ ;
 wire \reg_module/_05991_ ;
 wire \reg_module/_05992_ ;
 wire \reg_module/_05993_ ;
 wire \reg_module/_05994_ ;
 wire \reg_module/_05995_ ;
 wire \reg_module/_05996_ ;
 wire \reg_module/_05997_ ;
 wire \reg_module/_05998_ ;
 wire \reg_module/_05999_ ;
 wire \reg_module/_06000_ ;
 wire \reg_module/_06001_ ;
 wire \reg_module/_06002_ ;
 wire \reg_module/_06003_ ;
 wire \reg_module/_06004_ ;
 wire \reg_module/_06005_ ;
 wire \reg_module/_06006_ ;
 wire \reg_module/_06007_ ;
 wire \reg_module/_06008_ ;
 wire \reg_module/_06009_ ;
 wire \reg_module/_06010_ ;
 wire \reg_module/_06011_ ;
 wire \reg_module/_06012_ ;
 wire \reg_module/_06013_ ;
 wire \reg_module/_06014_ ;
 wire \reg_module/_06015_ ;
 wire \reg_module/_06016_ ;
 wire \reg_module/_06017_ ;
 wire \reg_module/_06018_ ;
 wire \reg_module/_06019_ ;
 wire \reg_module/_06020_ ;
 wire \reg_module/_06021_ ;
 wire \reg_module/_06022_ ;
 wire \reg_module/_06023_ ;
 wire \reg_module/_06024_ ;
 wire \reg_module/_06025_ ;
 wire \reg_module/_06026_ ;
 wire \reg_module/_06027_ ;
 wire \reg_module/_06028_ ;
 wire \reg_module/_06029_ ;
 wire \reg_module/_06030_ ;
 wire \reg_module/_06031_ ;
 wire \reg_module/_06032_ ;
 wire \reg_module/_06033_ ;
 wire \reg_module/_06034_ ;
 wire \reg_module/_06035_ ;
 wire \reg_module/_06036_ ;
 wire \reg_module/_06037_ ;
 wire \reg_module/_06038_ ;
 wire \reg_module/_06039_ ;
 wire \reg_module/_06040_ ;
 wire \reg_module/_06041_ ;
 wire \reg_module/_06042_ ;
 wire \reg_module/_06043_ ;
 wire \reg_module/_06044_ ;
 wire \reg_module/_06045_ ;
 wire \reg_module/_06046_ ;
 wire \reg_module/_06047_ ;
 wire \reg_module/_06048_ ;
 wire \reg_module/_06049_ ;
 wire \reg_module/_06050_ ;
 wire \reg_module/_06051_ ;
 wire \reg_module/_06052_ ;
 wire \reg_module/_06053_ ;
 wire \reg_module/_06054_ ;
 wire \reg_module/_06055_ ;
 wire \reg_module/_06056_ ;
 wire \reg_module/_06057_ ;
 wire \reg_module/_06058_ ;
 wire \reg_module/_06059_ ;
 wire \reg_module/_06060_ ;
 wire \reg_module/_06061_ ;
 wire \reg_module/_06062_ ;
 wire \reg_module/_06063_ ;
 wire \reg_module/_06064_ ;
 wire \reg_module/_06065_ ;
 wire \reg_module/_06066_ ;
 wire \reg_module/_06067_ ;
 wire \reg_module/_06068_ ;
 wire \reg_module/_06069_ ;
 wire \reg_module/_06070_ ;
 wire \reg_module/_06071_ ;
 wire \reg_module/_06072_ ;
 wire \reg_module/_06073_ ;
 wire \reg_module/_06074_ ;
 wire \reg_module/_06075_ ;
 wire \reg_module/_06076_ ;
 wire \reg_module/_06077_ ;
 wire \reg_module/_06078_ ;
 wire \reg_module/_06079_ ;
 wire \reg_module/_06080_ ;
 wire \reg_module/_06081_ ;
 wire \reg_module/_06082_ ;
 wire \reg_module/_06083_ ;
 wire \reg_module/_06084_ ;
 wire \reg_module/_06085_ ;
 wire \reg_module/_06086_ ;
 wire \reg_module/_06087_ ;
 wire \reg_module/_06088_ ;
 wire \reg_module/_06089_ ;
 wire \reg_module/_06090_ ;
 wire \reg_module/_06091_ ;
 wire \reg_module/_06092_ ;
 wire \reg_module/_06093_ ;
 wire \reg_module/_06094_ ;
 wire \reg_module/_06095_ ;
 wire \reg_module/_06096_ ;
 wire \reg_module/_06097_ ;
 wire \reg_module/_06098_ ;
 wire \reg_module/_06099_ ;
 wire \reg_module/_06100_ ;
 wire \reg_module/_06101_ ;
 wire \reg_module/_06102_ ;
 wire \reg_module/_06103_ ;
 wire \reg_module/_06104_ ;
 wire \reg_module/_06105_ ;
 wire \reg_module/_06106_ ;
 wire \reg_module/_06107_ ;
 wire \reg_module/_06108_ ;
 wire \reg_module/_06109_ ;
 wire \reg_module/_06110_ ;
 wire \reg_module/_06111_ ;
 wire \reg_module/_06112_ ;
 wire \reg_module/_06113_ ;
 wire \reg_module/_06114_ ;
 wire \reg_module/_06115_ ;
 wire \reg_module/_06116_ ;
 wire \reg_module/_06117_ ;
 wire \reg_module/_06118_ ;
 wire \reg_module/_06119_ ;
 wire \reg_module/_06120_ ;
 wire \reg_module/_06121_ ;
 wire \reg_module/_06122_ ;
 wire \reg_module/_06123_ ;
 wire \reg_module/_06124_ ;
 wire \reg_module/_06125_ ;
 wire \reg_module/_06126_ ;
 wire \reg_module/_06127_ ;
 wire \reg_module/_06128_ ;
 wire \reg_module/_06129_ ;
 wire \reg_module/_06130_ ;
 wire \reg_module/_06131_ ;
 wire \reg_module/_06132_ ;
 wire \reg_module/_06133_ ;
 wire \reg_module/_06134_ ;
 wire \reg_module/_06135_ ;
 wire \reg_module/_06136_ ;
 wire \reg_module/_06137_ ;
 wire \reg_module/_06138_ ;
 wire \reg_module/_06139_ ;
 wire \reg_module/_06140_ ;
 wire \reg_module/_06141_ ;
 wire \reg_module/_06142_ ;
 wire \reg_module/_06143_ ;
 wire \reg_module/_06144_ ;
 wire \reg_module/_06145_ ;
 wire \reg_module/_06146_ ;
 wire \reg_module/_06147_ ;
 wire \reg_module/_06148_ ;
 wire \reg_module/_06149_ ;
 wire \reg_module/_06150_ ;
 wire \reg_module/_06151_ ;
 wire \reg_module/_06152_ ;
 wire \reg_module/_06153_ ;
 wire \reg_module/_06154_ ;
 wire \reg_module/_06155_ ;
 wire \reg_module/_06156_ ;
 wire \reg_module/_06157_ ;
 wire \reg_module/_06158_ ;
 wire \reg_module/_06159_ ;
 wire \reg_module/_06160_ ;
 wire \reg_module/_06161_ ;
 wire \reg_module/_06162_ ;
 wire \reg_module/_06163_ ;
 wire \reg_module/_06164_ ;
 wire \reg_module/_06165_ ;
 wire \reg_module/_06166_ ;
 wire \reg_module/_06167_ ;
 wire \reg_module/_06168_ ;
 wire \reg_module/_06169_ ;
 wire \reg_module/_06170_ ;
 wire \reg_module/_06171_ ;
 wire \reg_module/_06172_ ;
 wire \reg_module/_06173_ ;
 wire \reg_module/_06174_ ;
 wire \reg_module/_06175_ ;
 wire \reg_module/_06176_ ;
 wire \reg_module/_06177_ ;
 wire \reg_module/_06178_ ;
 wire \reg_module/_06179_ ;
 wire \reg_module/_06180_ ;
 wire \reg_module/_06181_ ;
 wire \reg_module/_06182_ ;
 wire \reg_module/_06183_ ;
 wire \reg_module/_06184_ ;
 wire \reg_module/_06185_ ;
 wire \reg_module/_06186_ ;
 wire \reg_module/_06187_ ;
 wire \reg_module/_06188_ ;
 wire \reg_module/_06189_ ;
 wire \reg_module/_06190_ ;
 wire \reg_module/_06191_ ;
 wire \reg_module/_06192_ ;
 wire \reg_module/_06193_ ;
 wire \reg_module/_06194_ ;
 wire \reg_module/_06195_ ;
 wire \reg_module/_06196_ ;
 wire \reg_module/_06197_ ;
 wire \reg_module/_06198_ ;
 wire \reg_module/_06199_ ;
 wire \reg_module/_06200_ ;
 wire \reg_module/_06201_ ;
 wire \reg_module/_06202_ ;
 wire \reg_module/_06203_ ;
 wire \reg_module/_06204_ ;
 wire \reg_module/_06205_ ;
 wire \reg_module/_06206_ ;
 wire \reg_module/_06207_ ;
 wire \reg_module/_06208_ ;
 wire \reg_module/_06209_ ;
 wire \reg_module/_06210_ ;
 wire \reg_module/_06211_ ;
 wire \reg_module/_06212_ ;
 wire \reg_module/_06213_ ;
 wire \reg_module/_06214_ ;
 wire \reg_module/_06215_ ;
 wire \reg_module/_06216_ ;
 wire \reg_module/_06217_ ;
 wire \reg_module/_06218_ ;
 wire \reg_module/_06219_ ;
 wire \reg_module/_06220_ ;
 wire \reg_module/_06221_ ;
 wire \reg_module/_06222_ ;
 wire \reg_module/_06223_ ;
 wire \reg_module/_06224_ ;
 wire \reg_module/_06225_ ;
 wire \reg_module/_06226_ ;
 wire \reg_module/_06227_ ;
 wire \reg_module/_06228_ ;
 wire \reg_module/_06229_ ;
 wire \reg_module/_06230_ ;
 wire \reg_module/_06231_ ;
 wire \reg_module/_06232_ ;
 wire \reg_module/_06233_ ;
 wire \reg_module/_06234_ ;
 wire \reg_module/_06235_ ;
 wire \reg_module/_06236_ ;
 wire \reg_module/_06237_ ;
 wire \reg_module/_06238_ ;
 wire \reg_module/_06239_ ;
 wire \reg_module/_06240_ ;
 wire \reg_module/_06241_ ;
 wire \reg_module/_06242_ ;
 wire \reg_module/_06243_ ;
 wire \reg_module/_06244_ ;
 wire \reg_module/_06245_ ;
 wire \reg_module/_06246_ ;
 wire \reg_module/_06247_ ;
 wire \reg_module/_06248_ ;
 wire \reg_module/_06249_ ;
 wire \reg_module/_06250_ ;
 wire \reg_module/_06251_ ;
 wire \reg_module/_06252_ ;
 wire \reg_module/_06253_ ;
 wire \reg_module/_06254_ ;
 wire \reg_module/_06255_ ;
 wire \reg_module/_06256_ ;
 wire \reg_module/_06257_ ;
 wire \reg_module/_06258_ ;
 wire \reg_module/_06259_ ;
 wire \reg_module/_06260_ ;
 wire \reg_module/_06261_ ;
 wire \reg_module/_06262_ ;
 wire \reg_module/_06263_ ;
 wire \reg_module/_06264_ ;
 wire \reg_module/_06265_ ;
 wire \reg_module/_06266_ ;
 wire \reg_module/_06267_ ;
 wire \reg_module/_06268_ ;
 wire \reg_module/_06269_ ;
 wire \reg_module/_06270_ ;
 wire \reg_module/_06271_ ;
 wire \reg_module/_06272_ ;
 wire \reg_module/_06273_ ;
 wire \reg_module/_06274_ ;
 wire \reg_module/_06275_ ;
 wire \reg_module/_06276_ ;
 wire \reg_module/_06277_ ;
 wire \reg_module/_06278_ ;
 wire \reg_module/_06279_ ;
 wire \reg_module/_06280_ ;
 wire \reg_module/_06281_ ;
 wire \reg_module/_06282_ ;
 wire \reg_module/_06283_ ;
 wire \reg_module/_06284_ ;
 wire \reg_module/_06285_ ;
 wire \reg_module/_06286_ ;
 wire \reg_module/_06287_ ;
 wire \reg_module/_06288_ ;
 wire \reg_module/_06289_ ;
 wire \reg_module/_06290_ ;
 wire \reg_module/_06291_ ;
 wire \reg_module/_06292_ ;
 wire \reg_module/_06293_ ;
 wire \reg_module/_06294_ ;
 wire \reg_module/_06295_ ;
 wire \reg_module/_06296_ ;
 wire \reg_module/_06297_ ;
 wire \reg_module/_06298_ ;
 wire \reg_module/_06299_ ;
 wire \reg_module/_06300_ ;
 wire \reg_module/_06301_ ;
 wire \reg_module/_06302_ ;
 wire \reg_module/_06303_ ;
 wire \reg_module/_06304_ ;
 wire \reg_module/_06305_ ;
 wire \reg_module/_06306_ ;
 wire \reg_module/_06307_ ;
 wire \reg_module/_06308_ ;
 wire \reg_module/_06309_ ;
 wire \reg_module/_06310_ ;
 wire \reg_module/_06311_ ;
 wire \reg_module/_06312_ ;
 wire \reg_module/_06313_ ;
 wire \reg_module/_06314_ ;
 wire \reg_module/_06315_ ;
 wire \reg_module/_06316_ ;
 wire \reg_module/_06317_ ;
 wire \reg_module/_06318_ ;
 wire \reg_module/_06319_ ;
 wire \reg_module/_06320_ ;
 wire \reg_module/_06321_ ;
 wire \reg_module/_06322_ ;
 wire \reg_module/_06323_ ;
 wire \reg_module/_06324_ ;
 wire \reg_module/_06325_ ;
 wire \reg_module/_06326_ ;
 wire \reg_module/_06327_ ;
 wire \reg_module/_06328_ ;
 wire \reg_module/_06329_ ;
 wire \reg_module/_06330_ ;
 wire \reg_module/_06331_ ;
 wire \reg_module/_06332_ ;
 wire \reg_module/_06333_ ;
 wire \reg_module/_06334_ ;
 wire \reg_module/_06335_ ;
 wire \reg_module/_06336_ ;
 wire \reg_module/_06337_ ;
 wire \reg_module/_06338_ ;
 wire \reg_module/_06339_ ;
 wire \reg_module/_06340_ ;
 wire \reg_module/_06341_ ;
 wire \reg_module/_06342_ ;
 wire \reg_module/_06343_ ;
 wire \reg_module/_06344_ ;
 wire \reg_module/_06345_ ;
 wire \reg_module/_06346_ ;
 wire \reg_module/_06347_ ;
 wire \reg_module/_06348_ ;
 wire \reg_module/_06349_ ;
 wire \reg_module/_06350_ ;
 wire \reg_module/_06351_ ;
 wire \reg_module/_06352_ ;
 wire \reg_module/_06353_ ;
 wire \reg_module/_06354_ ;
 wire \reg_module/_06355_ ;
 wire \reg_module/_06356_ ;
 wire \reg_module/_06357_ ;
 wire \reg_module/_06358_ ;
 wire \reg_module/_06359_ ;
 wire \reg_module/_06360_ ;
 wire \reg_module/_06361_ ;
 wire \reg_module/_06362_ ;
 wire \reg_module/_06363_ ;
 wire \reg_module/_06364_ ;
 wire \reg_module/_06365_ ;
 wire \reg_module/_06366_ ;
 wire \reg_module/_06367_ ;
 wire \reg_module/_06368_ ;
 wire \reg_module/_06369_ ;
 wire \reg_module/_06370_ ;
 wire \reg_module/_06371_ ;
 wire \reg_module/_06372_ ;
 wire \reg_module/_06373_ ;
 wire \reg_module/_06374_ ;
 wire \reg_module/_06375_ ;
 wire \reg_module/_06376_ ;
 wire \reg_module/_06377_ ;
 wire \reg_module/_06378_ ;
 wire \reg_module/_06379_ ;
 wire \reg_module/_06380_ ;
 wire \reg_module/_06381_ ;
 wire \reg_module/_06382_ ;
 wire \reg_module/_06383_ ;
 wire \reg_module/_06384_ ;
 wire \reg_module/_06385_ ;
 wire \reg_module/_06386_ ;
 wire \reg_module/_06387_ ;
 wire \reg_module/_06388_ ;
 wire \reg_module/_06389_ ;
 wire \reg_module/_06390_ ;
 wire \reg_module/_06391_ ;
 wire \reg_module/_06392_ ;
 wire \reg_module/_06393_ ;
 wire \reg_module/_06394_ ;
 wire \reg_module/_06395_ ;
 wire \reg_module/_06396_ ;
 wire \reg_module/_06397_ ;
 wire \reg_module/_06398_ ;
 wire \reg_module/_06399_ ;
 wire \reg_module/_06400_ ;
 wire \reg_module/_06401_ ;
 wire \reg_module/_06402_ ;
 wire \reg_module/_06403_ ;
 wire \reg_module/_06404_ ;
 wire \reg_module/_06405_ ;
 wire \reg_module/_06406_ ;
 wire \reg_module/_06407_ ;
 wire \reg_module/_06408_ ;
 wire \reg_module/_06409_ ;
 wire \reg_module/_06410_ ;
 wire \reg_module/_06411_ ;
 wire \reg_module/_06412_ ;
 wire \reg_module/_06413_ ;
 wire \reg_module/_06414_ ;
 wire \reg_module/_06415_ ;
 wire \reg_module/_06416_ ;
 wire \reg_module/_06417_ ;
 wire \reg_module/_06418_ ;
 wire \reg_module/_06419_ ;
 wire \reg_module/_06420_ ;
 wire \reg_module/_06421_ ;
 wire \reg_module/_06422_ ;
 wire \reg_module/_06423_ ;
 wire \reg_module/_06424_ ;
 wire \reg_module/_06425_ ;
 wire \reg_module/_06426_ ;
 wire \reg_module/_06427_ ;
 wire \reg_module/_06428_ ;
 wire \reg_module/_06429_ ;
 wire \reg_module/_06430_ ;
 wire \reg_module/_06431_ ;
 wire \reg_module/_06432_ ;
 wire \reg_module/_06433_ ;
 wire \reg_module/_06434_ ;
 wire \reg_module/_06435_ ;
 wire \reg_module/_06436_ ;
 wire \reg_module/_06437_ ;
 wire \reg_module/_06438_ ;
 wire \reg_module/_06439_ ;
 wire \reg_module/_06440_ ;
 wire \reg_module/_06441_ ;
 wire \reg_module/_06442_ ;
 wire \reg_module/_06443_ ;
 wire \reg_module/_06444_ ;
 wire \reg_module/_06445_ ;
 wire \reg_module/_06446_ ;
 wire \reg_module/_06447_ ;
 wire \reg_module/_06448_ ;
 wire \reg_module/_06449_ ;
 wire \reg_module/_06450_ ;
 wire \reg_module/_06451_ ;
 wire \reg_module/_06452_ ;
 wire \reg_module/_06453_ ;
 wire \reg_module/_06454_ ;
 wire \reg_module/_06455_ ;
 wire \reg_module/_06456_ ;
 wire \reg_module/_06457_ ;
 wire \reg_module/_06458_ ;
 wire \reg_module/_06459_ ;
 wire \reg_module/_06460_ ;
 wire \reg_module/_06461_ ;
 wire \reg_module/_06462_ ;
 wire \reg_module/_06463_ ;
 wire \reg_module/_06464_ ;
 wire \reg_module/_06465_ ;
 wire \reg_module/_06466_ ;
 wire \reg_module/_06467_ ;
 wire \reg_module/_06468_ ;
 wire \reg_module/_06469_ ;
 wire \reg_module/_06470_ ;
 wire \reg_module/_06471_ ;
 wire \reg_module/_06472_ ;
 wire \reg_module/_06473_ ;
 wire \reg_module/_06474_ ;
 wire \reg_module/_06475_ ;
 wire \reg_module/_06476_ ;
 wire \reg_module/_06477_ ;
 wire \reg_module/_06478_ ;
 wire \reg_module/_06479_ ;
 wire \reg_module/_06480_ ;
 wire \reg_module/_06481_ ;
 wire \reg_module/_06482_ ;
 wire \reg_module/_06483_ ;
 wire \reg_module/_06484_ ;
 wire \reg_module/_06485_ ;
 wire \reg_module/_06486_ ;
 wire \reg_module/_06487_ ;
 wire \reg_module/_06488_ ;
 wire \reg_module/_06489_ ;
 wire \reg_module/_06490_ ;
 wire \reg_module/_06491_ ;
 wire \reg_module/_06492_ ;
 wire \reg_module/_06493_ ;
 wire \reg_module/_06494_ ;
 wire \reg_module/_06495_ ;
 wire \reg_module/_06496_ ;
 wire \reg_module/_06497_ ;
 wire \reg_module/_06498_ ;
 wire \reg_module/_06499_ ;
 wire \reg_module/_06500_ ;
 wire \reg_module/_06501_ ;
 wire \reg_module/_06502_ ;
 wire \reg_module/_06503_ ;
 wire \reg_module/_06504_ ;
 wire \reg_module/_06505_ ;
 wire \reg_module/_06506_ ;
 wire \reg_module/_06507_ ;
 wire \reg_module/_06508_ ;
 wire \reg_module/_06509_ ;
 wire \reg_module/_06510_ ;
 wire \reg_module/_06511_ ;
 wire \reg_module/_06512_ ;
 wire \reg_module/_06513_ ;
 wire \reg_module/_06514_ ;
 wire \reg_module/_06515_ ;
 wire \reg_module/_06516_ ;
 wire \reg_module/_06517_ ;
 wire \reg_module/_06518_ ;
 wire \reg_module/_06519_ ;
 wire \reg_module/_06520_ ;
 wire \reg_module/_06521_ ;
 wire \reg_module/_06522_ ;
 wire \reg_module/_06523_ ;
 wire \reg_module/_06524_ ;
 wire \reg_module/_06525_ ;
 wire \reg_module/_06526_ ;
 wire \reg_module/_06527_ ;
 wire \reg_module/_06528_ ;
 wire \reg_module/_06529_ ;
 wire \reg_module/_06530_ ;
 wire \reg_module/_06531_ ;
 wire \reg_module/_06532_ ;
 wire \reg_module/_06533_ ;
 wire \reg_module/_06534_ ;
 wire \reg_module/_06535_ ;
 wire \reg_module/_06536_ ;
 wire \reg_module/_06537_ ;
 wire \reg_module/_06538_ ;
 wire \reg_module/_06539_ ;
 wire \reg_module/_06540_ ;
 wire \reg_module/_06541_ ;
 wire \reg_module/_06542_ ;
 wire \reg_module/_06543_ ;
 wire \reg_module/_06544_ ;
 wire \reg_module/_06545_ ;
 wire \reg_module/_06546_ ;
 wire \reg_module/_06547_ ;
 wire \reg_module/_06548_ ;
 wire \reg_module/_06549_ ;
 wire \reg_module/_06550_ ;
 wire \reg_module/_06551_ ;
 wire \reg_module/_06552_ ;
 wire \reg_module/_06553_ ;
 wire \reg_module/_06554_ ;
 wire \reg_module/_06555_ ;
 wire \reg_module/_06556_ ;
 wire \reg_module/_06557_ ;
 wire \reg_module/_06558_ ;
 wire \reg_module/_06559_ ;
 wire \reg_module/_06560_ ;
 wire \reg_module/_06561_ ;
 wire \reg_module/_06562_ ;
 wire \reg_module/_06563_ ;
 wire \reg_module/_06564_ ;
 wire \reg_module/_06565_ ;
 wire \reg_module/_06566_ ;
 wire \reg_module/_06567_ ;
 wire \reg_module/_06568_ ;
 wire \reg_module/_06569_ ;
 wire \reg_module/_06570_ ;
 wire \reg_module/_06571_ ;
 wire \reg_module/_06572_ ;
 wire \reg_module/_06573_ ;
 wire \reg_module/_06574_ ;
 wire \reg_module/_06575_ ;
 wire \reg_module/_06576_ ;
 wire \reg_module/_06577_ ;
 wire \reg_module/_06578_ ;
 wire \reg_module/_06579_ ;
 wire \reg_module/_06580_ ;
 wire \reg_module/_06581_ ;
 wire \reg_module/_06582_ ;
 wire \reg_module/_06583_ ;
 wire \reg_module/_06584_ ;
 wire \reg_module/_06585_ ;
 wire \reg_module/_06586_ ;
 wire \reg_module/_06587_ ;
 wire \reg_module/_06588_ ;
 wire \reg_module/_06589_ ;
 wire \reg_module/_06590_ ;
 wire \reg_module/_06591_ ;
 wire \reg_module/_06592_ ;
 wire \reg_module/_06593_ ;
 wire \reg_module/_06594_ ;
 wire \reg_module/_06595_ ;
 wire \reg_module/_06596_ ;
 wire \reg_module/_06597_ ;
 wire \reg_module/_06598_ ;
 wire \reg_module/_06599_ ;
 wire \reg_module/_06600_ ;
 wire \reg_module/_06601_ ;
 wire \reg_module/_06602_ ;
 wire \reg_module/_06603_ ;
 wire \reg_module/_06604_ ;
 wire \reg_module/_06605_ ;
 wire \reg_module/_06606_ ;
 wire \reg_module/_06607_ ;
 wire \reg_module/_06608_ ;
 wire \reg_module/_06609_ ;
 wire \reg_module/_06610_ ;
 wire \reg_module/_06611_ ;
 wire \reg_module/_06612_ ;
 wire \reg_module/_06613_ ;
 wire \reg_module/_06614_ ;
 wire \reg_module/_06615_ ;
 wire \reg_module/_06616_ ;
 wire \reg_module/_06617_ ;
 wire \reg_module/_06618_ ;
 wire \reg_module/_06619_ ;
 wire \reg_module/_06620_ ;
 wire \reg_module/_06621_ ;
 wire \reg_module/_06622_ ;
 wire \reg_module/_06623_ ;
 wire \reg_module/_06624_ ;
 wire \reg_module/_06625_ ;
 wire \reg_module/_06626_ ;
 wire \reg_module/_06627_ ;
 wire \reg_module/_06628_ ;
 wire \reg_module/_06629_ ;
 wire \reg_module/_06630_ ;
 wire \reg_module/_06631_ ;
 wire \reg_module/_06632_ ;
 wire \reg_module/_06633_ ;
 wire \reg_module/_06634_ ;
 wire \reg_module/_06635_ ;
 wire \reg_module/_06636_ ;
 wire \reg_module/_06637_ ;
 wire \reg_module/_06638_ ;
 wire \reg_module/_06639_ ;
 wire \reg_module/_06640_ ;
 wire \reg_module/_06641_ ;
 wire \reg_module/_06642_ ;
 wire \reg_module/_06643_ ;
 wire \reg_module/_06644_ ;
 wire \reg_module/_06645_ ;
 wire \reg_module/_06646_ ;
 wire \reg_module/_06647_ ;
 wire \reg_module/_06648_ ;
 wire \reg_module/_06649_ ;
 wire \reg_module/_06650_ ;
 wire \reg_module/_06651_ ;
 wire \reg_module/_06652_ ;
 wire \reg_module/_06653_ ;
 wire \reg_module/_06654_ ;
 wire \reg_module/_06655_ ;
 wire \reg_module/_06656_ ;
 wire \reg_module/_06657_ ;
 wire \reg_module/_06658_ ;
 wire \reg_module/_06659_ ;
 wire \reg_module/_06660_ ;
 wire \reg_module/_06661_ ;
 wire \reg_module/_06662_ ;
 wire \reg_module/_06663_ ;
 wire \reg_module/_06664_ ;
 wire \reg_module/_06665_ ;
 wire \reg_module/_06666_ ;
 wire \reg_module/_06667_ ;
 wire \reg_module/_06668_ ;
 wire \reg_module/_06669_ ;
 wire \reg_module/_06670_ ;
 wire \reg_module/_06671_ ;
 wire \reg_module/_06672_ ;
 wire \reg_module/_06673_ ;
 wire \reg_module/_06674_ ;
 wire \reg_module/_06675_ ;
 wire \reg_module/_06676_ ;
 wire \reg_module/_06677_ ;
 wire \reg_module/_06678_ ;
 wire \reg_module/_06679_ ;
 wire \reg_module/_06680_ ;
 wire \reg_module/_06681_ ;
 wire \reg_module/_06682_ ;
 wire \reg_module/_06683_ ;
 wire \reg_module/_06684_ ;
 wire \reg_module/_06685_ ;
 wire \reg_module/_06686_ ;
 wire \reg_module/_06687_ ;
 wire \reg_module/_06688_ ;
 wire \reg_module/_06689_ ;
 wire \reg_module/_06690_ ;
 wire \reg_module/_06691_ ;
 wire \reg_module/_06692_ ;
 wire \reg_module/_06693_ ;
 wire \reg_module/_06694_ ;
 wire \reg_module/_06695_ ;
 wire \reg_module/_06696_ ;
 wire \reg_module/_06697_ ;
 wire \reg_module/_06698_ ;
 wire \reg_module/_06699_ ;
 wire \reg_module/_06700_ ;
 wire \reg_module/_06701_ ;
 wire \reg_module/_06702_ ;
 wire \reg_module/_06703_ ;
 wire \reg_module/_06704_ ;
 wire \reg_module/_06705_ ;
 wire \reg_module/_06706_ ;
 wire \reg_module/_06707_ ;
 wire \reg_module/_06708_ ;
 wire \reg_module/_06709_ ;
 wire \reg_module/_06710_ ;
 wire \reg_module/_06711_ ;
 wire \reg_module/_06712_ ;
 wire \reg_module/_06713_ ;
 wire \reg_module/_06714_ ;
 wire \reg_module/_06715_ ;
 wire \reg_module/_06716_ ;
 wire \reg_module/_06717_ ;
 wire \reg_module/_06718_ ;
 wire \reg_module/_06719_ ;
 wire \reg_module/_06720_ ;
 wire \reg_module/_06721_ ;
 wire \reg_module/_06722_ ;
 wire \reg_module/_06723_ ;
 wire \reg_module/_06724_ ;
 wire \reg_module/_06725_ ;
 wire \reg_module/_06726_ ;
 wire \reg_module/_06727_ ;
 wire \reg_module/_06728_ ;
 wire \reg_module/_06729_ ;
 wire \reg_module/_06730_ ;
 wire \reg_module/_06731_ ;
 wire \reg_module/_06732_ ;
 wire \reg_module/_06733_ ;
 wire \reg_module/_06734_ ;
 wire \reg_module/_06735_ ;
 wire \reg_module/_06736_ ;
 wire \reg_module/_06737_ ;
 wire \reg_module/_06738_ ;
 wire \reg_module/_06739_ ;
 wire \reg_module/_06740_ ;
 wire \reg_module/_06741_ ;
 wire \reg_module/_06742_ ;
 wire \reg_module/_06743_ ;
 wire \reg_module/_06744_ ;
 wire \reg_module/_06745_ ;
 wire \reg_module/_06746_ ;
 wire \reg_module/_06747_ ;
 wire \reg_module/_06748_ ;
 wire \reg_module/_06749_ ;
 wire \reg_module/_06750_ ;
 wire \reg_module/_06751_ ;
 wire \reg_module/_06752_ ;
 wire \reg_module/_06753_ ;
 wire \reg_module/_06754_ ;
 wire \reg_module/_06755_ ;
 wire \reg_module/_06756_ ;
 wire \reg_module/_06757_ ;
 wire \reg_module/_06758_ ;
 wire \reg_module/_06759_ ;
 wire \reg_module/_06760_ ;
 wire \reg_module/_06761_ ;
 wire \reg_module/_06762_ ;
 wire \reg_module/_06763_ ;
 wire \reg_module/_06764_ ;
 wire \reg_module/_06765_ ;
 wire \reg_module/_06766_ ;
 wire \reg_module/_06767_ ;
 wire \reg_module/_06768_ ;
 wire \reg_module/_06769_ ;
 wire \reg_module/_06770_ ;
 wire \reg_module/_06771_ ;
 wire \reg_module/_06772_ ;
 wire \reg_module/_06773_ ;
 wire \reg_module/_06774_ ;
 wire \reg_module/_06775_ ;
 wire \reg_module/_06776_ ;
 wire \reg_module/_06777_ ;
 wire \reg_module/_06778_ ;
 wire \reg_module/_06779_ ;
 wire \reg_module/_06780_ ;
 wire \reg_module/_06781_ ;
 wire \reg_module/_06782_ ;
 wire \reg_module/_06783_ ;
 wire \reg_module/_06784_ ;
 wire \reg_module/_06785_ ;
 wire \reg_module/_06786_ ;
 wire \reg_module/_06787_ ;
 wire \reg_module/_06788_ ;
 wire \reg_module/_06789_ ;
 wire \reg_module/_06790_ ;
 wire \reg_module/_06791_ ;
 wire \reg_module/_06792_ ;
 wire \reg_module/_06793_ ;
 wire \reg_module/_06794_ ;
 wire \reg_module/_06795_ ;
 wire \reg_module/_06796_ ;
 wire \reg_module/_06797_ ;
 wire \reg_module/_06798_ ;
 wire \reg_module/_06799_ ;
 wire \reg_module/_06800_ ;
 wire \reg_module/_06801_ ;
 wire \reg_module/_06802_ ;
 wire \reg_module/_06803_ ;
 wire \reg_module/_06804_ ;
 wire \reg_module/_06805_ ;
 wire \reg_module/_06806_ ;
 wire \reg_module/_06807_ ;
 wire \reg_module/_06808_ ;
 wire \reg_module/_06809_ ;
 wire \reg_module/_06810_ ;
 wire \reg_module/_06811_ ;
 wire \reg_module/_06812_ ;
 wire \reg_module/_06813_ ;
 wire \reg_module/_06814_ ;
 wire \reg_module/_06815_ ;
 wire \reg_module/_06816_ ;
 wire \reg_module/_06817_ ;
 wire \reg_module/_06818_ ;
 wire \reg_module/_06819_ ;
 wire \reg_module/_06820_ ;
 wire \reg_module/_06821_ ;
 wire \reg_module/_06822_ ;
 wire \reg_module/_06823_ ;
 wire \reg_module/_06824_ ;
 wire \reg_module/_06825_ ;
 wire \reg_module/_06826_ ;
 wire \reg_module/_06827_ ;
 wire \reg_module/_06828_ ;
 wire \reg_module/_06829_ ;
 wire \reg_module/_06830_ ;
 wire \reg_module/_06831_ ;
 wire \reg_module/_06832_ ;
 wire \reg_module/_06833_ ;
 wire \reg_module/_06834_ ;
 wire \reg_module/_06835_ ;
 wire \reg_module/_06836_ ;
 wire \reg_module/_06837_ ;
 wire \reg_module/_06838_ ;
 wire \reg_module/_06839_ ;
 wire \reg_module/_06840_ ;
 wire \reg_module/_06841_ ;
 wire \reg_module/_06842_ ;
 wire \reg_module/_06843_ ;
 wire \reg_module/_06844_ ;
 wire \reg_module/_06845_ ;
 wire \reg_module/_06846_ ;
 wire \reg_module/_06847_ ;
 wire \reg_module/_06848_ ;
 wire \reg_module/_06849_ ;
 wire \reg_module/_06850_ ;
 wire \reg_module/_06851_ ;
 wire \reg_module/_06852_ ;
 wire \reg_module/_06853_ ;
 wire \reg_module/_06854_ ;
 wire \reg_module/_06855_ ;
 wire \reg_module/_06856_ ;
 wire \reg_module/_06857_ ;
 wire \reg_module/_06858_ ;
 wire \reg_module/_06859_ ;
 wire \reg_module/_06860_ ;
 wire \reg_module/_06861_ ;
 wire \reg_module/_06862_ ;
 wire \reg_module/_06863_ ;
 wire \reg_module/_06864_ ;
 wire \reg_module/_06865_ ;
 wire \reg_module/_06866_ ;
 wire \reg_module/_06867_ ;
 wire \reg_module/_06868_ ;
 wire \reg_module/_06869_ ;
 wire \reg_module/_06870_ ;
 wire \reg_module/_06871_ ;
 wire \reg_module/_06872_ ;
 wire \reg_module/_06873_ ;
 wire \reg_module/_06874_ ;
 wire \reg_module/_06875_ ;
 wire \reg_module/_06876_ ;
 wire \reg_module/_06877_ ;
 wire \reg_module/_06878_ ;
 wire \reg_module/_06879_ ;
 wire \reg_module/_06880_ ;
 wire \reg_module/_06881_ ;
 wire \reg_module/_06882_ ;
 wire \reg_module/_06883_ ;
 wire \reg_module/_06884_ ;
 wire \reg_module/_06885_ ;
 wire \reg_module/_06886_ ;
 wire \reg_module/_06887_ ;
 wire \reg_module/_06888_ ;
 wire \reg_module/_06889_ ;
 wire \reg_module/_06890_ ;
 wire \reg_module/_06891_ ;
 wire \reg_module/_06892_ ;
 wire \reg_module/_06893_ ;
 wire \reg_module/_06894_ ;
 wire \reg_module/_06895_ ;
 wire \reg_module/_06896_ ;
 wire \reg_module/_06897_ ;
 wire \reg_module/_06898_ ;
 wire \reg_module/_06899_ ;
 wire \reg_module/_06900_ ;
 wire \reg_module/_06901_ ;
 wire \reg_module/_06902_ ;
 wire \reg_module/_06903_ ;
 wire \reg_module/_06904_ ;
 wire \reg_module/_06905_ ;
 wire \reg_module/_06906_ ;
 wire \reg_module/_06907_ ;
 wire \reg_module/_06908_ ;
 wire \reg_module/_06909_ ;
 wire \reg_module/_06910_ ;
 wire \reg_module/_06911_ ;
 wire \reg_module/_06912_ ;
 wire \reg_module/_06913_ ;
 wire \reg_module/_06914_ ;
 wire \reg_module/_06915_ ;
 wire \reg_module/_06916_ ;
 wire \reg_module/_06917_ ;
 wire \reg_module/_06918_ ;
 wire \reg_module/_06919_ ;
 wire \reg_module/_06920_ ;
 wire \reg_module/_06921_ ;
 wire \reg_module/_06922_ ;
 wire \reg_module/_06923_ ;
 wire \reg_module/_06924_ ;
 wire \reg_module/_06925_ ;
 wire \reg_module/_06926_ ;
 wire \reg_module/_06927_ ;
 wire \reg_module/_06928_ ;
 wire \reg_module/_06929_ ;
 wire \reg_module/_06930_ ;
 wire \reg_module/_06931_ ;
 wire \reg_module/_06932_ ;
 wire \reg_module/_06933_ ;
 wire \reg_module/_06934_ ;
 wire \reg_module/_06935_ ;
 wire \reg_module/_06936_ ;
 wire \reg_module/_06937_ ;
 wire \reg_module/_06938_ ;
 wire \reg_module/_06939_ ;
 wire \reg_module/_06940_ ;
 wire \reg_module/_06941_ ;
 wire \reg_module/_06942_ ;
 wire \reg_module/_06943_ ;
 wire \reg_module/_06944_ ;
 wire \reg_module/_06945_ ;
 wire \reg_module/_06946_ ;
 wire \reg_module/_06947_ ;
 wire \reg_module/_06948_ ;
 wire \reg_module/_06949_ ;
 wire \reg_module/_06950_ ;
 wire \reg_module/_06951_ ;
 wire \reg_module/_06952_ ;
 wire \reg_module/_06953_ ;
 wire \reg_module/_06954_ ;
 wire \reg_module/_06955_ ;
 wire \reg_module/_06956_ ;
 wire \reg_module/_06957_ ;
 wire \reg_module/_06958_ ;
 wire \reg_module/_06959_ ;
 wire \reg_module/_06960_ ;
 wire \reg_module/_06961_ ;
 wire \reg_module/_06962_ ;
 wire \reg_module/_06963_ ;
 wire \reg_module/_06964_ ;
 wire \reg_module/_06965_ ;
 wire \reg_module/_06966_ ;
 wire \reg_module/_06967_ ;
 wire \reg_module/_06968_ ;
 wire \reg_module/_06969_ ;
 wire \reg_module/_06970_ ;
 wire \reg_module/_06971_ ;
 wire \reg_module/_06972_ ;
 wire \reg_module/_06973_ ;
 wire \reg_module/_06974_ ;
 wire \reg_module/_06975_ ;
 wire \reg_module/_06976_ ;
 wire \reg_module/_06977_ ;
 wire \reg_module/_06978_ ;
 wire \reg_module/_06979_ ;
 wire \reg_module/_06980_ ;
 wire \reg_module/_06981_ ;
 wire \reg_module/_06982_ ;
 wire \reg_module/_06983_ ;
 wire \reg_module/_06984_ ;
 wire \reg_module/_06985_ ;
 wire \reg_module/_06986_ ;
 wire \reg_module/_06987_ ;
 wire \reg_module/_06988_ ;
 wire \reg_module/_06989_ ;
 wire \reg_module/_06990_ ;
 wire \reg_module/_06991_ ;
 wire \reg_module/_06992_ ;
 wire \reg_module/_06993_ ;
 wire \reg_module/_06994_ ;
 wire \reg_module/_06995_ ;
 wire \reg_module/_06996_ ;
 wire \reg_module/_06997_ ;
 wire \reg_module/_06998_ ;
 wire \reg_module/_06999_ ;
 wire \reg_module/_07000_ ;
 wire \reg_module/_07001_ ;
 wire \reg_module/_07002_ ;
 wire \reg_module/_07003_ ;
 wire \reg_module/_07004_ ;
 wire \reg_module/_07005_ ;
 wire \reg_module/_07006_ ;
 wire \reg_module/_07007_ ;
 wire \reg_module/_07008_ ;
 wire \reg_module/_07009_ ;
 wire \reg_module/_07010_ ;
 wire \reg_module/_07011_ ;
 wire \reg_module/_07012_ ;
 wire \reg_module/_07013_ ;
 wire \reg_module/_07014_ ;
 wire \reg_module/_07015_ ;
 wire \reg_module/_07016_ ;
 wire \reg_module/_07017_ ;
 wire \reg_module/_07018_ ;
 wire \reg_module/_07019_ ;
 wire \reg_module/_07020_ ;
 wire \reg_module/_07021_ ;
 wire \reg_module/_07022_ ;
 wire \reg_module/_07023_ ;
 wire \reg_module/_07024_ ;
 wire \reg_module/_07025_ ;
 wire \reg_module/_07026_ ;
 wire \reg_module/_07027_ ;
 wire \reg_module/_07028_ ;
 wire \reg_module/_07029_ ;
 wire \reg_module/_07030_ ;
 wire \reg_module/_07031_ ;
 wire \reg_module/_07032_ ;
 wire \reg_module/_07033_ ;
 wire \reg_module/_07034_ ;
 wire \reg_module/_07035_ ;
 wire \reg_module/_07036_ ;
 wire \reg_module/_07037_ ;
 wire \reg_module/_07038_ ;
 wire \reg_module/_07039_ ;
 wire \reg_module/_07040_ ;
 wire \reg_module/_07041_ ;
 wire \reg_module/_07042_ ;
 wire \reg_module/_07043_ ;
 wire \reg_module/_07044_ ;
 wire \reg_module/_07045_ ;
 wire \reg_module/_07046_ ;
 wire \reg_module/_07047_ ;
 wire \reg_module/_07048_ ;
 wire \reg_module/_07049_ ;
 wire \reg_module/_07050_ ;
 wire \reg_module/_07051_ ;
 wire \reg_module/_07052_ ;
 wire \reg_module/_07053_ ;
 wire \reg_module/_07054_ ;
 wire \reg_module/_07055_ ;
 wire \reg_module/_07056_ ;
 wire \reg_module/_07057_ ;
 wire \reg_module/_07058_ ;
 wire \reg_module/_07059_ ;
 wire \reg_module/_07060_ ;
 wire \reg_module/_07061_ ;
 wire \reg_module/_07062_ ;
 wire \reg_module/_07063_ ;
 wire \reg_module/_07064_ ;
 wire \reg_module/_07065_ ;
 wire \reg_module/_07066_ ;
 wire \reg_module/_07067_ ;
 wire \reg_module/_07068_ ;
 wire \reg_module/_07069_ ;
 wire \reg_module/_07070_ ;
 wire \reg_module/_07071_ ;
 wire \reg_module/_07072_ ;
 wire \reg_module/_07073_ ;
 wire \reg_module/_07074_ ;
 wire \reg_module/_07075_ ;
 wire \reg_module/_07076_ ;
 wire \reg_module/_07077_ ;
 wire \reg_module/_07078_ ;
 wire \reg_module/_07079_ ;
 wire \reg_module/_07080_ ;
 wire \reg_module/_07081_ ;
 wire \reg_module/_07082_ ;
 wire \reg_module/_07083_ ;
 wire \reg_module/_07084_ ;
 wire \reg_module/_07085_ ;
 wire \reg_module/_07086_ ;
 wire \reg_module/_07087_ ;
 wire \reg_module/_07088_ ;
 wire \reg_module/_07089_ ;
 wire \reg_module/_07090_ ;
 wire \reg_module/_07091_ ;
 wire \reg_module/_07092_ ;
 wire \reg_module/_07093_ ;
 wire \reg_module/_07094_ ;
 wire \reg_module/_07095_ ;
 wire \reg_module/_07096_ ;
 wire \reg_module/_07097_ ;
 wire \reg_module/_07098_ ;
 wire \reg_module/_07099_ ;
 wire \reg_module/_07100_ ;
 wire \reg_module/_07101_ ;
 wire \reg_module/_07102_ ;
 wire \reg_module/_07103_ ;
 wire \reg_module/_07104_ ;
 wire \reg_module/_07105_ ;
 wire \reg_module/_07106_ ;
 wire \reg_module/_07107_ ;
 wire \reg_module/_07108_ ;
 wire \reg_module/_07109_ ;
 wire \reg_module/_07110_ ;
 wire \reg_module/_07111_ ;
 wire \reg_module/_07112_ ;
 wire \reg_module/_07113_ ;
 wire \reg_module/_07114_ ;
 wire \reg_module/_07115_ ;
 wire \reg_module/_07116_ ;
 wire \reg_module/_07117_ ;
 wire \reg_module/_07118_ ;
 wire \reg_module/_07119_ ;
 wire \reg_module/_07120_ ;
 wire \reg_module/_07121_ ;
 wire \reg_module/_07122_ ;
 wire \reg_module/_07123_ ;
 wire \reg_module/_07124_ ;
 wire \reg_module/_07125_ ;
 wire \reg_module/_07126_ ;
 wire \reg_module/_07127_ ;
 wire \reg_module/_07128_ ;
 wire \reg_module/_07129_ ;
 wire \reg_module/_07130_ ;
 wire \reg_module/_07131_ ;
 wire \reg_module/_07132_ ;
 wire \reg_module/_07133_ ;
 wire \reg_module/_07134_ ;
 wire \reg_module/_07135_ ;
 wire \reg_module/_07136_ ;
 wire \reg_module/_07137_ ;
 wire \reg_module/_07138_ ;
 wire \reg_module/_07139_ ;
 wire \reg_module/_07140_ ;
 wire \reg_module/_07141_ ;
 wire \reg_module/_07142_ ;
 wire \reg_module/_07143_ ;
 wire \reg_module/_07144_ ;
 wire \reg_module/_07145_ ;
 wire \reg_module/_07146_ ;
 wire \reg_module/_07147_ ;
 wire \reg_module/_07148_ ;
 wire \reg_module/_07149_ ;
 wire \reg_module/_07150_ ;
 wire \reg_module/_07151_ ;
 wire \reg_module/_07152_ ;
 wire \reg_module/_07153_ ;
 wire \reg_module/_07154_ ;
 wire \reg_module/_07155_ ;
 wire \reg_module/_07156_ ;
 wire \reg_module/_07157_ ;
 wire \reg_module/_07158_ ;
 wire \reg_module/_07159_ ;
 wire \reg_module/_07160_ ;
 wire \reg_module/_07161_ ;
 wire \reg_module/_07162_ ;
 wire \reg_module/_07163_ ;
 wire \reg_module/_07164_ ;
 wire \reg_module/_07165_ ;
 wire \reg_module/_07166_ ;
 wire \reg_module/_07167_ ;
 wire \reg_module/_07168_ ;
 wire \reg_module/_07169_ ;
 wire \reg_module/_07170_ ;
 wire \reg_module/_07171_ ;
 wire \reg_module/_07172_ ;
 wire \reg_module/_07173_ ;
 wire \reg_module/_07174_ ;
 wire \reg_module/_07175_ ;
 wire \reg_module/_07176_ ;
 wire \reg_module/_07177_ ;
 wire \reg_module/_07178_ ;
 wire \reg_module/_07179_ ;
 wire \reg_module/_07180_ ;
 wire \reg_module/_07181_ ;
 wire \reg_module/_07182_ ;
 wire \reg_module/_07183_ ;
 wire \reg_module/_07184_ ;
 wire \reg_module/_07185_ ;
 wire \reg_module/_07186_ ;
 wire \reg_module/_07187_ ;
 wire \reg_module/_07188_ ;
 wire \reg_module/_07189_ ;
 wire \reg_module/_07190_ ;
 wire \reg_module/_07191_ ;
 wire \reg_module/_07192_ ;
 wire \reg_module/_07193_ ;
 wire \reg_module/_07194_ ;
 wire \reg_module/_07195_ ;
 wire \reg_module/_07196_ ;
 wire \reg_module/_07197_ ;
 wire \reg_module/_07198_ ;
 wire \reg_module/_07199_ ;
 wire \reg_module/_07200_ ;
 wire \reg_module/_07201_ ;
 wire \reg_module/_07202_ ;
 wire \reg_module/_07203_ ;
 wire \reg_module/_07204_ ;
 wire \reg_module/_07205_ ;
 wire \reg_module/_07206_ ;
 wire \reg_module/_07207_ ;
 wire \reg_module/_07208_ ;
 wire \reg_module/_07209_ ;
 wire \reg_module/_07210_ ;
 wire \reg_module/_07211_ ;
 wire \reg_module/_07212_ ;
 wire \reg_module/_07213_ ;
 wire \reg_module/_07214_ ;
 wire \reg_module/_07215_ ;
 wire \reg_module/_07216_ ;
 wire \reg_module/_07217_ ;
 wire \reg_module/_07218_ ;
 wire \reg_module/_07219_ ;
 wire \reg_module/_07220_ ;
 wire \reg_module/_07221_ ;
 wire \reg_module/_07222_ ;
 wire \reg_module/_07223_ ;
 wire \reg_module/_07224_ ;
 wire \reg_module/_07225_ ;
 wire \reg_module/_07226_ ;
 wire \reg_module/_07227_ ;
 wire \reg_module/_07228_ ;
 wire \reg_module/_07229_ ;
 wire \reg_module/_07230_ ;
 wire \reg_module/_07231_ ;
 wire \reg_module/_07232_ ;
 wire \reg_module/_07233_ ;
 wire \reg_module/_07234_ ;
 wire \reg_module/_07235_ ;
 wire \reg_module/_07236_ ;
 wire \reg_module/_07237_ ;
 wire \reg_module/_07238_ ;
 wire \reg_module/_07239_ ;
 wire \reg_module/_07240_ ;
 wire \reg_module/_07241_ ;
 wire \reg_module/_07242_ ;
 wire \reg_module/_07243_ ;
 wire \reg_module/_07244_ ;
 wire \reg_module/_07245_ ;
 wire \reg_module/_07246_ ;
 wire \reg_module/_07247_ ;
 wire \reg_module/_07248_ ;
 wire \reg_module/_07249_ ;
 wire \reg_module/_07250_ ;
 wire \reg_module/_07251_ ;
 wire \reg_module/_07252_ ;
 wire \reg_module/_07253_ ;
 wire \reg_module/_07254_ ;
 wire \reg_module/_07255_ ;
 wire \reg_module/_07256_ ;
 wire \reg_module/_07257_ ;
 wire \reg_module/_07258_ ;
 wire \reg_module/_07259_ ;
 wire \reg_module/_07260_ ;
 wire \reg_module/_07261_ ;
 wire \reg_module/_07262_ ;
 wire \reg_module/_07263_ ;
 wire \reg_module/_07264_ ;
 wire \reg_module/_07265_ ;
 wire \reg_module/_07266_ ;
 wire \reg_module/_07267_ ;
 wire \reg_module/_07268_ ;
 wire \reg_module/_07269_ ;
 wire \reg_module/_07270_ ;
 wire \reg_module/_07271_ ;
 wire \reg_module/_07272_ ;
 wire \reg_module/_07273_ ;
 wire \reg_module/_07274_ ;
 wire \reg_module/_07275_ ;
 wire \reg_module/_07276_ ;
 wire \reg_module/_07277_ ;
 wire \reg_module/_07278_ ;
 wire \reg_module/_07279_ ;
 wire \reg_module/_07280_ ;
 wire \reg_module/_07281_ ;
 wire \reg_module/_07282_ ;
 wire \reg_module/_07283_ ;
 wire \reg_module/_07284_ ;
 wire \reg_module/_07285_ ;
 wire \reg_module/_07286_ ;
 wire \reg_module/_07287_ ;
 wire \reg_module/_07288_ ;
 wire \reg_module/_07289_ ;
 wire \reg_module/_07290_ ;
 wire \reg_module/_07291_ ;
 wire \reg_module/_07292_ ;
 wire \reg_module/_07293_ ;
 wire \reg_module/_07294_ ;
 wire \reg_module/_07295_ ;
 wire \reg_module/_07296_ ;
 wire \reg_module/_07297_ ;
 wire \reg_module/_07298_ ;
 wire \reg_module/_07299_ ;
 wire \reg_module/_07300_ ;
 wire \reg_module/_07301_ ;
 wire \reg_module/_07302_ ;
 wire \reg_module/_07303_ ;
 wire \reg_module/_07304_ ;
 wire \reg_module/_07305_ ;
 wire \reg_module/_07306_ ;
 wire \reg_module/_07307_ ;
 wire \reg_module/_07308_ ;
 wire \reg_module/_07309_ ;
 wire \reg_module/_07310_ ;
 wire \reg_module/_07311_ ;
 wire \reg_module/_07312_ ;
 wire \reg_module/_07313_ ;
 wire \reg_module/_07314_ ;
 wire \reg_module/_07315_ ;
 wire \reg_module/_07316_ ;
 wire \reg_module/_07317_ ;
 wire \reg_module/_07318_ ;
 wire \reg_module/_07319_ ;
 wire \reg_module/_07320_ ;
 wire \reg_module/_07321_ ;
 wire \reg_module/_07322_ ;
 wire \reg_module/_07323_ ;
 wire \reg_module/_07324_ ;
 wire \reg_module/_07325_ ;
 wire \reg_module/_07326_ ;
 wire \reg_module/_07327_ ;
 wire \reg_module/_07328_ ;
 wire \reg_module/_07329_ ;
 wire \reg_module/_07330_ ;
 wire \reg_module/_07331_ ;
 wire \reg_module/_07332_ ;
 wire \reg_module/_07333_ ;
 wire \reg_module/_07334_ ;
 wire \reg_module/_07335_ ;
 wire \reg_module/_07336_ ;
 wire \reg_module/_07337_ ;
 wire \reg_module/_07338_ ;
 wire \reg_module/_07339_ ;
 wire \reg_module/_07340_ ;
 wire \reg_module/_07341_ ;
 wire \reg_module/_07342_ ;
 wire \reg_module/_07343_ ;
 wire \reg_module/_07344_ ;
 wire \reg_module/_07345_ ;
 wire \reg_module/_07346_ ;
 wire \reg_module/_07347_ ;
 wire \reg_module/_07348_ ;
 wire \reg_module/_07349_ ;
 wire \reg_module/_07350_ ;
 wire \reg_module/_07351_ ;
 wire \reg_module/_07352_ ;
 wire \reg_module/_07353_ ;
 wire \reg_module/_07354_ ;
 wire \reg_module/_07355_ ;
 wire \reg_module/_07356_ ;
 wire \reg_module/_07357_ ;
 wire \reg_module/_07358_ ;
 wire \reg_module/_07359_ ;
 wire \reg_module/_07360_ ;
 wire \reg_module/_07361_ ;
 wire \reg_module/_07362_ ;
 wire \reg_module/_07363_ ;
 wire \reg_module/_07364_ ;
 wire \reg_module/_07365_ ;
 wire \reg_module/_07366_ ;
 wire \reg_module/_07367_ ;
 wire \reg_module/_07368_ ;
 wire \reg_module/_07369_ ;
 wire \reg_module/_07370_ ;
 wire \reg_module/_07371_ ;
 wire \reg_module/_07372_ ;
 wire \reg_module/_07373_ ;
 wire \reg_module/_07374_ ;
 wire \reg_module/_07375_ ;
 wire \reg_module/_07376_ ;
 wire \reg_module/_07377_ ;
 wire \reg_module/_07378_ ;
 wire \reg_module/_07379_ ;
 wire \reg_module/_07380_ ;
 wire \reg_module/_07381_ ;
 wire \reg_module/_07382_ ;
 wire \reg_module/_07383_ ;
 wire \reg_module/_07384_ ;
 wire \reg_module/_07385_ ;
 wire \reg_module/_07386_ ;
 wire \reg_module/_07387_ ;
 wire \reg_module/_07388_ ;
 wire \reg_module/_07389_ ;
 wire \reg_module/_07390_ ;
 wire \reg_module/_07391_ ;
 wire \reg_module/_07392_ ;
 wire \reg_module/_07393_ ;
 wire \reg_module/_07394_ ;
 wire \reg_module/_07395_ ;
 wire \reg_module/_07396_ ;
 wire \reg_module/_07397_ ;
 wire \reg_module/_07398_ ;
 wire \reg_module/_07399_ ;
 wire \reg_module/_07400_ ;
 wire \reg_module/_07401_ ;
 wire \reg_module/_07402_ ;
 wire \reg_module/_07403_ ;
 wire \reg_module/_07404_ ;
 wire \reg_module/_07405_ ;
 wire \reg_module/_07406_ ;
 wire \reg_module/_07407_ ;
 wire \reg_module/_07408_ ;
 wire \reg_module/_07409_ ;
 wire \reg_module/_07410_ ;
 wire \reg_module/_07411_ ;
 wire \reg_module/_07412_ ;
 wire \reg_module/_07413_ ;
 wire \reg_module/_07414_ ;
 wire \reg_module/_07415_ ;
 wire \reg_module/_07416_ ;
 wire \reg_module/_07417_ ;
 wire \reg_module/_07418_ ;
 wire \reg_module/_07419_ ;
 wire \reg_module/_07420_ ;
 wire \reg_module/_07421_ ;
 wire \reg_module/_07422_ ;
 wire \reg_module/_07423_ ;
 wire \reg_module/_07424_ ;
 wire \reg_module/_07425_ ;
 wire \reg_module/_07426_ ;
 wire \reg_module/_07427_ ;
 wire \reg_module/_07428_ ;
 wire \reg_module/_07429_ ;
 wire \reg_module/_07430_ ;
 wire \reg_module/_07431_ ;
 wire \reg_module/_07432_ ;
 wire \reg_module/_07433_ ;
 wire \reg_module/_07434_ ;
 wire \reg_module/_07435_ ;
 wire \reg_module/_07436_ ;
 wire \reg_module/_07437_ ;
 wire \reg_module/_07438_ ;
 wire \reg_module/_07439_ ;
 wire \reg_module/_07440_ ;
 wire \reg_module/_07441_ ;
 wire \reg_module/_07442_ ;
 wire \reg_module/_07443_ ;
 wire \reg_module/_07444_ ;
 wire \reg_module/_07445_ ;
 wire \reg_module/_07446_ ;
 wire \reg_module/_07447_ ;
 wire \reg_module/_07448_ ;
 wire \reg_module/_07449_ ;
 wire \reg_module/_07450_ ;
 wire \reg_module/_07451_ ;
 wire \reg_module/_07452_ ;
 wire \reg_module/_07453_ ;
 wire \reg_module/_07454_ ;
 wire \reg_module/_07455_ ;
 wire \reg_module/_07456_ ;
 wire \reg_module/_07457_ ;
 wire \reg_module/_07458_ ;
 wire \reg_module/_07459_ ;
 wire \reg_module/_07460_ ;
 wire \reg_module/_07461_ ;
 wire \reg_module/_07462_ ;
 wire \reg_module/_07463_ ;
 wire \reg_module/_07464_ ;
 wire \reg_module/_07465_ ;
 wire \reg_module/_07466_ ;
 wire \reg_module/_07467_ ;
 wire \reg_module/_07468_ ;
 wire \reg_module/_07469_ ;
 wire \reg_module/_07470_ ;
 wire \reg_module/_07471_ ;
 wire \reg_module/_07472_ ;
 wire \reg_module/_07473_ ;
 wire \reg_module/_07474_ ;
 wire \reg_module/_07475_ ;
 wire \reg_module/_07476_ ;
 wire \reg_module/_07477_ ;
 wire \reg_module/_07478_ ;
 wire \reg_module/_07479_ ;
 wire \reg_module/_07480_ ;
 wire \reg_module/_07481_ ;
 wire \reg_module/_07482_ ;
 wire \reg_module/_07483_ ;
 wire \reg_module/_07484_ ;
 wire \reg_module/_07485_ ;
 wire \reg_module/_07486_ ;
 wire \reg_module/_07487_ ;
 wire \reg_module/_07488_ ;
 wire \reg_module/_07489_ ;
 wire \reg_module/_07490_ ;
 wire \reg_module/_07491_ ;
 wire \reg_module/_07492_ ;
 wire \reg_module/_07493_ ;
 wire \reg_module/_07494_ ;
 wire \reg_module/_07495_ ;
 wire \reg_module/_07496_ ;
 wire \reg_module/_07497_ ;
 wire \reg_module/_07498_ ;
 wire \reg_module/_07499_ ;
 wire \reg_module/_07500_ ;
 wire \reg_module/_07501_ ;
 wire \reg_module/_07502_ ;
 wire \reg_module/_07503_ ;
 wire \reg_module/_07504_ ;
 wire \reg_module/_07505_ ;
 wire \reg_module/_07506_ ;
 wire \reg_module/_07507_ ;
 wire \reg_module/_07508_ ;
 wire \reg_module/_07509_ ;
 wire \reg_module/_07510_ ;
 wire \reg_module/_07511_ ;
 wire \reg_module/_07512_ ;
 wire \reg_module/_07513_ ;
 wire \reg_module/_07514_ ;
 wire \reg_module/_07515_ ;
 wire \reg_module/_07516_ ;
 wire \reg_module/_07517_ ;
 wire \reg_module/_07518_ ;
 wire \reg_module/_07519_ ;
 wire \reg_module/_07520_ ;
 wire \reg_module/_07521_ ;
 wire \reg_module/_07522_ ;
 wire \reg_module/_07523_ ;
 wire \reg_module/_07524_ ;
 wire \reg_module/_07525_ ;
 wire \reg_module/_07526_ ;
 wire \reg_module/_07527_ ;
 wire \reg_module/_07528_ ;
 wire \reg_module/_07529_ ;
 wire \reg_module/_07530_ ;
 wire \reg_module/_07531_ ;
 wire \reg_module/_07532_ ;
 wire \reg_module/_07533_ ;
 wire \reg_module/_07534_ ;
 wire \reg_module/_07535_ ;
 wire \reg_module/_07536_ ;
 wire \reg_module/_07537_ ;
 wire \reg_module/_07538_ ;
 wire \reg_module/_07539_ ;
 wire \reg_module/_07540_ ;
 wire \reg_module/_07541_ ;
 wire \reg_module/_07542_ ;
 wire \reg_module/_07543_ ;
 wire \reg_module/_07544_ ;
 wire \reg_module/_07545_ ;
 wire \reg_module/_07546_ ;
 wire \reg_module/_07547_ ;
 wire \reg_module/_07548_ ;
 wire \reg_module/_07549_ ;
 wire \reg_module/_07550_ ;
 wire \reg_module/_07551_ ;
 wire \reg_module/_07552_ ;
 wire \reg_module/_07553_ ;
 wire \reg_module/_07554_ ;
 wire \reg_module/_07555_ ;
 wire \reg_module/_07556_ ;
 wire \reg_module/_07557_ ;
 wire \reg_module/_07558_ ;
 wire \reg_module/_07559_ ;
 wire \reg_module/_07560_ ;
 wire \reg_module/_07561_ ;
 wire \reg_module/_07562_ ;
 wire \reg_module/_07563_ ;
 wire \reg_module/_07564_ ;
 wire \reg_module/_07565_ ;
 wire \reg_module/_07566_ ;
 wire \reg_module/_07567_ ;
 wire \reg_module/_07568_ ;
 wire \reg_module/_07569_ ;
 wire \reg_module/_07570_ ;
 wire \reg_module/_07571_ ;
 wire \reg_module/_07572_ ;
 wire \reg_module/_07573_ ;
 wire \reg_module/_07574_ ;
 wire \reg_module/_07575_ ;
 wire \reg_module/_07576_ ;
 wire \reg_module/_07577_ ;
 wire \reg_module/_07578_ ;
 wire \reg_module/_07579_ ;
 wire \reg_module/_07580_ ;
 wire \reg_module/_07581_ ;
 wire \reg_module/_07582_ ;
 wire \reg_module/_07583_ ;
 wire \reg_module/_07584_ ;
 wire \reg_module/_07585_ ;
 wire \reg_module/_07586_ ;
 wire \reg_module/_07587_ ;
 wire \reg_module/_07588_ ;
 wire \reg_module/_07589_ ;
 wire \reg_module/_07590_ ;
 wire \reg_module/_07591_ ;
 wire \reg_module/_07592_ ;
 wire \reg_module/_07593_ ;
 wire \reg_module/_07594_ ;
 wire \reg_module/_07595_ ;
 wire \reg_module/_07596_ ;
 wire \reg_module/_07597_ ;
 wire \reg_module/_07598_ ;
 wire \reg_module/_07599_ ;
 wire \reg_module/_07600_ ;
 wire \reg_module/_07601_ ;
 wire \reg_module/_07602_ ;
 wire \reg_module/_07603_ ;
 wire \reg_module/_07604_ ;
 wire \reg_module/_07605_ ;
 wire \reg_module/_07606_ ;
 wire \reg_module/_07607_ ;
 wire \reg_module/_07608_ ;
 wire \reg_module/_07609_ ;
 wire \reg_module/_07610_ ;
 wire \reg_module/_07611_ ;
 wire \reg_module/_07612_ ;
 wire \reg_module/_07613_ ;
 wire \reg_module/_07614_ ;
 wire \reg_module/_07615_ ;
 wire \reg_module/_07616_ ;
 wire \reg_module/_07617_ ;
 wire \reg_module/_07618_ ;
 wire \reg_module/_07619_ ;
 wire \reg_module/_07620_ ;
 wire \reg_module/_07621_ ;
 wire \reg_module/_07622_ ;
 wire \reg_module/_07623_ ;
 wire \reg_module/_07624_ ;
 wire \reg_module/_07625_ ;
 wire \reg_module/_07626_ ;
 wire \reg_module/_07627_ ;
 wire \reg_module/_07628_ ;
 wire \reg_module/_07629_ ;
 wire \reg_module/_07630_ ;
 wire \reg_module/_07631_ ;
 wire \reg_module/_07632_ ;
 wire \reg_module/_07633_ ;
 wire \reg_module/_07634_ ;
 wire \reg_module/_07635_ ;
 wire \reg_module/_07636_ ;
 wire \reg_module/_07637_ ;
 wire \reg_module/_07638_ ;
 wire \reg_module/_07639_ ;
 wire \reg_module/_07640_ ;
 wire \reg_module/_07641_ ;
 wire \reg_module/_07642_ ;
 wire \reg_module/_07643_ ;
 wire \reg_module/_07644_ ;
 wire \reg_module/_07645_ ;
 wire \reg_module/_07646_ ;
 wire \reg_module/_07647_ ;
 wire \reg_module/_07648_ ;
 wire \reg_module/_07649_ ;
 wire \reg_module/_07650_ ;
 wire \reg_module/_07651_ ;
 wire \reg_module/_07652_ ;
 wire \reg_module/_07653_ ;
 wire \reg_module/_07654_ ;
 wire \reg_module/_07655_ ;
 wire \reg_module/_07656_ ;
 wire \reg_module/_07657_ ;
 wire \reg_module/_07658_ ;
 wire \reg_module/_07659_ ;
 wire \reg_module/_07660_ ;
 wire \reg_module/_07661_ ;
 wire \reg_module/_07662_ ;
 wire \reg_module/_07663_ ;
 wire \reg_module/_07664_ ;
 wire \reg_module/_07665_ ;
 wire \reg_module/_07666_ ;
 wire \reg_module/_07667_ ;
 wire \reg_module/_07668_ ;
 wire \reg_module/_07669_ ;
 wire \reg_module/_07670_ ;
 wire \reg_module/_07671_ ;
 wire \reg_module/_07672_ ;
 wire \reg_module/_07673_ ;
 wire \reg_module/_07674_ ;
 wire \reg_module/_07675_ ;
 wire \reg_module/_07676_ ;
 wire \reg_module/_07677_ ;
 wire \reg_module/_07678_ ;
 wire \reg_module/_07679_ ;
 wire \reg_module/_07680_ ;
 wire \reg_module/_07681_ ;
 wire \reg_module/_07682_ ;
 wire \reg_module/_07683_ ;
 wire \reg_module/_07684_ ;
 wire \reg_module/_07685_ ;
 wire \reg_module/_07686_ ;
 wire \reg_module/_07687_ ;
 wire \reg_module/_07688_ ;
 wire \reg_module/_07689_ ;
 wire \reg_module/_07690_ ;
 wire \reg_module/_07691_ ;
 wire \reg_module/_07692_ ;
 wire \reg_module/_07693_ ;
 wire \reg_module/_07694_ ;
 wire \reg_module/_07695_ ;
 wire \reg_module/_07696_ ;
 wire \reg_module/_07697_ ;
 wire \reg_module/_07698_ ;
 wire \reg_module/_07699_ ;
 wire \reg_module/_07700_ ;
 wire \reg_module/_07701_ ;
 wire \reg_module/_07702_ ;
 wire \reg_module/_07703_ ;
 wire \reg_module/_07704_ ;
 wire \reg_module/_07705_ ;
 wire \reg_module/_07706_ ;
 wire \reg_module/_07707_ ;
 wire \reg_module/_07708_ ;
 wire \reg_module/_07709_ ;
 wire \reg_module/_07710_ ;
 wire \reg_module/_07711_ ;
 wire \reg_module/_07712_ ;
 wire \reg_module/_07713_ ;
 wire \reg_module/_07714_ ;
 wire \reg_module/_07715_ ;
 wire \reg_module/_07716_ ;
 wire \reg_module/_07717_ ;
 wire \reg_module/_07718_ ;
 wire \reg_module/_07719_ ;
 wire \reg_module/_07720_ ;
 wire \reg_module/_07721_ ;
 wire \reg_module/_07722_ ;
 wire \reg_module/_07723_ ;
 wire \reg_module/_07724_ ;
 wire \reg_module/_07725_ ;
 wire \reg_module/_07726_ ;
 wire \reg_module/_07727_ ;
 wire \reg_module/_07728_ ;
 wire \reg_module/_07729_ ;
 wire \reg_module/_07730_ ;
 wire \reg_module/_07731_ ;
 wire \reg_module/_07732_ ;
 wire \reg_module/_07733_ ;
 wire \reg_module/_07734_ ;
 wire \reg_module/_07735_ ;
 wire \reg_module/_07736_ ;
 wire \reg_module/_07737_ ;
 wire \reg_module/_07738_ ;
 wire \reg_module/_07739_ ;
 wire \reg_module/_07740_ ;
 wire \reg_module/_07741_ ;
 wire \reg_module/_07742_ ;
 wire \reg_module/_07743_ ;
 wire \reg_module/_07744_ ;
 wire \reg_module/_07745_ ;
 wire \reg_module/_07746_ ;
 wire \reg_module/_07747_ ;
 wire \reg_module/_07748_ ;
 wire \reg_module/_07749_ ;
 wire \reg_module/_07750_ ;
 wire \reg_module/_07751_ ;
 wire \reg_module/_07752_ ;
 wire \reg_module/_07753_ ;
 wire \reg_module/_07754_ ;
 wire \reg_module/_07755_ ;
 wire \reg_module/_07756_ ;
 wire \reg_module/_07757_ ;
 wire \reg_module/_07758_ ;
 wire \reg_module/_07759_ ;
 wire \reg_module/_07760_ ;
 wire \reg_module/_07761_ ;
 wire \reg_module/_07762_ ;
 wire \reg_module/_07763_ ;
 wire \reg_module/_07764_ ;
 wire \reg_module/_07765_ ;
 wire \reg_module/_07766_ ;
 wire \reg_module/_07767_ ;
 wire \reg_module/_07768_ ;
 wire \reg_module/_07769_ ;
 wire \reg_module/_07770_ ;
 wire \reg_module/_07771_ ;
 wire \reg_module/_07772_ ;
 wire \reg_module/_07773_ ;
 wire \reg_module/_07774_ ;
 wire \reg_module/_07775_ ;
 wire \reg_module/_07776_ ;
 wire \reg_module/_07777_ ;
 wire \reg_module/_07778_ ;
 wire \reg_module/_07779_ ;
 wire \reg_module/_07780_ ;
 wire \reg_module/_07781_ ;
 wire \reg_module/_07782_ ;
 wire \reg_module/_07783_ ;
 wire \reg_module/_07784_ ;
 wire \reg_module/_07785_ ;
 wire \reg_module/_07786_ ;
 wire \reg_module/_07787_ ;
 wire \reg_module/_07788_ ;
 wire \reg_module/_07789_ ;
 wire \reg_module/_07790_ ;
 wire \reg_module/_07791_ ;
 wire \reg_module/_07792_ ;
 wire \reg_module/_07793_ ;
 wire \reg_module/_07794_ ;
 wire \reg_module/_07795_ ;
 wire \reg_module/_07796_ ;
 wire \reg_module/_07797_ ;
 wire \reg_module/_07798_ ;
 wire \reg_module/_07799_ ;
 wire \reg_module/_07800_ ;
 wire \reg_module/_07801_ ;
 wire \reg_module/_07802_ ;
 wire \reg_module/_07803_ ;
 wire \reg_module/_07804_ ;
 wire \reg_module/_07805_ ;
 wire \reg_module/_07806_ ;
 wire \reg_module/_07807_ ;
 wire \reg_module/_07808_ ;
 wire \reg_module/_07809_ ;
 wire \reg_module/_07810_ ;
 wire \reg_module/_07811_ ;
 wire \reg_module/_07812_ ;
 wire \reg_module/_07813_ ;
 wire \reg_module/_07814_ ;
 wire \reg_module/_07815_ ;
 wire \reg_module/_07816_ ;
 wire \reg_module/_07817_ ;
 wire \reg_module/_07818_ ;
 wire \reg_module/_07819_ ;
 wire \reg_module/_07820_ ;
 wire \reg_module/_07821_ ;
 wire \reg_module/_07822_ ;
 wire \reg_module/_07823_ ;
 wire \reg_module/_07824_ ;
 wire \reg_module/_07825_ ;
 wire \reg_module/_07826_ ;
 wire \reg_module/_07827_ ;
 wire \reg_module/_07828_ ;
 wire \reg_module/_07829_ ;
 wire \reg_module/_07830_ ;
 wire \reg_module/_07831_ ;
 wire \reg_module/_07832_ ;
 wire \reg_module/_07833_ ;
 wire \reg_module/_07834_ ;
 wire \reg_module/_07835_ ;
 wire \reg_module/_07836_ ;
 wire \reg_module/_07837_ ;
 wire \reg_module/_07838_ ;
 wire \reg_module/_07839_ ;
 wire \reg_module/_07840_ ;
 wire \reg_module/_07841_ ;
 wire \reg_module/_07842_ ;
 wire \reg_module/_07843_ ;
 wire \reg_module/_07844_ ;
 wire \reg_module/_07845_ ;
 wire \reg_module/_07846_ ;
 wire \reg_module/_07847_ ;
 wire \reg_module/_07848_ ;
 wire \reg_module/_07849_ ;
 wire \reg_module/_07850_ ;
 wire \reg_module/_07851_ ;
 wire \reg_module/_07852_ ;
 wire \reg_module/_07853_ ;
 wire \reg_module/_07854_ ;
 wire \reg_module/_07855_ ;
 wire \reg_module/_07856_ ;
 wire \reg_module/_07857_ ;
 wire \reg_module/_07858_ ;
 wire \reg_module/_07859_ ;
 wire \reg_module/_07860_ ;
 wire \reg_module/_07861_ ;
 wire \reg_module/_07862_ ;
 wire \reg_module/_07863_ ;
 wire \reg_module/_07864_ ;
 wire \reg_module/_07865_ ;
 wire \reg_module/_07866_ ;
 wire \reg_module/_07867_ ;
 wire \reg_module/_07868_ ;
 wire \reg_module/_07869_ ;
 wire \reg_module/_07870_ ;
 wire \reg_module/_07871_ ;
 wire \reg_module/_07872_ ;
 wire \reg_module/_07873_ ;
 wire \reg_module/_07874_ ;
 wire \reg_module/_07875_ ;
 wire \reg_module/_07876_ ;
 wire \reg_module/_07877_ ;
 wire \reg_module/_07878_ ;
 wire \reg_module/_07879_ ;
 wire \reg_module/_07880_ ;
 wire \reg_module/_07881_ ;
 wire \reg_module/_07882_ ;
 wire \reg_module/_07883_ ;
 wire \reg_module/_07884_ ;
 wire \reg_module/_07885_ ;
 wire \reg_module/_07886_ ;
 wire \reg_module/_07887_ ;
 wire \reg_module/_07888_ ;
 wire \reg_module/_07889_ ;
 wire \reg_module/_07890_ ;
 wire \reg_module/_07891_ ;
 wire \reg_module/_07892_ ;
 wire \reg_module/_07893_ ;
 wire \reg_module/_07894_ ;
 wire \reg_module/_07895_ ;
 wire \reg_module/_07896_ ;
 wire \reg_module/_07897_ ;
 wire \reg_module/_07898_ ;
 wire \reg_module/_07899_ ;
 wire \reg_module/_07900_ ;
 wire \reg_module/_07901_ ;
 wire \reg_module/_07902_ ;
 wire \reg_module/_07903_ ;
 wire \reg_module/_07904_ ;
 wire \reg_module/_07905_ ;
 wire \reg_module/_07906_ ;
 wire \reg_module/_07907_ ;
 wire \reg_module/_07908_ ;
 wire \reg_module/_07909_ ;
 wire \reg_module/_07910_ ;
 wire \reg_module/_07911_ ;
 wire \reg_module/_07912_ ;
 wire \reg_module/_07913_ ;
 wire \reg_module/_07914_ ;
 wire \reg_module/_07915_ ;
 wire \reg_module/_07916_ ;
 wire \reg_module/_07917_ ;
 wire \reg_module/_07918_ ;
 wire \reg_module/_07919_ ;
 wire \reg_module/_07920_ ;
 wire \reg_module/_07921_ ;
 wire \reg_module/_07922_ ;
 wire \reg_module/_07923_ ;
 wire \reg_module/_07924_ ;
 wire \reg_module/_07925_ ;
 wire \reg_module/_07926_ ;
 wire \reg_module/_07927_ ;
 wire \reg_module/_07928_ ;
 wire \reg_module/_07929_ ;
 wire \reg_module/_07930_ ;
 wire \reg_module/_07931_ ;
 wire \reg_module/_07932_ ;
 wire \reg_module/_07933_ ;
 wire \reg_module/_07934_ ;
 wire \reg_module/_07935_ ;
 wire \reg_module/_07936_ ;
 wire \reg_module/_07937_ ;
 wire \reg_module/_07938_ ;
 wire \reg_module/_07939_ ;
 wire \reg_module/_07940_ ;
 wire \reg_module/_07941_ ;
 wire \reg_module/_07942_ ;
 wire \reg_module/_07943_ ;
 wire \reg_module/_07944_ ;
 wire \reg_module/_07945_ ;
 wire \reg_module/_07946_ ;
 wire \reg_module/_07947_ ;
 wire \reg_module/_07948_ ;
 wire \reg_module/_07949_ ;
 wire \reg_module/_07950_ ;
 wire \reg_module/_07951_ ;
 wire \reg_module/_07952_ ;
 wire \reg_module/_07953_ ;
 wire \reg_module/_07954_ ;
 wire \reg_module/_07955_ ;
 wire \reg_module/_07956_ ;
 wire \reg_module/_07957_ ;
 wire \reg_module/_07958_ ;
 wire \reg_module/_07959_ ;
 wire \reg_module/_07960_ ;
 wire \reg_module/_07961_ ;
 wire \reg_module/_07962_ ;
 wire \reg_module/_07963_ ;
 wire \reg_module/_07964_ ;
 wire \reg_module/_07965_ ;
 wire \reg_module/_07966_ ;
 wire \reg_module/_07967_ ;
 wire \reg_module/_07968_ ;
 wire \reg_module/_07969_ ;
 wire \reg_module/_07970_ ;
 wire \reg_module/_07971_ ;
 wire \reg_module/_07972_ ;
 wire \reg_module/_07973_ ;
 wire \reg_module/_07974_ ;
 wire \reg_module/_07975_ ;
 wire \reg_module/_07976_ ;
 wire \reg_module/_07977_ ;
 wire \reg_module/_07978_ ;
 wire \reg_module/_07979_ ;
 wire \reg_module/_07980_ ;
 wire \reg_module/_07981_ ;
 wire \reg_module/_07982_ ;
 wire \reg_module/_07983_ ;
 wire \reg_module/_07984_ ;
 wire \reg_module/_07985_ ;
 wire \reg_module/_07986_ ;
 wire \reg_module/_07987_ ;
 wire \reg_module/_07988_ ;
 wire \reg_module/_07989_ ;
 wire \reg_module/_07990_ ;
 wire \reg_module/_07991_ ;
 wire \reg_module/_07992_ ;
 wire \reg_module/_07993_ ;
 wire \reg_module/_07994_ ;
 wire \reg_module/_07995_ ;
 wire \reg_module/_07996_ ;
 wire \reg_module/_07997_ ;
 wire \reg_module/_07998_ ;
 wire \reg_module/_07999_ ;
 wire \reg_module/_08000_ ;
 wire \reg_module/_08001_ ;
 wire \reg_module/_08002_ ;
 wire \reg_module/_08003_ ;
 wire \reg_module/_08004_ ;
 wire \reg_module/_08005_ ;
 wire \reg_module/_08006_ ;
 wire \reg_module/_08007_ ;
 wire \reg_module/_08008_ ;
 wire \reg_module/_08009_ ;
 wire \reg_module/_08010_ ;
 wire \reg_module/_08011_ ;
 wire \reg_module/_08012_ ;
 wire \reg_module/_08013_ ;
 wire \reg_module/_08014_ ;
 wire \reg_module/_08015_ ;
 wire \reg_module/_08016_ ;
 wire \reg_module/_08017_ ;
 wire \reg_module/_08018_ ;
 wire \reg_module/_08019_ ;
 wire \reg_module/_08020_ ;
 wire \reg_module/_08021_ ;
 wire \reg_module/_08022_ ;
 wire \reg_module/_08023_ ;
 wire \reg_module/_08024_ ;
 wire \reg_module/_08025_ ;
 wire \reg_module/_08026_ ;
 wire \reg_module/_08027_ ;
 wire \reg_module/_08028_ ;
 wire \reg_module/_08029_ ;
 wire \reg_module/_08030_ ;
 wire \reg_module/_08031_ ;
 wire \reg_module/_08032_ ;
 wire \reg_module/_08033_ ;
 wire \reg_module/_08034_ ;
 wire \reg_module/_08035_ ;
 wire \reg_module/_08036_ ;
 wire \reg_module/_08037_ ;
 wire \reg_module/_08038_ ;
 wire \reg_module/_08039_ ;
 wire \reg_module/_08040_ ;
 wire \reg_module/_08041_ ;
 wire \reg_module/_08042_ ;
 wire \reg_module/_08043_ ;
 wire \reg_module/_08044_ ;
 wire \reg_module/_08045_ ;
 wire \reg_module/_08046_ ;
 wire \reg_module/_08047_ ;
 wire \reg_module/_08048_ ;
 wire \reg_module/_08049_ ;
 wire \reg_module/_08050_ ;
 wire \reg_module/_08051_ ;
 wire \reg_module/_08052_ ;
 wire \reg_module/_08053_ ;
 wire \reg_module/_08054_ ;
 wire \reg_module/_08055_ ;
 wire \reg_module/_08056_ ;
 wire \reg_module/_08057_ ;
 wire \reg_module/_08058_ ;
 wire \reg_module/_08059_ ;
 wire \reg_module/_08060_ ;
 wire \reg_module/_08061_ ;
 wire \reg_module/_08062_ ;
 wire \reg_module/_08063_ ;
 wire \reg_module/_08064_ ;
 wire \reg_module/_08065_ ;
 wire \reg_module/_08066_ ;
 wire \reg_module/_08067_ ;
 wire \reg_module/_08068_ ;
 wire \reg_module/_08069_ ;
 wire \reg_module/_08070_ ;
 wire \reg_module/_08071_ ;
 wire \reg_module/_08072_ ;
 wire \reg_module/_08073_ ;
 wire \reg_module/_08074_ ;
 wire \reg_module/_08075_ ;
 wire \reg_module/_08076_ ;
 wire \reg_module/_08077_ ;
 wire \reg_module/_08078_ ;
 wire \reg_module/_08079_ ;
 wire \reg_module/_08080_ ;
 wire \reg_module/_08081_ ;
 wire \reg_module/_08082_ ;
 wire \reg_module/_08083_ ;
 wire \reg_module/_08084_ ;
 wire \reg_module/_08085_ ;
 wire \reg_module/_08086_ ;
 wire \reg_module/_08087_ ;
 wire \reg_module/_08088_ ;
 wire \reg_module/_08089_ ;
 wire \reg_module/_08090_ ;
 wire \reg_module/_08091_ ;
 wire \reg_module/_08092_ ;
 wire \reg_module/_08093_ ;
 wire \reg_module/_08094_ ;
 wire \reg_module/_08095_ ;
 wire \reg_module/_08096_ ;
 wire \reg_module/_08097_ ;
 wire \reg_module/_08098_ ;
 wire \reg_module/_08099_ ;
 wire \reg_module/_08100_ ;
 wire \reg_module/_08101_ ;
 wire \reg_module/_08102_ ;
 wire \reg_module/_08103_ ;
 wire \reg_module/_08104_ ;
 wire \reg_module/_08105_ ;
 wire \reg_module/_08106_ ;
 wire \reg_module/_08107_ ;
 wire \reg_module/_08108_ ;
 wire \reg_module/_08109_ ;
 wire \reg_module/_08110_ ;
 wire \reg_module/_08111_ ;
 wire \reg_module/_08112_ ;
 wire \reg_module/_08113_ ;
 wire \reg_module/_08114_ ;
 wire \reg_module/_08115_ ;
 wire \reg_module/_08116_ ;
 wire \reg_module/_08117_ ;
 wire \reg_module/_08118_ ;
 wire \reg_module/_08119_ ;
 wire \reg_module/_08120_ ;
 wire \reg_module/_08121_ ;
 wire \reg_module/_08122_ ;
 wire \reg_module/_08123_ ;
 wire \reg_module/_08124_ ;
 wire \reg_module/_08125_ ;
 wire \reg_module/_08126_ ;
 wire \reg_module/_08127_ ;
 wire \reg_module/_08128_ ;
 wire \reg_module/_08129_ ;
 wire \reg_module/_08130_ ;
 wire \reg_module/_08131_ ;
 wire \reg_module/_08132_ ;
 wire \reg_module/_08133_ ;
 wire \reg_module/_08134_ ;
 wire \reg_module/_08135_ ;
 wire \reg_module/_08136_ ;
 wire \reg_module/_08137_ ;
 wire \reg_module/_08138_ ;
 wire \reg_module/_08139_ ;
 wire \reg_module/_08140_ ;
 wire \reg_module/_08141_ ;
 wire \reg_module/_08142_ ;
 wire \reg_module/_08143_ ;
 wire \reg_module/_08144_ ;
 wire \reg_module/_08145_ ;
 wire \reg_module/_08146_ ;
 wire \reg_module/_08147_ ;
 wire \reg_module/_08148_ ;
 wire \reg_module/_08149_ ;
 wire \reg_module/_08150_ ;
 wire \reg_module/_08151_ ;
 wire \reg_module/_08152_ ;
 wire \reg_module/_08153_ ;
 wire \reg_module/_08154_ ;
 wire \reg_module/_08155_ ;
 wire \reg_module/_08156_ ;
 wire \reg_module/_08157_ ;
 wire \reg_module/_08158_ ;
 wire \reg_module/_08159_ ;
 wire \reg_module/_08160_ ;
 wire \reg_module/_08161_ ;
 wire \reg_module/_08162_ ;
 wire \reg_module/_08163_ ;
 wire \reg_module/_08164_ ;
 wire \reg_module/_08165_ ;
 wire \reg_module/_08166_ ;
 wire \reg_module/_08167_ ;
 wire \reg_module/_08168_ ;
 wire \reg_module/_08169_ ;
 wire \reg_module/_08170_ ;
 wire \reg_module/_08171_ ;
 wire \reg_module/_08172_ ;
 wire \reg_module/_08173_ ;
 wire \reg_module/_08174_ ;
 wire \reg_module/_08175_ ;
 wire \reg_module/_08176_ ;
 wire \reg_module/_08177_ ;
 wire \reg_module/_08178_ ;
 wire \reg_module/_08179_ ;
 wire \reg_module/_08180_ ;
 wire \reg_module/_08181_ ;
 wire \reg_module/_08182_ ;
 wire \reg_module/_08183_ ;
 wire \reg_module/_08184_ ;
 wire \reg_module/_08185_ ;
 wire \reg_module/_08186_ ;
 wire \reg_module/_08187_ ;
 wire \reg_module/_08188_ ;
 wire \reg_module/_08189_ ;
 wire \reg_module/_08190_ ;
 wire \reg_module/_08191_ ;
 wire \reg_module/_08192_ ;
 wire \reg_module/_08193_ ;
 wire \reg_module/_08194_ ;
 wire \reg_module/_08195_ ;
 wire \reg_module/_08196_ ;
 wire \reg_module/_08197_ ;
 wire \reg_module/_08198_ ;
 wire \reg_module/_08199_ ;
 wire \reg_module/_08200_ ;
 wire \reg_module/_08201_ ;
 wire \reg_module/_08202_ ;
 wire \reg_module/_08203_ ;
 wire \reg_module/_08204_ ;
 wire \reg_module/_08205_ ;
 wire \reg_module/_08206_ ;
 wire \reg_module/_08207_ ;
 wire \reg_module/_08208_ ;
 wire \reg_module/_08209_ ;
 wire \reg_module/_08210_ ;
 wire \reg_module/_08211_ ;
 wire \reg_module/_08212_ ;
 wire \reg_module/_08213_ ;
 wire \reg_module/_08214_ ;
 wire \reg_module/_08215_ ;
 wire \reg_module/_08216_ ;
 wire \reg_module/_08217_ ;
 wire \reg_module/_08218_ ;
 wire \reg_module/_08219_ ;
 wire \reg_module/_08220_ ;
 wire \reg_module/_08221_ ;
 wire \reg_module/_08222_ ;
 wire \reg_module/_08223_ ;
 wire \reg_module/_08224_ ;
 wire \reg_module/_08225_ ;
 wire \reg_module/_08226_ ;
 wire \reg_module/_08227_ ;
 wire \reg_module/_08228_ ;
 wire \reg_module/_08229_ ;
 wire \reg_module/_08230_ ;
 wire \reg_module/_08231_ ;
 wire \reg_module/_08232_ ;
 wire \reg_module/_08233_ ;
 wire \reg_module/_08234_ ;
 wire \reg_module/_08235_ ;
 wire \reg_module/_08236_ ;
 wire \reg_module/_08237_ ;
 wire \reg_module/_08238_ ;
 wire \reg_module/_08239_ ;
 wire \reg_module/_08240_ ;
 wire \reg_module/_08241_ ;
 wire \reg_module/_08242_ ;
 wire \reg_module/_08243_ ;
 wire \reg_module/_08244_ ;
 wire \reg_module/_08245_ ;
 wire \reg_module/_08246_ ;
 wire \reg_module/_08247_ ;
 wire \reg_module/_08248_ ;
 wire \reg_module/_08249_ ;
 wire \reg_module/_08250_ ;
 wire \reg_module/_08251_ ;
 wire \reg_module/_08252_ ;
 wire \reg_module/_08253_ ;
 wire \reg_module/_08254_ ;
 wire \reg_module/_08255_ ;
 wire \reg_module/_08256_ ;
 wire \reg_module/_08257_ ;
 wire \reg_module/_08258_ ;
 wire \reg_module/_08259_ ;
 wire \reg_module/_08260_ ;
 wire \reg_module/_08261_ ;
 wire \reg_module/_08262_ ;
 wire \reg_module/_08263_ ;
 wire \reg_module/_08264_ ;
 wire \reg_module/_08265_ ;
 wire \reg_module/_08266_ ;
 wire \reg_module/_08267_ ;
 wire \reg_module/_08268_ ;
 wire \reg_module/_08269_ ;
 wire \reg_module/_08270_ ;
 wire \reg_module/_08271_ ;
 wire \reg_module/_08272_ ;
 wire \reg_module/_08273_ ;
 wire \reg_module/_08274_ ;
 wire \reg_module/_08275_ ;
 wire \reg_module/_08276_ ;
 wire \reg_module/_08277_ ;
 wire \reg_module/_08278_ ;
 wire \reg_module/_08279_ ;
 wire \reg_module/_08280_ ;
 wire \reg_module/_08281_ ;
 wire \reg_module/_08282_ ;
 wire \reg_module/_08283_ ;
 wire \reg_module/_08284_ ;
 wire \reg_module/_08285_ ;
 wire \reg_module/_08286_ ;
 wire \reg_module/_08287_ ;
 wire \reg_module/_08288_ ;
 wire \reg_module/_08289_ ;
 wire \reg_module/_08290_ ;
 wire \reg_module/_08291_ ;
 wire \reg_module/_08292_ ;
 wire \reg_module/_08293_ ;
 wire \reg_module/_08294_ ;
 wire \reg_module/_08295_ ;
 wire \reg_module/_08296_ ;
 wire \reg_module/_08297_ ;
 wire \reg_module/_08298_ ;
 wire \reg_module/_08299_ ;
 wire \reg_module/_08300_ ;
 wire \reg_module/_08301_ ;
 wire \reg_module/_08302_ ;
 wire \reg_module/_08303_ ;
 wire \reg_module/_08304_ ;
 wire \reg_module/_08305_ ;
 wire \reg_module/_08306_ ;
 wire \reg_module/_08307_ ;
 wire \reg_module/_08308_ ;
 wire \reg_module/_08309_ ;
 wire \reg_module/_08310_ ;
 wire \reg_module/_08311_ ;
 wire \reg_module/_08312_ ;
 wire \reg_module/_08313_ ;
 wire \reg_module/_08314_ ;
 wire \reg_module/_08315_ ;
 wire \reg_module/_08316_ ;
 wire \reg_module/_08317_ ;
 wire \reg_module/_08318_ ;
 wire \reg_module/_08319_ ;
 wire \reg_module/_08320_ ;
 wire \reg_module/_08321_ ;
 wire \reg_module/_08322_ ;
 wire \reg_module/_08323_ ;
 wire \reg_module/_08324_ ;
 wire \reg_module/_08325_ ;
 wire \reg_module/_08326_ ;
 wire \reg_module/_08327_ ;
 wire \reg_module/_08328_ ;
 wire \reg_module/_08329_ ;
 wire \reg_module/_08330_ ;
 wire \reg_module/_08331_ ;
 wire \reg_module/_08332_ ;
 wire \reg_module/_08333_ ;
 wire \reg_module/_08334_ ;
 wire \reg_module/_08335_ ;
 wire \reg_module/_08336_ ;
 wire \reg_module/_08337_ ;
 wire \reg_module/_08338_ ;
 wire \reg_module/_08339_ ;
 wire \reg_module/_08340_ ;
 wire \reg_module/_08341_ ;
 wire \reg_module/_08342_ ;
 wire \reg_module/_08343_ ;
 wire \reg_module/_08344_ ;
 wire \reg_module/_08345_ ;
 wire \reg_module/_08346_ ;
 wire \reg_module/_08347_ ;
 wire \reg_module/_08348_ ;
 wire \reg_module/_08349_ ;
 wire \reg_module/_08350_ ;
 wire \reg_module/_08351_ ;
 wire \reg_module/_08352_ ;
 wire \reg_module/_08353_ ;
 wire \reg_module/_08354_ ;
 wire \reg_module/_08355_ ;
 wire \reg_module/_08356_ ;
 wire \reg_module/_08357_ ;
 wire \reg_module/_08358_ ;
 wire \reg_module/_08359_ ;
 wire \reg_module/_08360_ ;
 wire \reg_module/_08361_ ;
 wire \reg_module/_08362_ ;
 wire \reg_module/_08363_ ;
 wire \reg_module/_08364_ ;
 wire \reg_module/_08365_ ;
 wire \reg_module/_08366_ ;
 wire \reg_module/_08367_ ;
 wire \reg_module/_08368_ ;
 wire \reg_module/_08369_ ;
 wire \reg_module/_08370_ ;
 wire \reg_module/_08371_ ;
 wire \reg_module/_08372_ ;
 wire \reg_module/_08373_ ;
 wire \reg_module/_08374_ ;
 wire \reg_module/_08375_ ;
 wire \reg_module/_08376_ ;
 wire \reg_module/_08377_ ;
 wire \reg_module/_08378_ ;
 wire \reg_module/_08379_ ;
 wire \reg_module/_08380_ ;
 wire \reg_module/_08381_ ;
 wire \reg_module/_08382_ ;
 wire \reg_module/_08383_ ;
 wire \reg_module/_08384_ ;
 wire \reg_module/_08385_ ;
 wire \reg_module/_08386_ ;
 wire \reg_module/_08387_ ;
 wire \reg_module/_08388_ ;
 wire \reg_module/_08389_ ;
 wire \reg_module/_08390_ ;
 wire \reg_module/_08391_ ;
 wire \reg_module/_08392_ ;
 wire \reg_module/_08393_ ;
 wire \reg_module/_08394_ ;
 wire \reg_module/_08395_ ;
 wire \reg_module/_08396_ ;
 wire \reg_module/_08397_ ;
 wire \reg_module/_08398_ ;
 wire \reg_module/_08399_ ;
 wire \reg_module/_08400_ ;
 wire \reg_module/_08401_ ;
 wire \reg_module/_08402_ ;
 wire \reg_module/_08403_ ;
 wire \reg_module/_08404_ ;
 wire \reg_module/_08405_ ;
 wire \reg_module/_08406_ ;
 wire \reg_module/_08407_ ;
 wire \reg_module/_08408_ ;
 wire \reg_module/_08409_ ;
 wire \reg_module/_08410_ ;
 wire \reg_module/_08411_ ;
 wire \reg_module/_08412_ ;
 wire \reg_module/_08413_ ;
 wire \reg_module/_08414_ ;
 wire \reg_module/_08415_ ;
 wire \reg_module/_08416_ ;
 wire \reg_module/_08417_ ;
 wire \reg_module/_08418_ ;
 wire \reg_module/_08419_ ;
 wire \reg_module/_08420_ ;
 wire \reg_module/_08421_ ;
 wire \reg_module/_08422_ ;
 wire \reg_module/_08423_ ;
 wire \reg_module/_08424_ ;
 wire \reg_module/_08425_ ;
 wire \reg_module/_08426_ ;
 wire \reg_module/_08427_ ;
 wire \reg_module/_08428_ ;
 wire \reg_module/_08429_ ;
 wire \reg_module/_08430_ ;
 wire \reg_module/_08431_ ;
 wire \reg_module/_08432_ ;
 wire \reg_module/_08433_ ;
 wire \reg_module/_08434_ ;
 wire \reg_module/_08435_ ;
 wire \reg_module/_08436_ ;
 wire \reg_module/_08437_ ;
 wire \reg_module/_08438_ ;
 wire \reg_module/_08439_ ;
 wire \reg_module/_08440_ ;
 wire \reg_module/_08441_ ;
 wire \reg_module/_08442_ ;
 wire \reg_module/_08443_ ;
 wire \reg_module/_08444_ ;
 wire \reg_module/_08445_ ;
 wire \reg_module/_08446_ ;
 wire \reg_module/_08447_ ;
 wire \reg_module/_08448_ ;
 wire \reg_module/_08449_ ;
 wire \reg_module/_08450_ ;
 wire \reg_module/_08451_ ;
 wire \reg_module/_08452_ ;
 wire \reg_module/_08453_ ;
 wire \reg_module/_08454_ ;
 wire \reg_module/_08455_ ;
 wire \reg_module/_08456_ ;
 wire \reg_module/_08457_ ;
 wire \reg_module/_08458_ ;
 wire \reg_module/_08459_ ;
 wire \reg_module/_08460_ ;
 wire \reg_module/_08461_ ;
 wire \reg_module/_08462_ ;
 wire \reg_module/_08463_ ;
 wire \reg_module/_08464_ ;
 wire \reg_module/_08465_ ;
 wire \reg_module/_08466_ ;
 wire \reg_module/_08467_ ;
 wire \reg_module/_08468_ ;
 wire \reg_module/_08469_ ;
 wire \reg_module/_08470_ ;
 wire \reg_module/_08471_ ;
 wire \reg_module/_08472_ ;
 wire \reg_module/_08473_ ;
 wire \reg_module/_08474_ ;
 wire \reg_module/_08475_ ;
 wire \reg_module/_08476_ ;
 wire \reg_module/_08477_ ;
 wire \reg_module/_08478_ ;
 wire \reg_module/_08479_ ;
 wire \reg_module/_08480_ ;
 wire \reg_module/_08481_ ;
 wire \reg_module/_08482_ ;
 wire \reg_module/_08483_ ;
 wire \reg_module/_08484_ ;
 wire \reg_module/_08485_ ;
 wire \reg_module/_08486_ ;
 wire \reg_module/_08487_ ;
 wire \reg_module/_08488_ ;
 wire \reg_module/_08489_ ;
 wire \reg_module/_08490_ ;
 wire \reg_module/_08491_ ;
 wire \reg_module/_08492_ ;
 wire \reg_module/_08493_ ;
 wire \reg_module/_08494_ ;
 wire \reg_module/_08495_ ;
 wire \reg_module/_08496_ ;
 wire \reg_module/_08497_ ;
 wire \reg_module/_08498_ ;
 wire \reg_module/_08499_ ;
 wire \reg_module/_08500_ ;
 wire \reg_module/_08501_ ;
 wire \reg_module/_08502_ ;
 wire \reg_module/_08503_ ;
 wire \reg_module/_08504_ ;
 wire \reg_module/_08505_ ;
 wire \reg_module/_08506_ ;
 wire \reg_module/_08507_ ;
 wire \reg_module/_08508_ ;
 wire \reg_module/_08509_ ;
 wire \reg_module/_08510_ ;
 wire \reg_module/_08511_ ;
 wire \reg_module/_08512_ ;
 wire \reg_module/_08513_ ;
 wire \reg_module/_08514_ ;
 wire \reg_module/_08515_ ;
 wire \reg_module/_08516_ ;
 wire \reg_module/_08517_ ;
 wire \reg_module/_08518_ ;
 wire \reg_module/_08519_ ;
 wire \reg_module/_08520_ ;
 wire \reg_module/_08521_ ;
 wire \reg_module/_08522_ ;
 wire \reg_module/_08523_ ;
 wire \reg_module/_08524_ ;
 wire \reg_module/_08525_ ;
 wire \reg_module/_08526_ ;
 wire \reg_module/_08527_ ;
 wire \reg_module/_08528_ ;
 wire \reg_module/_08529_ ;
 wire \reg_module/_08530_ ;
 wire \reg_module/_08531_ ;
 wire \reg_module/_08532_ ;
 wire \reg_module/_08533_ ;
 wire \reg_module/_08534_ ;
 wire \reg_module/_08535_ ;
 wire \reg_module/_08536_ ;
 wire \reg_module/_08537_ ;
 wire \reg_module/_08538_ ;
 wire \reg_module/_08539_ ;
 wire \reg_module/_08540_ ;
 wire \reg_module/_08541_ ;
 wire \reg_module/_08542_ ;
 wire \reg_module/_08543_ ;
 wire \reg_module/_08544_ ;
 wire \reg_module/_08545_ ;
 wire \reg_module/_08546_ ;
 wire \reg_module/_08547_ ;
 wire \reg_module/_08548_ ;
 wire \reg_module/_08549_ ;
 wire \reg_module/_08550_ ;
 wire \reg_module/_08551_ ;
 wire \reg_module/_08552_ ;
 wire \reg_module/_08553_ ;
 wire \reg_module/_08554_ ;
 wire \reg_module/_08555_ ;
 wire \reg_module/_08556_ ;
 wire \reg_module/_08557_ ;
 wire \reg_module/_08558_ ;
 wire \reg_module/_08559_ ;
 wire \reg_module/_08560_ ;
 wire \reg_module/_08561_ ;
 wire \reg_module/_08562_ ;
 wire \reg_module/_08563_ ;
 wire \reg_module/_08564_ ;
 wire \reg_module/_08565_ ;
 wire \reg_module/_08566_ ;
 wire \reg_module/_08567_ ;
 wire \reg_module/_08568_ ;
 wire \reg_module/_08569_ ;
 wire \reg_module/_08570_ ;
 wire \reg_module/_08571_ ;
 wire \reg_module/_08572_ ;
 wire \reg_module/_08573_ ;
 wire \reg_module/_08574_ ;
 wire \reg_module/_08575_ ;
 wire \reg_module/_08576_ ;
 wire \reg_module/_08577_ ;
 wire \reg_module/_08578_ ;
 wire \reg_module/_08579_ ;
 wire \reg_module/_08580_ ;
 wire \reg_module/_08581_ ;
 wire \reg_module/_08582_ ;
 wire \reg_module/_08583_ ;
 wire \reg_module/_08584_ ;
 wire \reg_module/_08585_ ;
 wire \reg_module/_08586_ ;
 wire \reg_module/_08587_ ;
 wire \reg_module/_08588_ ;
 wire \reg_module/_08589_ ;
 wire \reg_module/_08590_ ;
 wire \reg_module/_08591_ ;
 wire \reg_module/_08592_ ;
 wire \reg_module/_08593_ ;
 wire \reg_module/_08594_ ;
 wire \reg_module/_08595_ ;
 wire \reg_module/_08596_ ;
 wire \reg_module/_08597_ ;
 wire \reg_module/_08598_ ;
 wire \reg_module/_08599_ ;
 wire \reg_module/_08600_ ;
 wire \reg_module/_08601_ ;
 wire \reg_module/_08602_ ;
 wire \reg_module/_08603_ ;
 wire \reg_module/_08604_ ;
 wire \reg_module/_08605_ ;
 wire \reg_module/_08606_ ;
 wire \reg_module/_08607_ ;
 wire \reg_module/_08608_ ;
 wire \reg_module/_08609_ ;
 wire \reg_module/_08610_ ;
 wire \reg_module/_08611_ ;
 wire \reg_module/_08612_ ;
 wire \reg_module/_08613_ ;
 wire \reg_module/_08614_ ;
 wire \reg_module/_08615_ ;
 wire \reg_module/_08616_ ;
 wire \reg_module/_08617_ ;
 wire \reg_module/_08618_ ;
 wire \reg_module/_08619_ ;
 wire \reg_module/_08620_ ;
 wire \reg_module/_08621_ ;
 wire \reg_module/_08622_ ;
 wire \reg_module/_08623_ ;
 wire \reg_module/_08624_ ;
 wire \reg_module/_08625_ ;
 wire \reg_module/_08626_ ;
 wire \reg_module/_08627_ ;
 wire \reg_module/_08628_ ;
 wire \reg_module/_08629_ ;
 wire \reg_module/_08630_ ;
 wire \reg_module/_08631_ ;
 wire \reg_module/_08632_ ;
 wire \reg_module/_08633_ ;
 wire \reg_module/_08634_ ;
 wire \reg_module/_08635_ ;
 wire \reg_module/_08636_ ;
 wire \reg_module/_08637_ ;
 wire \reg_module/_08638_ ;
 wire \reg_module/_08639_ ;
 wire \reg_module/_08640_ ;
 wire \reg_module/_08641_ ;
 wire \reg_module/_08642_ ;
 wire \reg_module/_08643_ ;
 wire \reg_module/_08644_ ;
 wire \reg_module/_08645_ ;
 wire \reg_module/_08646_ ;
 wire \reg_module/_08647_ ;
 wire \reg_module/_08648_ ;
 wire \reg_module/_08649_ ;
 wire \reg_module/_08650_ ;
 wire \reg_module/_08651_ ;
 wire \reg_module/_08652_ ;
 wire \reg_module/_08653_ ;
 wire \reg_module/_08654_ ;
 wire \reg_module/_08655_ ;
 wire \reg_module/_08656_ ;
 wire \reg_module/_08657_ ;
 wire \reg_module/_08658_ ;
 wire \reg_module/_08659_ ;
 wire \reg_module/_08660_ ;
 wire \reg_module/_08661_ ;
 wire \reg_module/_08662_ ;
 wire \reg_module/_08663_ ;
 wire \reg_module/_08664_ ;
 wire \reg_module/_08665_ ;
 wire \reg_module/_08666_ ;
 wire \reg_module/_08667_ ;
 wire \reg_module/_08668_ ;
 wire \reg_module/_08669_ ;
 wire \reg_module/_08670_ ;
 wire \reg_module/_08671_ ;
 wire \reg_module/_08672_ ;
 wire \reg_module/_08673_ ;
 wire \reg_module/_08674_ ;
 wire \reg_module/_08675_ ;
 wire \reg_module/_08676_ ;
 wire \reg_module/_08677_ ;
 wire \reg_module/_08678_ ;
 wire \reg_module/_08679_ ;
 wire \reg_module/_08680_ ;
 wire \reg_module/_08681_ ;
 wire \reg_module/_08682_ ;
 wire \reg_module/_08683_ ;
 wire \reg_module/_08684_ ;
 wire \reg_module/_08685_ ;
 wire \reg_module/_08686_ ;
 wire \reg_module/_08687_ ;
 wire \reg_module/_08688_ ;
 wire \reg_module/_08689_ ;
 wire \reg_module/_08690_ ;
 wire \reg_module/_08691_ ;
 wire \reg_module/_08692_ ;
 wire \reg_module/_08693_ ;
 wire \reg_module/_08694_ ;
 wire \reg_module/_08695_ ;
 wire \reg_module/_08696_ ;
 wire \reg_module/_08697_ ;
 wire \reg_module/_08698_ ;
 wire \reg_module/_08699_ ;
 wire \reg_module/_08700_ ;
 wire \reg_module/_08701_ ;
 wire \reg_module/_08702_ ;
 wire \reg_module/_08703_ ;
 wire \reg_module/_08704_ ;
 wire \reg_module/_08705_ ;
 wire \reg_module/_08706_ ;
 wire \reg_module/_08707_ ;
 wire \reg_module/_08708_ ;
 wire \reg_module/_08709_ ;
 wire \reg_module/_08710_ ;
 wire \reg_module/_08711_ ;
 wire \reg_module/_08712_ ;
 wire \reg_module/_08713_ ;
 wire \reg_module/_08714_ ;
 wire \reg_module/_08715_ ;
 wire \reg_module/_08716_ ;
 wire \reg_module/_08717_ ;
 wire \reg_module/_08718_ ;
 wire \reg_module/_08719_ ;
 wire \reg_module/_08720_ ;
 wire \reg_module/_08721_ ;
 wire \reg_module/_08722_ ;
 wire \reg_module/_08723_ ;
 wire \reg_module/_08724_ ;
 wire \reg_module/_08725_ ;
 wire \reg_module/_08726_ ;
 wire \reg_module/_08727_ ;
 wire \reg_module/_08728_ ;
 wire \reg_module/_08729_ ;
 wire \reg_module/_08730_ ;
 wire \reg_module/_08731_ ;
 wire \reg_module/_08732_ ;
 wire \reg_module/_08733_ ;
 wire \reg_module/_08734_ ;
 wire \reg_module/_08735_ ;
 wire \reg_module/_08736_ ;
 wire \reg_module/_08737_ ;
 wire \reg_module/_08738_ ;
 wire \reg_module/_08739_ ;
 wire \reg_module/_08740_ ;
 wire \reg_module/_08741_ ;
 wire \reg_module/_08742_ ;
 wire \reg_module/_08743_ ;
 wire \reg_module/_08744_ ;
 wire \reg_module/_08745_ ;
 wire \reg_module/_08746_ ;
 wire \reg_module/_08747_ ;
 wire \reg_module/_08748_ ;
 wire \reg_module/_08749_ ;
 wire \reg_module/_08750_ ;
 wire \reg_module/_08751_ ;
 wire \reg_module/_08752_ ;
 wire \reg_module/_08753_ ;
 wire \reg_module/_08754_ ;
 wire \reg_module/_08755_ ;
 wire \reg_module/_08756_ ;
 wire \reg_module/_08757_ ;
 wire \reg_module/_08758_ ;
 wire \reg_module/_08759_ ;
 wire \reg_module/_08760_ ;
 wire \reg_module/_08761_ ;
 wire \reg_module/_08762_ ;
 wire \reg_module/_08763_ ;
 wire \reg_module/_08764_ ;
 wire \reg_module/_08765_ ;
 wire \reg_module/_08766_ ;
 wire \reg_module/_08767_ ;
 wire \reg_module/_08768_ ;
 wire \reg_module/_08769_ ;
 wire \reg_module/_08770_ ;
 wire \reg_module/_08771_ ;
 wire \reg_module/_08772_ ;
 wire \reg_module/_08773_ ;
 wire \reg_module/_08774_ ;
 wire \reg_module/_08775_ ;
 wire \reg_module/_08776_ ;
 wire \reg_module/_08777_ ;
 wire \reg_module/_08778_ ;
 wire \reg_module/_08779_ ;
 wire \reg_module/_08780_ ;
 wire \reg_module/_08781_ ;
 wire \reg_module/_08782_ ;
 wire \reg_module/_08783_ ;
 wire \reg_module/_08784_ ;
 wire \reg_module/_08785_ ;
 wire \reg_module/_08786_ ;
 wire \reg_module/_08787_ ;
 wire \reg_module/_08788_ ;
 wire \reg_module/_08789_ ;
 wire \reg_module/_08790_ ;
 wire \reg_module/_08791_ ;
 wire \reg_module/_08792_ ;
 wire \reg_module/_08793_ ;
 wire \reg_module/_08794_ ;
 wire \reg_module/_08795_ ;
 wire \reg_module/_08796_ ;
 wire \reg_module/_08797_ ;
 wire \reg_module/_08798_ ;
 wire \reg_module/_08799_ ;
 wire \reg_module/_08800_ ;
 wire \reg_module/_08801_ ;
 wire \reg_module/_08802_ ;
 wire \reg_module/_08803_ ;
 wire \reg_module/_08804_ ;
 wire \reg_module/_08805_ ;
 wire \reg_module/_08806_ ;
 wire \reg_module/_08807_ ;
 wire \reg_module/_08808_ ;
 wire \reg_module/_08809_ ;
 wire \reg_module/_08810_ ;
 wire \reg_module/_08811_ ;
 wire \reg_module/_08812_ ;
 wire \reg_module/_08813_ ;
 wire \reg_module/_08814_ ;
 wire \reg_module/_08815_ ;
 wire \reg_module/_08816_ ;
 wire \reg_module/_08817_ ;
 wire \reg_module/_08818_ ;
 wire \reg_module/_08819_ ;
 wire \reg_module/_08820_ ;
 wire \reg_module/_08821_ ;
 wire \reg_module/_08822_ ;
 wire \reg_module/_08823_ ;
 wire \reg_module/_08824_ ;
 wire \reg_module/_08825_ ;
 wire \reg_module/_08826_ ;
 wire \reg_module/_08827_ ;
 wire \reg_module/_08828_ ;
 wire \reg_module/_08829_ ;
 wire \reg_module/_08830_ ;
 wire \reg_module/_08831_ ;
 wire \reg_module/_08832_ ;
 wire \reg_module/_08833_ ;
 wire \reg_module/_08834_ ;
 wire \reg_module/_08835_ ;
 wire \reg_module/_08836_ ;
 wire \reg_module/_08837_ ;
 wire \reg_module/_08838_ ;
 wire \reg_module/_08839_ ;
 wire \reg_module/_08840_ ;
 wire \reg_module/_08841_ ;
 wire \reg_module/_08842_ ;
 wire \reg_module/_08843_ ;
 wire \reg_module/_08844_ ;
 wire \reg_module/_08845_ ;
 wire \reg_module/_08846_ ;
 wire \reg_module/_08847_ ;
 wire \reg_module/_08848_ ;
 wire \reg_module/_08849_ ;
 wire \reg_module/_08850_ ;
 wire \reg_module/_08851_ ;
 wire \reg_module/_08852_ ;
 wire \reg_module/_08853_ ;
 wire \reg_module/_08854_ ;
 wire \reg_module/_08855_ ;
 wire \reg_module/_08856_ ;
 wire \reg_module/_08857_ ;
 wire \reg_module/_08858_ ;
 wire \reg_module/_08859_ ;
 wire \reg_module/_08860_ ;
 wire \reg_module/_08861_ ;
 wire \reg_module/_08862_ ;
 wire \reg_module/_08863_ ;
 wire \reg_module/_08864_ ;
 wire \reg_module/_08865_ ;
 wire \reg_module/_08866_ ;
 wire \reg_module/_08867_ ;
 wire \reg_module/_08868_ ;
 wire \reg_module/_08869_ ;
 wire \reg_module/_08870_ ;
 wire \reg_module/_08871_ ;
 wire \reg_module/_08872_ ;
 wire \reg_module/_08873_ ;
 wire \reg_module/_08874_ ;
 wire \reg_module/_08875_ ;
 wire \reg_module/_08876_ ;
 wire \reg_module/_08877_ ;
 wire \reg_module/_08878_ ;
 wire \reg_module/_08879_ ;
 wire \reg_module/_08880_ ;
 wire \reg_module/_08881_ ;
 wire \reg_module/_08882_ ;
 wire \reg_module/_08883_ ;
 wire \reg_module/_08884_ ;
 wire \reg_module/_08885_ ;
 wire \reg_module/_08886_ ;
 wire \reg_module/_08887_ ;
 wire \reg_module/_08888_ ;
 wire \reg_module/_08889_ ;
 wire \reg_module/_08890_ ;
 wire \reg_module/_08891_ ;
 wire \reg_module/_08892_ ;
 wire \reg_module/_08893_ ;
 wire \reg_module/_08894_ ;
 wire \reg_module/_08895_ ;
 wire \reg_module/_08896_ ;
 wire \reg_module/_08897_ ;
 wire \reg_module/_08898_ ;
 wire \reg_module/_08899_ ;
 wire \reg_module/_08900_ ;
 wire \reg_module/_08901_ ;
 wire \reg_module/_08902_ ;
 wire \reg_module/_08903_ ;
 wire \reg_module/_08904_ ;
 wire \reg_module/_08905_ ;
 wire \reg_module/_08906_ ;
 wire \reg_module/_08907_ ;
 wire \reg_module/_08908_ ;
 wire \reg_module/_08909_ ;
 wire \reg_module/_08910_ ;
 wire \reg_module/_08911_ ;
 wire \reg_module/_08912_ ;
 wire \reg_module/_08913_ ;
 wire \reg_module/_08914_ ;
 wire \reg_module/_08915_ ;
 wire \reg_module/_08916_ ;
 wire \reg_module/_08917_ ;
 wire \reg_module/_08918_ ;
 wire \reg_module/_08919_ ;
 wire \reg_module/_08920_ ;
 wire \reg_module/_08921_ ;
 wire \reg_module/_08922_ ;
 wire \reg_module/_08923_ ;
 wire \reg_module/_08924_ ;
 wire \reg_module/_08925_ ;
 wire \reg_module/_08926_ ;
 wire \reg_module/_08927_ ;
 wire \reg_module/_08928_ ;
 wire \reg_module/_08929_ ;
 wire \reg_module/_08930_ ;
 wire \reg_module/_08931_ ;
 wire \reg_module/_08932_ ;
 wire \reg_module/_08933_ ;
 wire \reg_module/_08934_ ;
 wire \reg_module/_08935_ ;
 wire \reg_module/_08936_ ;
 wire \reg_module/_08937_ ;
 wire \reg_module/_08938_ ;
 wire \reg_module/_08939_ ;
 wire \reg_module/_08940_ ;
 wire \reg_module/_08941_ ;
 wire \reg_module/_08942_ ;
 wire \reg_module/_08943_ ;
 wire \reg_module/_08944_ ;
 wire \reg_module/_08945_ ;
 wire \reg_module/_08946_ ;
 wire \reg_module/_08947_ ;
 wire \reg_module/_08948_ ;
 wire \reg_module/_08949_ ;
 wire \reg_module/_08950_ ;
 wire \reg_module/_08951_ ;
 wire \reg_module/_08952_ ;
 wire \reg_module/_08953_ ;
 wire \reg_module/_08954_ ;
 wire \reg_module/_08955_ ;
 wire \reg_module/_08956_ ;
 wire \reg_module/_08957_ ;
 wire \reg_module/_08958_ ;
 wire \reg_module/_08959_ ;
 wire \reg_module/_08960_ ;
 wire \reg_module/_08961_ ;
 wire \reg_module/_08962_ ;
 wire \reg_module/_08963_ ;
 wire \reg_module/_08964_ ;
 wire \reg_module/_08965_ ;
 wire \reg_module/_08966_ ;
 wire \reg_module/_08967_ ;
 wire \reg_module/_08968_ ;
 wire \reg_module/_08969_ ;
 wire \reg_module/_08970_ ;
 wire \reg_module/_08971_ ;
 wire \reg_module/_08972_ ;
 wire \reg_module/_08973_ ;
 wire \reg_module/_08974_ ;
 wire \reg_module/_08975_ ;
 wire \reg_module/_08976_ ;
 wire \reg_module/_08977_ ;
 wire \reg_module/_08978_ ;
 wire \reg_module/_08979_ ;
 wire \reg_module/_08980_ ;
 wire \reg_module/_08981_ ;
 wire \reg_module/_08982_ ;
 wire \reg_module/_08983_ ;
 wire \reg_module/_08984_ ;
 wire \reg_module/_08985_ ;
 wire \reg_module/_08986_ ;
 wire \reg_module/_08987_ ;
 wire \reg_module/_08988_ ;
 wire \reg_module/_08989_ ;
 wire \reg_module/_08990_ ;
 wire \reg_module/_08991_ ;
 wire \reg_module/_08992_ ;
 wire \reg_module/_08993_ ;
 wire \reg_module/_08994_ ;
 wire \reg_module/_08995_ ;
 wire \reg_module/_08996_ ;
 wire \reg_module/_08997_ ;
 wire \reg_module/_08998_ ;
 wire \reg_module/_08999_ ;
 wire \reg_module/_09000_ ;
 wire \reg_module/_09001_ ;
 wire \reg_module/_09002_ ;
 wire \reg_module/_09003_ ;
 wire \reg_module/_09004_ ;
 wire \reg_module/_09005_ ;
 wire \reg_module/_09006_ ;
 wire \reg_module/_09007_ ;
 wire \reg_module/_09008_ ;
 wire \reg_module/_09009_ ;
 wire \reg_module/_09010_ ;
 wire \reg_module/_09011_ ;
 wire \reg_module/_09012_ ;
 wire \reg_module/_09013_ ;
 wire \reg_module/_09014_ ;
 wire \reg_module/_09015_ ;
 wire \reg_module/_09016_ ;
 wire \reg_module/_09017_ ;
 wire \reg_module/_09018_ ;
 wire \reg_module/_09019_ ;
 wire \reg_module/_09020_ ;
 wire \reg_module/_09021_ ;
 wire \reg_module/_09022_ ;
 wire \reg_module/_09023_ ;
 wire \reg_module/_09024_ ;
 wire \reg_module/_09025_ ;
 wire \reg_module/_09026_ ;
 wire \reg_module/_09027_ ;
 wire \reg_module/_09028_ ;
 wire \reg_module/_09029_ ;
 wire \reg_module/_09030_ ;
 wire \reg_module/_09031_ ;
 wire \reg_module/_09032_ ;
 wire \reg_module/_09033_ ;
 wire \reg_module/_09034_ ;
 wire \reg_module/_09035_ ;
 wire \reg_module/_09036_ ;
 wire \reg_module/_09037_ ;
 wire \reg_module/_09038_ ;
 wire \reg_module/_09039_ ;
 wire \reg_module/_09040_ ;
 wire \reg_module/_09041_ ;
 wire \reg_module/_09042_ ;
 wire \reg_module/_09043_ ;
 wire \reg_module/_09044_ ;
 wire \reg_module/_09045_ ;
 wire \reg_module/_09046_ ;
 wire \reg_module/_09047_ ;
 wire \reg_module/_09048_ ;
 wire \reg_module/_09049_ ;
 wire \reg_module/_09050_ ;
 wire \reg_module/_09051_ ;
 wire \reg_module/_09052_ ;
 wire \reg_module/_09053_ ;
 wire \reg_module/_09054_ ;
 wire \reg_module/_09055_ ;
 wire \reg_module/_09056_ ;
 wire \reg_module/_09057_ ;
 wire \reg_module/_09058_ ;
 wire \reg_module/_09059_ ;
 wire \reg_module/_09060_ ;
 wire \reg_module/_09061_ ;
 wire \reg_module/_09062_ ;
 wire \reg_module/_09063_ ;
 wire \reg_module/_09064_ ;
 wire \reg_module/_09065_ ;
 wire \reg_module/_09066_ ;
 wire \reg_module/_09067_ ;
 wire \reg_module/_09068_ ;
 wire \reg_module/_09069_ ;
 wire \reg_module/_09070_ ;
 wire \reg_module/_09071_ ;
 wire \reg_module/_09072_ ;
 wire \reg_module/_09073_ ;
 wire \reg_module/_09074_ ;
 wire \reg_module/_09075_ ;
 wire \reg_module/_09076_ ;
 wire \reg_module/_09077_ ;
 wire \reg_module/_09078_ ;
 wire \reg_module/_09079_ ;
 wire \reg_module/_09080_ ;
 wire \reg_module/_09081_ ;
 wire \reg_module/_09082_ ;
 wire \reg_module/_09083_ ;
 wire \reg_module/_09084_ ;
 wire \reg_module/_09085_ ;
 wire \reg_module/_09086_ ;
 wire \reg_module/_09087_ ;
 wire \reg_module/_09088_ ;
 wire \reg_module/_09089_ ;
 wire \reg_module/_09090_ ;
 wire \reg_module/_09091_ ;
 wire \reg_module/_09092_ ;
 wire \reg_module/_09093_ ;
 wire \reg_module/_09094_ ;
 wire \reg_module/_09095_ ;
 wire \reg_module/_09096_ ;
 wire \reg_module/_09097_ ;
 wire \reg_module/_09098_ ;
 wire \reg_module/_09099_ ;
 wire \reg_module/_09100_ ;
 wire \reg_module/_09101_ ;
 wire \reg_module/_09102_ ;
 wire \reg_module/_09103_ ;
 wire \reg_module/_09104_ ;
 wire \reg_module/_09105_ ;
 wire \reg_module/_09106_ ;
 wire \reg_module/_09107_ ;
 wire \reg_module/_09108_ ;
 wire \reg_module/_09109_ ;
 wire \reg_module/_09110_ ;
 wire \reg_module/_09111_ ;
 wire \reg_module/_09112_ ;
 wire \reg_module/_09113_ ;
 wire \reg_module/_09114_ ;
 wire \reg_module/_09115_ ;
 wire \reg_module/_09116_ ;
 wire \reg_module/_09117_ ;
 wire \reg_module/_09118_ ;
 wire \reg_module/_09119_ ;
 wire \reg_module/_09120_ ;
 wire \reg_module/_09121_ ;
 wire \reg_module/_09122_ ;
 wire \reg_module/_09123_ ;
 wire \reg_module/_09124_ ;
 wire \reg_module/_09125_ ;
 wire \reg_module/_09126_ ;
 wire \reg_module/_09127_ ;
 wire \reg_module/_09128_ ;
 wire \reg_module/_09129_ ;
 wire \reg_module/_09130_ ;
 wire \reg_module/_09131_ ;
 wire \reg_module/_09132_ ;
 wire \reg_module/_09133_ ;
 wire \reg_module/_09134_ ;
 wire \reg_module/_09135_ ;
 wire \reg_module/_09136_ ;
 wire \reg_module/_09137_ ;
 wire \reg_module/_09138_ ;
 wire \reg_module/_09139_ ;
 wire \reg_module/_09140_ ;
 wire \reg_module/_09141_ ;
 wire \reg_module/_09142_ ;
 wire \reg_module/_09143_ ;
 wire \reg_module/_09144_ ;
 wire \reg_module/_09145_ ;
 wire \reg_module/_09146_ ;
 wire \reg_module/_09147_ ;
 wire \reg_module/_09148_ ;
 wire \reg_module/_09149_ ;
 wire \reg_module/_09150_ ;
 wire \reg_module/_09151_ ;
 wire \reg_module/_09152_ ;
 wire \reg_module/_09153_ ;
 wire \reg_module/_09154_ ;
 wire \reg_module/_09155_ ;
 wire \reg_module/_09156_ ;
 wire \reg_module/_09157_ ;
 wire \reg_module/_09158_ ;
 wire \reg_module/_09159_ ;
 wire \reg_module/_09160_ ;
 wire \reg_module/_09161_ ;
 wire \reg_module/_09162_ ;
 wire \reg_module/_09163_ ;
 wire \reg_module/_09164_ ;
 wire \reg_module/_09165_ ;
 wire \reg_module/_09166_ ;
 wire \reg_module/_09167_ ;
 wire \reg_module/_09168_ ;
 wire \reg_module/_09169_ ;
 wire \reg_module/_09170_ ;
 wire \reg_module/_09171_ ;
 wire \reg_module/_09172_ ;
 wire \reg_module/_09173_ ;
 wire \reg_module/_09174_ ;
 wire \reg_module/_09175_ ;
 wire \reg_module/_09176_ ;
 wire \reg_module/_09177_ ;
 wire \reg_module/_09178_ ;
 wire \reg_module/_09179_ ;
 wire \reg_module/_09180_ ;
 wire \reg_module/_09181_ ;
 wire \reg_module/_09182_ ;
 wire \reg_module/_09183_ ;
 wire \reg_module/_09184_ ;
 wire \reg_module/_09185_ ;
 wire \reg_module/_09186_ ;
 wire \reg_module/_09187_ ;
 wire \reg_module/_09188_ ;
 wire \reg_module/_09189_ ;
 wire \reg_module/_09190_ ;
 wire \reg_module/_09191_ ;
 wire \reg_module/_09192_ ;
 wire \reg_module/_09193_ ;
 wire \reg_module/_09194_ ;
 wire \reg_module/_09195_ ;
 wire \reg_module/_09196_ ;
 wire \reg_module/_09197_ ;
 wire \reg_module/_09198_ ;
 wire \reg_module/_09199_ ;
 wire \reg_module/_09200_ ;
 wire \reg_module/_09201_ ;
 wire \reg_module/_09202_ ;
 wire \reg_module/_09203_ ;
 wire \reg_module/_09204_ ;
 wire \reg_module/_09205_ ;
 wire \reg_module/_09206_ ;
 wire \reg_module/_09207_ ;
 wire \reg_module/_09208_ ;
 wire \reg_module/_09209_ ;
 wire \reg_module/_09210_ ;
 wire \reg_module/_09211_ ;
 wire \reg_module/_09212_ ;
 wire \reg_module/_09213_ ;
 wire \reg_module/_09214_ ;
 wire \reg_module/_09215_ ;
 wire \reg_module/_09216_ ;
 wire \reg_module/_09217_ ;
 wire \reg_module/_09218_ ;
 wire \reg_module/_09219_ ;
 wire \reg_module/_09220_ ;
 wire \reg_module/_09221_ ;
 wire \reg_module/_09222_ ;
 wire \reg_module/_09223_ ;
 wire \reg_module/_09224_ ;
 wire \reg_module/_09225_ ;
 wire \reg_module/_09226_ ;
 wire \reg_module/_09227_ ;
 wire \reg_module/_09228_ ;
 wire \reg_module/_09229_ ;
 wire \reg_module/_09230_ ;
 wire \reg_module/_09231_ ;
 wire \reg_module/_09232_ ;
 wire \reg_module/_09233_ ;
 wire \reg_module/_09234_ ;
 wire \reg_module/_09235_ ;
 wire \reg_module/_09236_ ;
 wire \reg_module/_09237_ ;
 wire \reg_module/_09238_ ;
 wire \reg_module/_09239_ ;
 wire \reg_module/_09240_ ;
 wire \reg_module/_09241_ ;
 wire \reg_module/_09242_ ;
 wire \reg_module/_09243_ ;
 wire \reg_module/_09244_ ;
 wire \reg_module/_09245_ ;
 wire \reg_module/_09246_ ;
 wire \reg_module/_09247_ ;
 wire \reg_module/_09248_ ;
 wire \reg_module/_09249_ ;
 wire \reg_module/_09250_ ;
 wire \reg_module/_09251_ ;
 wire \reg_module/_09252_ ;
 wire \reg_module/_09253_ ;
 wire \reg_module/_09254_ ;
 wire \reg_module/_09255_ ;
 wire \reg_module/_09256_ ;
 wire \reg_module/_09257_ ;
 wire \reg_module/_09258_ ;
 wire \reg_module/_09259_ ;
 wire \reg_module/_09260_ ;
 wire \reg_module/_09261_ ;
 wire \reg_module/_09262_ ;
 wire \reg_module/_09263_ ;
 wire \reg_module/_09264_ ;
 wire \reg_module/_09265_ ;
 wire \reg_module/_09266_ ;
 wire \reg_module/_09267_ ;
 wire \reg_module/_09268_ ;
 wire \reg_module/_09269_ ;
 wire \reg_module/_09270_ ;
 wire \reg_module/_09271_ ;
 wire \reg_module/_09272_ ;
 wire \reg_module/_09273_ ;
 wire \reg_module/_09274_ ;
 wire \reg_module/_09275_ ;
 wire \reg_module/_09276_ ;
 wire \reg_module/_09277_ ;
 wire \reg_module/_09278_ ;
 wire \reg_module/_09279_ ;
 wire \reg_module/_09280_ ;
 wire \reg_module/_09281_ ;
 wire \reg_module/_09282_ ;
 wire \reg_module/_09283_ ;
 wire \reg_module/_09284_ ;
 wire \reg_module/_09285_ ;
 wire \reg_module/_09286_ ;
 wire \reg_module/_09287_ ;
 wire \reg_module/_09288_ ;
 wire \reg_module/_09289_ ;
 wire \reg_module/_09290_ ;
 wire \reg_module/_09291_ ;
 wire \reg_module/_09292_ ;
 wire \reg_module/_09293_ ;
 wire \reg_module/_09294_ ;
 wire \reg_module/_09295_ ;
 wire \reg_module/_09296_ ;
 wire \reg_module/_09297_ ;
 wire \reg_module/_09298_ ;
 wire \reg_module/_09299_ ;
 wire \reg_module/_09300_ ;
 wire \reg_module/_09301_ ;
 wire \reg_module/_09302_ ;
 wire \reg_module/_09303_ ;
 wire \reg_module/_09304_ ;
 wire \reg_module/_09305_ ;
 wire \reg_module/_09306_ ;
 wire \reg_module/_09307_ ;
 wire \reg_module/_09308_ ;
 wire \reg_module/_09309_ ;
 wire \reg_module/_09310_ ;
 wire \reg_module/_09311_ ;
 wire \reg_module/_09312_ ;
 wire \reg_module/_09313_ ;
 wire \reg_module/_09314_ ;
 wire \reg_module/_09315_ ;
 wire \reg_module/_09316_ ;
 wire \reg_module/_09317_ ;
 wire \reg_module/_09318_ ;
 wire \reg_module/_09319_ ;
 wire \reg_module/_09320_ ;
 wire \reg_module/_09321_ ;
 wire \reg_module/_09322_ ;
 wire \reg_module/_09323_ ;
 wire \reg_module/_09324_ ;
 wire \reg_module/_09325_ ;
 wire \reg_module/_09326_ ;
 wire \reg_module/_09327_ ;
 wire \reg_module/_09328_ ;
 wire \reg_module/_09329_ ;
 wire \reg_module/_09330_ ;
 wire \reg_module/_09331_ ;
 wire \reg_module/_09332_ ;
 wire \reg_module/_09333_ ;
 wire \reg_module/_09334_ ;
 wire \reg_module/_09335_ ;
 wire \reg_module/_09336_ ;
 wire \reg_module/_09337_ ;
 wire \reg_module/_09338_ ;
 wire \reg_module/_09339_ ;
 wire \reg_module/_09340_ ;
 wire \reg_module/_09341_ ;
 wire \reg_module/_09342_ ;
 wire \reg_module/_09343_ ;
 wire \reg_module/_09344_ ;
 wire \reg_module/_09345_ ;
 wire \reg_module/_09346_ ;
 wire \reg_module/_09347_ ;
 wire \reg_module/_09348_ ;
 wire \reg_module/_09349_ ;
 wire \reg_module/_09350_ ;
 wire \reg_module/_09351_ ;
 wire \reg_module/_09352_ ;
 wire \reg_module/_09353_ ;
 wire \reg_module/_09354_ ;
 wire \reg_module/_09355_ ;
 wire \reg_module/_09356_ ;
 wire \reg_module/_09357_ ;
 wire \reg_module/_09358_ ;
 wire \reg_module/_09359_ ;
 wire \reg_module/_09360_ ;
 wire \reg_module/_09361_ ;
 wire \reg_module/_09362_ ;
 wire \reg_module/_09363_ ;
 wire \reg_module/_09364_ ;
 wire \reg_module/_09365_ ;
 wire \reg_module/_09366_ ;
 wire \reg_module/_09367_ ;
 wire \reg_module/_09368_ ;
 wire \reg_module/_09369_ ;
 wire \reg_module/_09370_ ;
 wire \reg_module/_09371_ ;
 wire \reg_module/_09372_ ;
 wire \reg_module/_09373_ ;
 wire \reg_module/_09374_ ;
 wire \reg_module/_09375_ ;
 wire \reg_module/_09376_ ;
 wire \reg_module/_09377_ ;
 wire \reg_module/_09378_ ;
 wire \reg_module/_09379_ ;
 wire \reg_module/_09380_ ;
 wire \reg_module/_09381_ ;
 wire \reg_module/_09382_ ;
 wire \reg_module/_09383_ ;
 wire \reg_module/_09384_ ;
 wire \reg_module/_09385_ ;
 wire \reg_module/_09386_ ;
 wire \reg_module/_09387_ ;
 wire \reg_module/_09388_ ;
 wire \reg_module/_09389_ ;
 wire \reg_module/_09390_ ;
 wire \reg_module/_09391_ ;
 wire \reg_module/_09392_ ;
 wire \reg_module/_09393_ ;
 wire \reg_module/_09394_ ;
 wire \reg_module/_09395_ ;
 wire \reg_module/_09396_ ;
 wire \reg_module/_09397_ ;
 wire \reg_module/_09398_ ;
 wire \reg_module/_09399_ ;
 wire \reg_module/_09400_ ;
 wire \reg_module/_09401_ ;
 wire \reg_module/_09402_ ;
 wire \reg_module/_09403_ ;
 wire \reg_module/_09404_ ;
 wire \reg_module/_09405_ ;
 wire \reg_module/_09406_ ;
 wire \reg_module/_09407_ ;
 wire \reg_module/_09408_ ;
 wire \reg_module/_09409_ ;
 wire \reg_module/_09410_ ;
 wire \reg_module/_09411_ ;
 wire \reg_module/_09412_ ;
 wire \reg_module/_09413_ ;
 wire \reg_module/_09414_ ;
 wire \reg_module/_09415_ ;
 wire \reg_module/_09416_ ;
 wire \reg_module/_09417_ ;
 wire \reg_module/_09418_ ;
 wire \reg_module/_09419_ ;
 wire \reg_module/_09420_ ;
 wire \reg_module/_09421_ ;
 wire \reg_module/_09422_ ;
 wire \reg_module/_09423_ ;
 wire \reg_module/_09424_ ;
 wire \reg_module/_09425_ ;
 wire \reg_module/_09426_ ;
 wire \reg_module/_09427_ ;
 wire \reg_module/_09428_ ;
 wire \reg_module/_09429_ ;
 wire \reg_module/_09430_ ;
 wire \reg_module/_09431_ ;
 wire \reg_module/_09432_ ;
 wire \reg_module/_09433_ ;
 wire \reg_module/_09434_ ;
 wire \reg_module/_09435_ ;
 wire \reg_module/_09436_ ;
 wire \reg_module/_09437_ ;
 wire \reg_module/_09438_ ;
 wire \reg_module/_09439_ ;
 wire \reg_module/_09440_ ;
 wire \reg_module/_09441_ ;
 wire \reg_module/_09442_ ;
 wire \reg_module/_09443_ ;
 wire \reg_module/_09444_ ;
 wire \reg_module/_09445_ ;
 wire \reg_module/_09446_ ;
 wire \reg_module/_09447_ ;
 wire \reg_module/_09448_ ;
 wire \reg_module/_09449_ ;
 wire \reg_module/_09450_ ;
 wire \reg_module/_09451_ ;
 wire \reg_module/_09452_ ;
 wire \reg_module/_09453_ ;
 wire \reg_module/_09454_ ;
 wire \reg_module/_09455_ ;
 wire \reg_module/_09456_ ;
 wire \reg_module/_09457_ ;
 wire \reg_module/_09458_ ;
 wire \reg_module/_09459_ ;
 wire \reg_module/_09460_ ;
 wire \reg_module/_09461_ ;
 wire \reg_module/_09462_ ;
 wire \reg_module/_09463_ ;
 wire \reg_module/_09464_ ;
 wire \reg_module/_09465_ ;
 wire \reg_module/_09466_ ;
 wire \reg_module/_09467_ ;
 wire \reg_module/_09468_ ;
 wire \reg_module/_09469_ ;
 wire \reg_module/_09470_ ;
 wire \reg_module/_09471_ ;
 wire \reg_module/_09472_ ;
 wire \reg_module/_09473_ ;
 wire \reg_module/_09474_ ;
 wire \reg_module/_09475_ ;
 wire \reg_module/_09476_ ;
 wire \reg_module/_09477_ ;
 wire \reg_module/_09478_ ;
 wire \reg_module/_09479_ ;
 wire \reg_module/_09480_ ;
 wire \reg_module/_09481_ ;
 wire \reg_module/_09482_ ;
 wire \reg_module/_09483_ ;
 wire \reg_module/_09484_ ;
 wire \reg_module/_09485_ ;
 wire \reg_module/_09486_ ;
 wire \reg_module/_09487_ ;
 wire \reg_module/_09488_ ;
 wire \reg_module/_09489_ ;
 wire \reg_module/_09490_ ;
 wire \reg_module/_09491_ ;
 wire \reg_module/_09492_ ;
 wire \reg_module/_09493_ ;
 wire \reg_module/_09494_ ;
 wire \reg_module/_09495_ ;
 wire \reg_module/_09496_ ;
 wire \reg_module/_09497_ ;
 wire \reg_module/_09498_ ;
 wire \reg_module/_09499_ ;
 wire \reg_module/_09500_ ;
 wire \reg_module/_09501_ ;
 wire \reg_module/_09502_ ;
 wire \reg_module/_09503_ ;
 wire \reg_module/_09504_ ;
 wire \reg_module/_09505_ ;
 wire \reg_module/_09506_ ;
 wire \reg_module/_09507_ ;
 wire \reg_module/_09508_ ;
 wire \reg_module/_09509_ ;
 wire \reg_module/_09510_ ;
 wire \reg_module/_09511_ ;
 wire \reg_module/_09512_ ;
 wire \reg_module/_09513_ ;
 wire \reg_module/_09514_ ;
 wire \reg_module/_09515_ ;
 wire \reg_module/_09516_ ;
 wire \reg_module/_09517_ ;
 wire \reg_module/_09518_ ;
 wire \reg_module/_09519_ ;
 wire \reg_module/_09520_ ;
 wire \reg_module/_09521_ ;
 wire \reg_module/_09522_ ;
 wire \reg_module/_09523_ ;
 wire \reg_module/_09524_ ;
 wire \reg_module/_09525_ ;
 wire \reg_module/_09526_ ;
 wire \reg_module/_09527_ ;
 wire \reg_module/_09528_ ;
 wire \reg_module/_09529_ ;
 wire \reg_module/_09530_ ;
 wire \reg_module/_09531_ ;
 wire \reg_module/_09532_ ;
 wire \reg_module/_09533_ ;
 wire \reg_module/_09534_ ;
 wire \reg_module/_09535_ ;
 wire \reg_module/_09536_ ;
 wire \reg_module/_09537_ ;
 wire \reg_module/_09538_ ;
 wire \reg_module/_09539_ ;
 wire \reg_module/_09540_ ;
 wire \reg_module/_09541_ ;
 wire \reg_module/_09542_ ;
 wire \reg_module/_09543_ ;
 wire \reg_module/_09544_ ;
 wire \reg_module/_09545_ ;
 wire \reg_module/_09546_ ;
 wire \reg_module/_09547_ ;
 wire \reg_module/_09548_ ;
 wire \reg_module/_09549_ ;
 wire \reg_module/_09550_ ;
 wire \reg_module/_09551_ ;
 wire \reg_module/_09552_ ;
 wire \reg_module/_09553_ ;
 wire \reg_module/_09554_ ;
 wire \reg_module/_09555_ ;
 wire \reg_module/_09556_ ;
 wire \reg_module/_09557_ ;
 wire \reg_module/_09558_ ;
 wire \reg_module/_09559_ ;
 wire \reg_module/_09560_ ;
 wire \reg_module/_09561_ ;
 wire \reg_module/_09562_ ;
 wire \reg_module/_09563_ ;
 wire \reg_module/_09564_ ;
 wire \reg_module/_09565_ ;
 wire \reg_module/_09566_ ;
 wire \reg_module/_09567_ ;
 wire \reg_module/_09568_ ;
 wire \reg_module/_09569_ ;
 wire \reg_module/_09570_ ;
 wire \reg_module/_09571_ ;
 wire \reg_module/_09572_ ;
 wire \reg_module/_09573_ ;
 wire \reg_module/_09574_ ;
 wire \reg_module/_09575_ ;
 wire \reg_module/_09576_ ;
 wire \reg_module/_09577_ ;
 wire \reg_module/_09578_ ;
 wire \reg_module/_09579_ ;
 wire \reg_module/_09580_ ;
 wire \reg_module/_09581_ ;
 wire \reg_module/_09582_ ;
 wire \reg_module/_09583_ ;
 wire \reg_module/_09584_ ;
 wire \reg_module/_09585_ ;
 wire \reg_module/_09586_ ;
 wire \reg_module/_09587_ ;
 wire \reg_module/_09588_ ;
 wire \reg_module/_09589_ ;
 wire \reg_module/_09590_ ;
 wire \reg_module/_09591_ ;
 wire \reg_module/_09592_ ;
 wire \reg_module/_09593_ ;
 wire \reg_module/_09594_ ;
 wire \reg_module/_09595_ ;
 wire \reg_module/_09596_ ;
 wire \reg_module/_09597_ ;
 wire \reg_module/_09598_ ;
 wire \reg_module/_09599_ ;
 wire \reg_module/_09600_ ;
 wire \reg_module/_09601_ ;
 wire \reg_module/_09602_ ;
 wire \reg_module/_09603_ ;
 wire \reg_module/_09604_ ;
 wire \reg_module/_09605_ ;
 wire \reg_module/_09606_ ;
 wire \reg_module/_09607_ ;
 wire \reg_module/_09608_ ;
 wire \reg_module/_09609_ ;
 wire \reg_module/_09610_ ;
 wire \reg_module/_09611_ ;
 wire \reg_module/_09612_ ;
 wire \reg_module/_09613_ ;
 wire \reg_module/_09614_ ;
 wire \reg_module/_09615_ ;
 wire \reg_module/_09616_ ;
 wire \reg_module/_09617_ ;
 wire \reg_module/_09618_ ;
 wire \reg_module/_09619_ ;
 wire \reg_module/_09620_ ;
 wire \reg_module/_09621_ ;
 wire \reg_module/_09622_ ;
 wire \reg_module/_09623_ ;
 wire \reg_module/_09624_ ;
 wire \reg_module/_09625_ ;
 wire \reg_module/_09626_ ;
 wire \reg_module/_09627_ ;
 wire \reg_module/_09628_ ;
 wire \reg_module/_09629_ ;
 wire \reg_module/_09630_ ;
 wire \reg_module/_09631_ ;
 wire \reg_module/_09632_ ;
 wire \reg_module/_09633_ ;
 wire \reg_module/_09634_ ;
 wire \reg_module/_09635_ ;
 wire \reg_module/_09636_ ;
 wire \reg_module/_09637_ ;
 wire \reg_module/_09638_ ;
 wire \reg_module/_09639_ ;
 wire \reg_module/_09640_ ;
 wire \reg_module/_09641_ ;
 wire \reg_module/_09642_ ;
 wire \reg_module/_09643_ ;
 wire \reg_module/_09644_ ;
 wire \reg_module/_09645_ ;
 wire \reg_module/_09646_ ;
 wire \reg_module/_09647_ ;
 wire \reg_module/_09648_ ;
 wire \reg_module/_09649_ ;
 wire \reg_module/_09650_ ;
 wire \reg_module/_09651_ ;
 wire \reg_module/_09652_ ;
 wire \reg_module/_09653_ ;
 wire \reg_module/_09654_ ;
 wire \reg_module/_09655_ ;
 wire \reg_module/_09656_ ;
 wire \reg_module/_09657_ ;
 wire \reg_module/_09658_ ;
 wire \reg_module/_09659_ ;
 wire \reg_module/_09660_ ;
 wire \reg_module/_09661_ ;
 wire \reg_module/_09662_ ;
 wire \reg_module/_09663_ ;
 wire \reg_module/_09664_ ;
 wire \reg_module/_09665_ ;
 wire \reg_module/_09666_ ;
 wire \reg_module/_09667_ ;
 wire \reg_module/_09668_ ;
 wire \reg_module/_09669_ ;
 wire \reg_module/_09670_ ;
 wire \reg_module/_09671_ ;
 wire \reg_module/_09672_ ;
 wire \reg_module/_09673_ ;
 wire \reg_module/_09674_ ;
 wire \reg_module/_09675_ ;
 wire \reg_module/_09676_ ;
 wire \reg_module/_09677_ ;
 wire \reg_module/_09678_ ;
 wire \reg_module/_09679_ ;
 wire \reg_module/_09680_ ;
 wire \reg_module/_09681_ ;
 wire \reg_module/_09682_ ;
 wire \reg_module/_09683_ ;
 wire \reg_module/_09684_ ;
 wire \reg_module/_09685_ ;
 wire \reg_module/_09686_ ;
 wire \reg_module/_09687_ ;
 wire \reg_module/_09688_ ;
 wire \reg_module/_09689_ ;
 wire \reg_module/_09690_ ;
 wire \reg_module/_09691_ ;
 wire \reg_module/_09692_ ;
 wire \reg_module/_09693_ ;
 wire \reg_module/_09694_ ;
 wire \reg_module/_09695_ ;
 wire \reg_module/_09696_ ;
 wire \reg_module/_09697_ ;
 wire \reg_module/_09698_ ;
 wire \reg_module/_09699_ ;
 wire \reg_module/_09700_ ;
 wire \reg_module/_09701_ ;
 wire \reg_module/_09702_ ;
 wire \reg_module/_09703_ ;
 wire \reg_module/_09704_ ;
 wire \reg_module/_09705_ ;
 wire \reg_module/_09706_ ;
 wire \reg_module/_09707_ ;
 wire \reg_module/_09708_ ;
 wire \reg_module/_09709_ ;
 wire \reg_module/_09710_ ;
 wire \reg_module/_09711_ ;
 wire \reg_module/_09712_ ;
 wire \reg_module/_09713_ ;
 wire \reg_module/_09714_ ;
 wire \reg_module/_09715_ ;
 wire \reg_module/_09716_ ;
 wire \reg_module/_09717_ ;
 wire \reg_module/_09718_ ;
 wire \reg_module/_09719_ ;
 wire \reg_module/_09720_ ;
 wire \reg_module/_09721_ ;
 wire \reg_module/_09722_ ;
 wire \reg_module/_09723_ ;
 wire \reg_module/_09724_ ;
 wire \reg_module/_09725_ ;
 wire \reg_module/_09726_ ;
 wire \reg_module/_09727_ ;
 wire \reg_module/_09728_ ;
 wire \reg_module/_09729_ ;
 wire \reg_module/_09730_ ;
 wire \reg_module/_09731_ ;
 wire \reg_module/_09732_ ;
 wire \reg_module/_09733_ ;
 wire \reg_module/_09734_ ;
 wire \reg_module/_09735_ ;
 wire \reg_module/_09736_ ;
 wire \reg_module/_09737_ ;
 wire \reg_module/_09738_ ;
 wire \reg_module/_09739_ ;
 wire \reg_module/_09740_ ;
 wire \reg_module/_09741_ ;
 wire \reg_module/_09742_ ;
 wire \reg_module/_09743_ ;
 wire \reg_module/_09744_ ;
 wire \reg_module/_09745_ ;
 wire \reg_module/_09746_ ;
 wire \reg_module/_09747_ ;
 wire \reg_module/_09748_ ;
 wire \reg_module/_09749_ ;
 wire \reg_module/_09750_ ;
 wire \reg_module/_09751_ ;
 wire \reg_module/_09752_ ;
 wire \reg_module/_09753_ ;
 wire \reg_module/_09754_ ;
 wire \reg_module/_09755_ ;
 wire \reg_module/_09756_ ;
 wire \reg_module/_09757_ ;
 wire \reg_module/_09758_ ;
 wire \reg_module/_09759_ ;
 wire \reg_module/gprf[0] ;
 wire \reg_module/gprf[1000] ;
 wire \reg_module/gprf[1001] ;
 wire \reg_module/gprf[1002] ;
 wire \reg_module/gprf[1003] ;
 wire \reg_module/gprf[1004] ;
 wire \reg_module/gprf[1005] ;
 wire \reg_module/gprf[1006] ;
 wire \reg_module/gprf[1007] ;
 wire \reg_module/gprf[1008] ;
 wire \reg_module/gprf[1009] ;
 wire \reg_module/gprf[100] ;
 wire \reg_module/gprf[1010] ;
 wire \reg_module/gprf[1011] ;
 wire \reg_module/gprf[1012] ;
 wire \reg_module/gprf[1013] ;
 wire \reg_module/gprf[1014] ;
 wire \reg_module/gprf[1015] ;
 wire \reg_module/gprf[1016] ;
 wire \reg_module/gprf[1017] ;
 wire \reg_module/gprf[1018] ;
 wire \reg_module/gprf[1019] ;
 wire \reg_module/gprf[101] ;
 wire \reg_module/gprf[1020] ;
 wire \reg_module/gprf[1021] ;
 wire \reg_module/gprf[1022] ;
 wire \reg_module/gprf[1023] ;
 wire \reg_module/gprf[102] ;
 wire \reg_module/gprf[103] ;
 wire \reg_module/gprf[104] ;
 wire \reg_module/gprf[105] ;
 wire \reg_module/gprf[106] ;
 wire \reg_module/gprf[107] ;
 wire \reg_module/gprf[108] ;
 wire \reg_module/gprf[109] ;
 wire \reg_module/gprf[10] ;
 wire \reg_module/gprf[110] ;
 wire \reg_module/gprf[111] ;
 wire \reg_module/gprf[112] ;
 wire \reg_module/gprf[113] ;
 wire \reg_module/gprf[114] ;
 wire \reg_module/gprf[115] ;
 wire \reg_module/gprf[116] ;
 wire \reg_module/gprf[117] ;
 wire \reg_module/gprf[118] ;
 wire \reg_module/gprf[119] ;
 wire \reg_module/gprf[11] ;
 wire \reg_module/gprf[120] ;
 wire \reg_module/gprf[121] ;
 wire \reg_module/gprf[122] ;
 wire \reg_module/gprf[123] ;
 wire \reg_module/gprf[124] ;
 wire \reg_module/gprf[125] ;
 wire \reg_module/gprf[126] ;
 wire \reg_module/gprf[127] ;
 wire \reg_module/gprf[128] ;
 wire \reg_module/gprf[129] ;
 wire \reg_module/gprf[12] ;
 wire \reg_module/gprf[130] ;
 wire \reg_module/gprf[131] ;
 wire \reg_module/gprf[132] ;
 wire \reg_module/gprf[133] ;
 wire \reg_module/gprf[134] ;
 wire \reg_module/gprf[135] ;
 wire \reg_module/gprf[136] ;
 wire \reg_module/gprf[137] ;
 wire \reg_module/gprf[138] ;
 wire \reg_module/gprf[139] ;
 wire \reg_module/gprf[13] ;
 wire \reg_module/gprf[140] ;
 wire \reg_module/gprf[141] ;
 wire \reg_module/gprf[142] ;
 wire \reg_module/gprf[143] ;
 wire \reg_module/gprf[144] ;
 wire \reg_module/gprf[145] ;
 wire \reg_module/gprf[146] ;
 wire \reg_module/gprf[147] ;
 wire \reg_module/gprf[148] ;
 wire \reg_module/gprf[149] ;
 wire \reg_module/gprf[14] ;
 wire \reg_module/gprf[150] ;
 wire \reg_module/gprf[151] ;
 wire \reg_module/gprf[152] ;
 wire \reg_module/gprf[153] ;
 wire \reg_module/gprf[154] ;
 wire \reg_module/gprf[155] ;
 wire \reg_module/gprf[156] ;
 wire \reg_module/gprf[157] ;
 wire \reg_module/gprf[158] ;
 wire \reg_module/gprf[159] ;
 wire \reg_module/gprf[15] ;
 wire \reg_module/gprf[160] ;
 wire \reg_module/gprf[161] ;
 wire \reg_module/gprf[162] ;
 wire \reg_module/gprf[163] ;
 wire \reg_module/gprf[164] ;
 wire \reg_module/gprf[165] ;
 wire \reg_module/gprf[166] ;
 wire \reg_module/gprf[167] ;
 wire \reg_module/gprf[168] ;
 wire \reg_module/gprf[169] ;
 wire \reg_module/gprf[16] ;
 wire \reg_module/gprf[170] ;
 wire \reg_module/gprf[171] ;
 wire \reg_module/gprf[172] ;
 wire \reg_module/gprf[173] ;
 wire \reg_module/gprf[174] ;
 wire \reg_module/gprf[175] ;
 wire \reg_module/gprf[176] ;
 wire \reg_module/gprf[177] ;
 wire \reg_module/gprf[178] ;
 wire \reg_module/gprf[179] ;
 wire \reg_module/gprf[17] ;
 wire \reg_module/gprf[180] ;
 wire \reg_module/gprf[181] ;
 wire \reg_module/gprf[182] ;
 wire \reg_module/gprf[183] ;
 wire \reg_module/gprf[184] ;
 wire \reg_module/gprf[185] ;
 wire \reg_module/gprf[186] ;
 wire \reg_module/gprf[187] ;
 wire \reg_module/gprf[188] ;
 wire \reg_module/gprf[189] ;
 wire \reg_module/gprf[18] ;
 wire \reg_module/gprf[190] ;
 wire \reg_module/gprf[191] ;
 wire \reg_module/gprf[192] ;
 wire \reg_module/gprf[193] ;
 wire \reg_module/gprf[194] ;
 wire \reg_module/gprf[195] ;
 wire \reg_module/gprf[196] ;
 wire \reg_module/gprf[197] ;
 wire \reg_module/gprf[198] ;
 wire \reg_module/gprf[199] ;
 wire \reg_module/gprf[19] ;
 wire \reg_module/gprf[1] ;
 wire \reg_module/gprf[200] ;
 wire \reg_module/gprf[201] ;
 wire \reg_module/gprf[202] ;
 wire \reg_module/gprf[203] ;
 wire \reg_module/gprf[204] ;
 wire \reg_module/gprf[205] ;
 wire \reg_module/gprf[206] ;
 wire \reg_module/gprf[207] ;
 wire \reg_module/gprf[208] ;
 wire \reg_module/gprf[209] ;
 wire \reg_module/gprf[20] ;
 wire \reg_module/gprf[210] ;
 wire \reg_module/gprf[211] ;
 wire \reg_module/gprf[212] ;
 wire \reg_module/gprf[213] ;
 wire \reg_module/gprf[214] ;
 wire \reg_module/gprf[215] ;
 wire \reg_module/gprf[216] ;
 wire \reg_module/gprf[217] ;
 wire \reg_module/gprf[218] ;
 wire \reg_module/gprf[219] ;
 wire \reg_module/gprf[21] ;
 wire \reg_module/gprf[220] ;
 wire \reg_module/gprf[221] ;
 wire \reg_module/gprf[222] ;
 wire \reg_module/gprf[223] ;
 wire \reg_module/gprf[224] ;
 wire \reg_module/gprf[225] ;
 wire \reg_module/gprf[226] ;
 wire \reg_module/gprf[227] ;
 wire \reg_module/gprf[228] ;
 wire \reg_module/gprf[229] ;
 wire \reg_module/gprf[22] ;
 wire \reg_module/gprf[230] ;
 wire \reg_module/gprf[231] ;
 wire \reg_module/gprf[232] ;
 wire \reg_module/gprf[233] ;
 wire \reg_module/gprf[234] ;
 wire \reg_module/gprf[235] ;
 wire \reg_module/gprf[236] ;
 wire \reg_module/gprf[237] ;
 wire \reg_module/gprf[238] ;
 wire \reg_module/gprf[239] ;
 wire \reg_module/gprf[23] ;
 wire \reg_module/gprf[240] ;
 wire \reg_module/gprf[241] ;
 wire \reg_module/gprf[242] ;
 wire \reg_module/gprf[243] ;
 wire \reg_module/gprf[244] ;
 wire \reg_module/gprf[245] ;
 wire \reg_module/gprf[246] ;
 wire \reg_module/gprf[247] ;
 wire \reg_module/gprf[248] ;
 wire \reg_module/gprf[249] ;
 wire \reg_module/gprf[24] ;
 wire \reg_module/gprf[250] ;
 wire \reg_module/gprf[251] ;
 wire \reg_module/gprf[252] ;
 wire \reg_module/gprf[253] ;
 wire \reg_module/gprf[254] ;
 wire \reg_module/gprf[255] ;
 wire \reg_module/gprf[256] ;
 wire \reg_module/gprf[257] ;
 wire \reg_module/gprf[258] ;
 wire \reg_module/gprf[259] ;
 wire \reg_module/gprf[25] ;
 wire \reg_module/gprf[260] ;
 wire \reg_module/gprf[261] ;
 wire \reg_module/gprf[262] ;
 wire \reg_module/gprf[263] ;
 wire \reg_module/gprf[264] ;
 wire \reg_module/gprf[265] ;
 wire \reg_module/gprf[266] ;
 wire \reg_module/gprf[267] ;
 wire \reg_module/gprf[268] ;
 wire \reg_module/gprf[269] ;
 wire \reg_module/gprf[26] ;
 wire \reg_module/gprf[270] ;
 wire \reg_module/gprf[271] ;
 wire \reg_module/gprf[272] ;
 wire \reg_module/gprf[273] ;
 wire \reg_module/gprf[274] ;
 wire \reg_module/gprf[275] ;
 wire \reg_module/gprf[276] ;
 wire \reg_module/gprf[277] ;
 wire \reg_module/gprf[278] ;
 wire \reg_module/gprf[279] ;
 wire \reg_module/gprf[27] ;
 wire \reg_module/gprf[280] ;
 wire \reg_module/gprf[281] ;
 wire \reg_module/gprf[282] ;
 wire \reg_module/gprf[283] ;
 wire \reg_module/gprf[284] ;
 wire \reg_module/gprf[285] ;
 wire \reg_module/gprf[286] ;
 wire \reg_module/gprf[287] ;
 wire \reg_module/gprf[288] ;
 wire \reg_module/gprf[289] ;
 wire \reg_module/gprf[28] ;
 wire \reg_module/gprf[290] ;
 wire \reg_module/gprf[291] ;
 wire \reg_module/gprf[292] ;
 wire \reg_module/gprf[293] ;
 wire \reg_module/gprf[294] ;
 wire \reg_module/gprf[295] ;
 wire \reg_module/gprf[296] ;
 wire \reg_module/gprf[297] ;
 wire \reg_module/gprf[298] ;
 wire \reg_module/gprf[299] ;
 wire \reg_module/gprf[29] ;
 wire \reg_module/gprf[2] ;
 wire \reg_module/gprf[300] ;
 wire \reg_module/gprf[301] ;
 wire \reg_module/gprf[302] ;
 wire \reg_module/gprf[303] ;
 wire \reg_module/gprf[304] ;
 wire \reg_module/gprf[305] ;
 wire \reg_module/gprf[306] ;
 wire \reg_module/gprf[307] ;
 wire \reg_module/gprf[308] ;
 wire \reg_module/gprf[309] ;
 wire \reg_module/gprf[30] ;
 wire \reg_module/gprf[310] ;
 wire \reg_module/gprf[311] ;
 wire \reg_module/gprf[312] ;
 wire \reg_module/gprf[313] ;
 wire \reg_module/gprf[314] ;
 wire \reg_module/gprf[315] ;
 wire \reg_module/gprf[316] ;
 wire \reg_module/gprf[317] ;
 wire \reg_module/gprf[318] ;
 wire \reg_module/gprf[319] ;
 wire \reg_module/gprf[31] ;
 wire \reg_module/gprf[320] ;
 wire \reg_module/gprf[321] ;
 wire \reg_module/gprf[322] ;
 wire \reg_module/gprf[323] ;
 wire \reg_module/gprf[324] ;
 wire \reg_module/gprf[325] ;
 wire \reg_module/gprf[326] ;
 wire \reg_module/gprf[327] ;
 wire \reg_module/gprf[328] ;
 wire \reg_module/gprf[329] ;
 wire \reg_module/gprf[32] ;
 wire \reg_module/gprf[330] ;
 wire \reg_module/gprf[331] ;
 wire \reg_module/gprf[332] ;
 wire \reg_module/gprf[333] ;
 wire \reg_module/gprf[334] ;
 wire \reg_module/gprf[335] ;
 wire \reg_module/gprf[336] ;
 wire \reg_module/gprf[337] ;
 wire \reg_module/gprf[338] ;
 wire \reg_module/gprf[339] ;
 wire \reg_module/gprf[33] ;
 wire \reg_module/gprf[340] ;
 wire \reg_module/gprf[341] ;
 wire \reg_module/gprf[342] ;
 wire \reg_module/gprf[343] ;
 wire \reg_module/gprf[344] ;
 wire \reg_module/gprf[345] ;
 wire \reg_module/gprf[346] ;
 wire \reg_module/gprf[347] ;
 wire \reg_module/gprf[348] ;
 wire \reg_module/gprf[349] ;
 wire \reg_module/gprf[34] ;
 wire \reg_module/gprf[350] ;
 wire \reg_module/gprf[351] ;
 wire \reg_module/gprf[352] ;
 wire \reg_module/gprf[353] ;
 wire \reg_module/gprf[354] ;
 wire \reg_module/gprf[355] ;
 wire \reg_module/gprf[356] ;
 wire \reg_module/gprf[357] ;
 wire \reg_module/gprf[358] ;
 wire \reg_module/gprf[359] ;
 wire \reg_module/gprf[35] ;
 wire \reg_module/gprf[360] ;
 wire \reg_module/gprf[361] ;
 wire \reg_module/gprf[362] ;
 wire \reg_module/gprf[363] ;
 wire \reg_module/gprf[364] ;
 wire \reg_module/gprf[365] ;
 wire \reg_module/gprf[366] ;
 wire \reg_module/gprf[367] ;
 wire \reg_module/gprf[368] ;
 wire \reg_module/gprf[369] ;
 wire \reg_module/gprf[36] ;
 wire \reg_module/gprf[370] ;
 wire \reg_module/gprf[371] ;
 wire \reg_module/gprf[372] ;
 wire \reg_module/gprf[373] ;
 wire \reg_module/gprf[374] ;
 wire \reg_module/gprf[375] ;
 wire \reg_module/gprf[376] ;
 wire \reg_module/gprf[377] ;
 wire \reg_module/gprf[378] ;
 wire \reg_module/gprf[379] ;
 wire \reg_module/gprf[37] ;
 wire \reg_module/gprf[380] ;
 wire \reg_module/gprf[381] ;
 wire \reg_module/gprf[382] ;
 wire \reg_module/gprf[383] ;
 wire \reg_module/gprf[384] ;
 wire \reg_module/gprf[385] ;
 wire \reg_module/gprf[386] ;
 wire \reg_module/gprf[387] ;
 wire \reg_module/gprf[388] ;
 wire \reg_module/gprf[389] ;
 wire \reg_module/gprf[38] ;
 wire \reg_module/gprf[390] ;
 wire \reg_module/gprf[391] ;
 wire \reg_module/gprf[392] ;
 wire \reg_module/gprf[393] ;
 wire \reg_module/gprf[394] ;
 wire \reg_module/gprf[395] ;
 wire \reg_module/gprf[396] ;
 wire \reg_module/gprf[397] ;
 wire \reg_module/gprf[398] ;
 wire \reg_module/gprf[399] ;
 wire \reg_module/gprf[39] ;
 wire \reg_module/gprf[3] ;
 wire \reg_module/gprf[400] ;
 wire \reg_module/gprf[401] ;
 wire \reg_module/gprf[402] ;
 wire \reg_module/gprf[403] ;
 wire \reg_module/gprf[404] ;
 wire \reg_module/gprf[405] ;
 wire \reg_module/gprf[406] ;
 wire \reg_module/gprf[407] ;
 wire \reg_module/gprf[408] ;
 wire \reg_module/gprf[409] ;
 wire \reg_module/gprf[40] ;
 wire \reg_module/gprf[410] ;
 wire \reg_module/gprf[411] ;
 wire \reg_module/gprf[412] ;
 wire \reg_module/gprf[413] ;
 wire \reg_module/gprf[414] ;
 wire \reg_module/gprf[415] ;
 wire \reg_module/gprf[416] ;
 wire \reg_module/gprf[417] ;
 wire \reg_module/gprf[418] ;
 wire \reg_module/gprf[419] ;
 wire \reg_module/gprf[41] ;
 wire \reg_module/gprf[420] ;
 wire \reg_module/gprf[421] ;
 wire \reg_module/gprf[422] ;
 wire \reg_module/gprf[423] ;
 wire \reg_module/gprf[424] ;
 wire \reg_module/gprf[425] ;
 wire \reg_module/gprf[426] ;
 wire \reg_module/gprf[427] ;
 wire \reg_module/gprf[428] ;
 wire \reg_module/gprf[429] ;
 wire \reg_module/gprf[42] ;
 wire \reg_module/gprf[430] ;
 wire \reg_module/gprf[431] ;
 wire \reg_module/gprf[432] ;
 wire \reg_module/gprf[433] ;
 wire \reg_module/gprf[434] ;
 wire \reg_module/gprf[435] ;
 wire \reg_module/gprf[436] ;
 wire \reg_module/gprf[437] ;
 wire \reg_module/gprf[438] ;
 wire \reg_module/gprf[439] ;
 wire \reg_module/gprf[43] ;
 wire \reg_module/gprf[440] ;
 wire \reg_module/gprf[441] ;
 wire \reg_module/gprf[442] ;
 wire \reg_module/gprf[443] ;
 wire \reg_module/gprf[444] ;
 wire \reg_module/gprf[445] ;
 wire \reg_module/gprf[446] ;
 wire \reg_module/gprf[447] ;
 wire \reg_module/gprf[448] ;
 wire \reg_module/gprf[449] ;
 wire \reg_module/gprf[44] ;
 wire \reg_module/gprf[450] ;
 wire \reg_module/gprf[451] ;
 wire \reg_module/gprf[452] ;
 wire \reg_module/gprf[453] ;
 wire \reg_module/gprf[454] ;
 wire \reg_module/gprf[455] ;
 wire \reg_module/gprf[456] ;
 wire \reg_module/gprf[457] ;
 wire \reg_module/gprf[458] ;
 wire \reg_module/gprf[459] ;
 wire \reg_module/gprf[45] ;
 wire \reg_module/gprf[460] ;
 wire \reg_module/gprf[461] ;
 wire \reg_module/gprf[462] ;
 wire \reg_module/gprf[463] ;
 wire \reg_module/gprf[464] ;
 wire \reg_module/gprf[465] ;
 wire \reg_module/gprf[466] ;
 wire \reg_module/gprf[467] ;
 wire \reg_module/gprf[468] ;
 wire \reg_module/gprf[469] ;
 wire \reg_module/gprf[46] ;
 wire \reg_module/gprf[470] ;
 wire \reg_module/gprf[471] ;
 wire \reg_module/gprf[472] ;
 wire \reg_module/gprf[473] ;
 wire \reg_module/gprf[474] ;
 wire \reg_module/gprf[475] ;
 wire \reg_module/gprf[476] ;
 wire \reg_module/gprf[477] ;
 wire \reg_module/gprf[478] ;
 wire \reg_module/gprf[479] ;
 wire \reg_module/gprf[47] ;
 wire \reg_module/gprf[480] ;
 wire \reg_module/gprf[481] ;
 wire \reg_module/gprf[482] ;
 wire \reg_module/gprf[483] ;
 wire \reg_module/gprf[484] ;
 wire \reg_module/gprf[485] ;
 wire \reg_module/gprf[486] ;
 wire \reg_module/gprf[487] ;
 wire \reg_module/gprf[488] ;
 wire \reg_module/gprf[489] ;
 wire \reg_module/gprf[48] ;
 wire \reg_module/gprf[490] ;
 wire \reg_module/gprf[491] ;
 wire \reg_module/gprf[492] ;
 wire \reg_module/gprf[493] ;
 wire \reg_module/gprf[494] ;
 wire \reg_module/gprf[495] ;
 wire \reg_module/gprf[496] ;
 wire \reg_module/gprf[497] ;
 wire \reg_module/gprf[498] ;
 wire \reg_module/gprf[499] ;
 wire \reg_module/gprf[49] ;
 wire \reg_module/gprf[4] ;
 wire \reg_module/gprf[500] ;
 wire \reg_module/gprf[501] ;
 wire \reg_module/gprf[502] ;
 wire \reg_module/gprf[503] ;
 wire \reg_module/gprf[504] ;
 wire \reg_module/gprf[505] ;
 wire \reg_module/gprf[506] ;
 wire \reg_module/gprf[507] ;
 wire \reg_module/gprf[508] ;
 wire \reg_module/gprf[509] ;
 wire \reg_module/gprf[50] ;
 wire \reg_module/gprf[510] ;
 wire \reg_module/gprf[511] ;
 wire \reg_module/gprf[512] ;
 wire \reg_module/gprf[513] ;
 wire \reg_module/gprf[514] ;
 wire \reg_module/gprf[515] ;
 wire \reg_module/gprf[516] ;
 wire \reg_module/gprf[517] ;
 wire \reg_module/gprf[518] ;
 wire \reg_module/gprf[519] ;
 wire \reg_module/gprf[51] ;
 wire \reg_module/gprf[520] ;
 wire \reg_module/gprf[521] ;
 wire \reg_module/gprf[522] ;
 wire \reg_module/gprf[523] ;
 wire \reg_module/gprf[524] ;
 wire \reg_module/gprf[525] ;
 wire \reg_module/gprf[526] ;
 wire \reg_module/gprf[527] ;
 wire \reg_module/gprf[528] ;
 wire \reg_module/gprf[529] ;
 wire \reg_module/gprf[52] ;
 wire \reg_module/gprf[530] ;
 wire \reg_module/gprf[531] ;
 wire \reg_module/gprf[532] ;
 wire \reg_module/gprf[533] ;
 wire \reg_module/gprf[534] ;
 wire \reg_module/gprf[535] ;
 wire \reg_module/gprf[536] ;
 wire \reg_module/gprf[537] ;
 wire \reg_module/gprf[538] ;
 wire \reg_module/gprf[539] ;
 wire \reg_module/gprf[53] ;
 wire \reg_module/gprf[540] ;
 wire \reg_module/gprf[541] ;
 wire \reg_module/gprf[542] ;
 wire \reg_module/gprf[543] ;
 wire \reg_module/gprf[544] ;
 wire \reg_module/gprf[545] ;
 wire \reg_module/gprf[546] ;
 wire \reg_module/gprf[547] ;
 wire \reg_module/gprf[548] ;
 wire \reg_module/gprf[549] ;
 wire \reg_module/gprf[54] ;
 wire \reg_module/gprf[550] ;
 wire \reg_module/gprf[551] ;
 wire \reg_module/gprf[552] ;
 wire \reg_module/gprf[553] ;
 wire \reg_module/gprf[554] ;
 wire \reg_module/gprf[555] ;
 wire \reg_module/gprf[556] ;
 wire \reg_module/gprf[557] ;
 wire \reg_module/gprf[558] ;
 wire \reg_module/gprf[559] ;
 wire \reg_module/gprf[55] ;
 wire \reg_module/gprf[560] ;
 wire \reg_module/gprf[561] ;
 wire \reg_module/gprf[562] ;
 wire \reg_module/gprf[563] ;
 wire \reg_module/gprf[564] ;
 wire \reg_module/gprf[565] ;
 wire \reg_module/gprf[566] ;
 wire \reg_module/gprf[567] ;
 wire \reg_module/gprf[568] ;
 wire \reg_module/gprf[569] ;
 wire \reg_module/gprf[56] ;
 wire \reg_module/gprf[570] ;
 wire \reg_module/gprf[571] ;
 wire \reg_module/gprf[572] ;
 wire \reg_module/gprf[573] ;
 wire \reg_module/gprf[574] ;
 wire \reg_module/gprf[575] ;
 wire \reg_module/gprf[576] ;
 wire \reg_module/gprf[577] ;
 wire \reg_module/gprf[578] ;
 wire \reg_module/gprf[579] ;
 wire \reg_module/gprf[57] ;
 wire \reg_module/gprf[580] ;
 wire \reg_module/gprf[581] ;
 wire \reg_module/gprf[582] ;
 wire \reg_module/gprf[583] ;
 wire \reg_module/gprf[584] ;
 wire \reg_module/gprf[585] ;
 wire \reg_module/gprf[586] ;
 wire \reg_module/gprf[587] ;
 wire \reg_module/gprf[588] ;
 wire \reg_module/gprf[589] ;
 wire \reg_module/gprf[58] ;
 wire \reg_module/gprf[590] ;
 wire \reg_module/gprf[591] ;
 wire \reg_module/gprf[592] ;
 wire \reg_module/gprf[593] ;
 wire \reg_module/gprf[594] ;
 wire \reg_module/gprf[595] ;
 wire \reg_module/gprf[596] ;
 wire \reg_module/gprf[597] ;
 wire \reg_module/gprf[598] ;
 wire \reg_module/gprf[599] ;
 wire \reg_module/gprf[59] ;
 wire \reg_module/gprf[5] ;
 wire \reg_module/gprf[600] ;
 wire \reg_module/gprf[601] ;
 wire \reg_module/gprf[602] ;
 wire \reg_module/gprf[603] ;
 wire \reg_module/gprf[604] ;
 wire \reg_module/gprf[605] ;
 wire \reg_module/gprf[606] ;
 wire \reg_module/gprf[607] ;
 wire \reg_module/gprf[608] ;
 wire \reg_module/gprf[609] ;
 wire \reg_module/gprf[60] ;
 wire \reg_module/gprf[610] ;
 wire \reg_module/gprf[611] ;
 wire \reg_module/gprf[612] ;
 wire \reg_module/gprf[613] ;
 wire \reg_module/gprf[614] ;
 wire \reg_module/gprf[615] ;
 wire \reg_module/gprf[616] ;
 wire \reg_module/gprf[617] ;
 wire \reg_module/gprf[618] ;
 wire \reg_module/gprf[619] ;
 wire \reg_module/gprf[61] ;
 wire \reg_module/gprf[620] ;
 wire \reg_module/gprf[621] ;
 wire \reg_module/gprf[622] ;
 wire \reg_module/gprf[623] ;
 wire \reg_module/gprf[624] ;
 wire \reg_module/gprf[625] ;
 wire \reg_module/gprf[626] ;
 wire \reg_module/gprf[627] ;
 wire \reg_module/gprf[628] ;
 wire \reg_module/gprf[629] ;
 wire \reg_module/gprf[62] ;
 wire \reg_module/gprf[630] ;
 wire \reg_module/gprf[631] ;
 wire \reg_module/gprf[632] ;
 wire \reg_module/gprf[633] ;
 wire \reg_module/gprf[634] ;
 wire \reg_module/gprf[635] ;
 wire \reg_module/gprf[636] ;
 wire \reg_module/gprf[637] ;
 wire \reg_module/gprf[638] ;
 wire \reg_module/gprf[639] ;
 wire \reg_module/gprf[63] ;
 wire \reg_module/gprf[640] ;
 wire \reg_module/gprf[641] ;
 wire \reg_module/gprf[642] ;
 wire \reg_module/gprf[643] ;
 wire \reg_module/gprf[644] ;
 wire \reg_module/gprf[645] ;
 wire \reg_module/gprf[646] ;
 wire \reg_module/gprf[647] ;
 wire \reg_module/gprf[648] ;
 wire \reg_module/gprf[649] ;
 wire \reg_module/gprf[64] ;
 wire \reg_module/gprf[650] ;
 wire \reg_module/gprf[651] ;
 wire \reg_module/gprf[652] ;
 wire \reg_module/gprf[653] ;
 wire \reg_module/gprf[654] ;
 wire \reg_module/gprf[655] ;
 wire \reg_module/gprf[656] ;
 wire \reg_module/gprf[657] ;
 wire \reg_module/gprf[658] ;
 wire \reg_module/gprf[659] ;
 wire \reg_module/gprf[65] ;
 wire \reg_module/gprf[660] ;
 wire \reg_module/gprf[661] ;
 wire \reg_module/gprf[662] ;
 wire \reg_module/gprf[663] ;
 wire \reg_module/gprf[664] ;
 wire \reg_module/gprf[665] ;
 wire \reg_module/gprf[666] ;
 wire \reg_module/gprf[667] ;
 wire \reg_module/gprf[668] ;
 wire \reg_module/gprf[669] ;
 wire \reg_module/gprf[66] ;
 wire \reg_module/gprf[670] ;
 wire \reg_module/gprf[671] ;
 wire \reg_module/gprf[672] ;
 wire \reg_module/gprf[673] ;
 wire \reg_module/gprf[674] ;
 wire \reg_module/gprf[675] ;
 wire \reg_module/gprf[676] ;
 wire \reg_module/gprf[677] ;
 wire \reg_module/gprf[678] ;
 wire \reg_module/gprf[679] ;
 wire \reg_module/gprf[67] ;
 wire \reg_module/gprf[680] ;
 wire \reg_module/gprf[681] ;
 wire \reg_module/gprf[682] ;
 wire \reg_module/gprf[683] ;
 wire \reg_module/gprf[684] ;
 wire \reg_module/gprf[685] ;
 wire \reg_module/gprf[686] ;
 wire \reg_module/gprf[687] ;
 wire \reg_module/gprf[688] ;
 wire \reg_module/gprf[689] ;
 wire \reg_module/gprf[68] ;
 wire \reg_module/gprf[690] ;
 wire \reg_module/gprf[691] ;
 wire \reg_module/gprf[692] ;
 wire \reg_module/gprf[693] ;
 wire \reg_module/gprf[694] ;
 wire \reg_module/gprf[695] ;
 wire \reg_module/gprf[696] ;
 wire \reg_module/gprf[697] ;
 wire \reg_module/gprf[698] ;
 wire \reg_module/gprf[699] ;
 wire \reg_module/gprf[69] ;
 wire \reg_module/gprf[6] ;
 wire \reg_module/gprf[700] ;
 wire \reg_module/gprf[701] ;
 wire \reg_module/gprf[702] ;
 wire \reg_module/gprf[703] ;
 wire \reg_module/gprf[704] ;
 wire \reg_module/gprf[705] ;
 wire \reg_module/gprf[706] ;
 wire \reg_module/gprf[707] ;
 wire \reg_module/gprf[708] ;
 wire \reg_module/gprf[709] ;
 wire \reg_module/gprf[70] ;
 wire \reg_module/gprf[710] ;
 wire \reg_module/gprf[711] ;
 wire \reg_module/gprf[712] ;
 wire \reg_module/gprf[713] ;
 wire \reg_module/gprf[714] ;
 wire \reg_module/gprf[715] ;
 wire \reg_module/gprf[716] ;
 wire \reg_module/gprf[717] ;
 wire \reg_module/gprf[718] ;
 wire \reg_module/gprf[719] ;
 wire \reg_module/gprf[71] ;
 wire \reg_module/gprf[720] ;
 wire \reg_module/gprf[721] ;
 wire \reg_module/gprf[722] ;
 wire \reg_module/gprf[723] ;
 wire \reg_module/gprf[724] ;
 wire \reg_module/gprf[725] ;
 wire \reg_module/gprf[726] ;
 wire \reg_module/gprf[727] ;
 wire \reg_module/gprf[728] ;
 wire \reg_module/gprf[729] ;
 wire \reg_module/gprf[72] ;
 wire \reg_module/gprf[730] ;
 wire \reg_module/gprf[731] ;
 wire \reg_module/gprf[732] ;
 wire \reg_module/gprf[733] ;
 wire \reg_module/gprf[734] ;
 wire \reg_module/gprf[735] ;
 wire \reg_module/gprf[736] ;
 wire \reg_module/gprf[737] ;
 wire \reg_module/gprf[738] ;
 wire \reg_module/gprf[739] ;
 wire \reg_module/gprf[73] ;
 wire \reg_module/gprf[740] ;
 wire \reg_module/gprf[741] ;
 wire \reg_module/gprf[742] ;
 wire \reg_module/gprf[743] ;
 wire \reg_module/gprf[744] ;
 wire \reg_module/gprf[745] ;
 wire \reg_module/gprf[746] ;
 wire \reg_module/gprf[747] ;
 wire \reg_module/gprf[748] ;
 wire \reg_module/gprf[749] ;
 wire \reg_module/gprf[74] ;
 wire \reg_module/gprf[750] ;
 wire \reg_module/gprf[751] ;
 wire \reg_module/gprf[752] ;
 wire \reg_module/gprf[753] ;
 wire \reg_module/gprf[754] ;
 wire \reg_module/gprf[755] ;
 wire \reg_module/gprf[756] ;
 wire \reg_module/gprf[757] ;
 wire \reg_module/gprf[758] ;
 wire \reg_module/gprf[759] ;
 wire \reg_module/gprf[75] ;
 wire \reg_module/gprf[760] ;
 wire \reg_module/gprf[761] ;
 wire \reg_module/gprf[762] ;
 wire \reg_module/gprf[763] ;
 wire \reg_module/gprf[764] ;
 wire \reg_module/gprf[765] ;
 wire \reg_module/gprf[766] ;
 wire \reg_module/gprf[767] ;
 wire \reg_module/gprf[768] ;
 wire \reg_module/gprf[769] ;
 wire \reg_module/gprf[76] ;
 wire \reg_module/gprf[770] ;
 wire \reg_module/gprf[771] ;
 wire \reg_module/gprf[772] ;
 wire \reg_module/gprf[773] ;
 wire \reg_module/gprf[774] ;
 wire \reg_module/gprf[775] ;
 wire \reg_module/gprf[776] ;
 wire \reg_module/gprf[777] ;
 wire \reg_module/gprf[778] ;
 wire \reg_module/gprf[779] ;
 wire \reg_module/gprf[77] ;
 wire \reg_module/gprf[780] ;
 wire \reg_module/gprf[781] ;
 wire \reg_module/gprf[782] ;
 wire \reg_module/gprf[783] ;
 wire \reg_module/gprf[784] ;
 wire \reg_module/gprf[785] ;
 wire \reg_module/gprf[786] ;
 wire \reg_module/gprf[787] ;
 wire \reg_module/gprf[788] ;
 wire \reg_module/gprf[789] ;
 wire \reg_module/gprf[78] ;
 wire \reg_module/gprf[790] ;
 wire \reg_module/gprf[791] ;
 wire \reg_module/gprf[792] ;
 wire \reg_module/gprf[793] ;
 wire \reg_module/gprf[794] ;
 wire \reg_module/gprf[795] ;
 wire \reg_module/gprf[796] ;
 wire \reg_module/gprf[797] ;
 wire \reg_module/gprf[798] ;
 wire \reg_module/gprf[799] ;
 wire \reg_module/gprf[79] ;
 wire \reg_module/gprf[7] ;
 wire \reg_module/gprf[800] ;
 wire \reg_module/gprf[801] ;
 wire \reg_module/gprf[802] ;
 wire \reg_module/gprf[803] ;
 wire \reg_module/gprf[804] ;
 wire \reg_module/gprf[805] ;
 wire \reg_module/gprf[806] ;
 wire \reg_module/gprf[807] ;
 wire \reg_module/gprf[808] ;
 wire \reg_module/gprf[809] ;
 wire \reg_module/gprf[80] ;
 wire \reg_module/gprf[810] ;
 wire \reg_module/gprf[811] ;
 wire \reg_module/gprf[812] ;
 wire \reg_module/gprf[813] ;
 wire \reg_module/gprf[814] ;
 wire \reg_module/gprf[815] ;
 wire \reg_module/gprf[816] ;
 wire \reg_module/gprf[817] ;
 wire \reg_module/gprf[818] ;
 wire \reg_module/gprf[819] ;
 wire \reg_module/gprf[81] ;
 wire \reg_module/gprf[820] ;
 wire \reg_module/gprf[821] ;
 wire \reg_module/gprf[822] ;
 wire \reg_module/gprf[823] ;
 wire \reg_module/gprf[824] ;
 wire \reg_module/gprf[825] ;
 wire \reg_module/gprf[826] ;
 wire \reg_module/gprf[827] ;
 wire \reg_module/gprf[828] ;
 wire \reg_module/gprf[829] ;
 wire \reg_module/gprf[82] ;
 wire \reg_module/gprf[830] ;
 wire \reg_module/gprf[831] ;
 wire \reg_module/gprf[832] ;
 wire \reg_module/gprf[833] ;
 wire \reg_module/gprf[834] ;
 wire \reg_module/gprf[835] ;
 wire \reg_module/gprf[836] ;
 wire \reg_module/gprf[837] ;
 wire \reg_module/gprf[838] ;
 wire \reg_module/gprf[839] ;
 wire \reg_module/gprf[83] ;
 wire \reg_module/gprf[840] ;
 wire \reg_module/gprf[841] ;
 wire \reg_module/gprf[842] ;
 wire \reg_module/gprf[843] ;
 wire \reg_module/gprf[844] ;
 wire \reg_module/gprf[845] ;
 wire \reg_module/gprf[846] ;
 wire \reg_module/gprf[847] ;
 wire \reg_module/gprf[848] ;
 wire \reg_module/gprf[849] ;
 wire \reg_module/gprf[84] ;
 wire \reg_module/gprf[850] ;
 wire \reg_module/gprf[851] ;
 wire \reg_module/gprf[852] ;
 wire \reg_module/gprf[853] ;
 wire \reg_module/gprf[854] ;
 wire \reg_module/gprf[855] ;
 wire \reg_module/gprf[856] ;
 wire \reg_module/gprf[857] ;
 wire \reg_module/gprf[858] ;
 wire \reg_module/gprf[859] ;
 wire \reg_module/gprf[85] ;
 wire \reg_module/gprf[860] ;
 wire \reg_module/gprf[861] ;
 wire \reg_module/gprf[862] ;
 wire \reg_module/gprf[863] ;
 wire \reg_module/gprf[864] ;
 wire \reg_module/gprf[865] ;
 wire \reg_module/gprf[866] ;
 wire \reg_module/gprf[867] ;
 wire \reg_module/gprf[868] ;
 wire \reg_module/gprf[869] ;
 wire \reg_module/gprf[86] ;
 wire \reg_module/gprf[870] ;
 wire \reg_module/gprf[871] ;
 wire \reg_module/gprf[872] ;
 wire \reg_module/gprf[873] ;
 wire \reg_module/gprf[874] ;
 wire \reg_module/gprf[875] ;
 wire \reg_module/gprf[876] ;
 wire \reg_module/gprf[877] ;
 wire \reg_module/gprf[878] ;
 wire \reg_module/gprf[879] ;
 wire \reg_module/gprf[87] ;
 wire \reg_module/gprf[880] ;
 wire \reg_module/gprf[881] ;
 wire \reg_module/gprf[882] ;
 wire \reg_module/gprf[883] ;
 wire \reg_module/gprf[884] ;
 wire \reg_module/gprf[885] ;
 wire \reg_module/gprf[886] ;
 wire \reg_module/gprf[887] ;
 wire \reg_module/gprf[888] ;
 wire \reg_module/gprf[889] ;
 wire \reg_module/gprf[88] ;
 wire \reg_module/gprf[890] ;
 wire \reg_module/gprf[891] ;
 wire \reg_module/gprf[892] ;
 wire \reg_module/gprf[893] ;
 wire \reg_module/gprf[894] ;
 wire \reg_module/gprf[895] ;
 wire \reg_module/gprf[896] ;
 wire \reg_module/gprf[897] ;
 wire \reg_module/gprf[898] ;
 wire \reg_module/gprf[899] ;
 wire \reg_module/gprf[89] ;
 wire \reg_module/gprf[8] ;
 wire \reg_module/gprf[900] ;
 wire \reg_module/gprf[901] ;
 wire \reg_module/gprf[902] ;
 wire \reg_module/gprf[903] ;
 wire \reg_module/gprf[904] ;
 wire \reg_module/gprf[905] ;
 wire \reg_module/gprf[906] ;
 wire \reg_module/gprf[907] ;
 wire \reg_module/gprf[908] ;
 wire \reg_module/gprf[909] ;
 wire \reg_module/gprf[90] ;
 wire \reg_module/gprf[910] ;
 wire \reg_module/gprf[911] ;
 wire \reg_module/gprf[912] ;
 wire \reg_module/gprf[913] ;
 wire \reg_module/gprf[914] ;
 wire \reg_module/gprf[915] ;
 wire \reg_module/gprf[916] ;
 wire \reg_module/gprf[917] ;
 wire \reg_module/gprf[918] ;
 wire \reg_module/gprf[919] ;
 wire \reg_module/gprf[91] ;
 wire \reg_module/gprf[920] ;
 wire \reg_module/gprf[921] ;
 wire \reg_module/gprf[922] ;
 wire \reg_module/gprf[923] ;
 wire \reg_module/gprf[924] ;
 wire \reg_module/gprf[925] ;
 wire \reg_module/gprf[926] ;
 wire \reg_module/gprf[927] ;
 wire \reg_module/gprf[928] ;
 wire \reg_module/gprf[929] ;
 wire \reg_module/gprf[92] ;
 wire \reg_module/gprf[930] ;
 wire \reg_module/gprf[931] ;
 wire \reg_module/gprf[932] ;
 wire \reg_module/gprf[933] ;
 wire \reg_module/gprf[934] ;
 wire \reg_module/gprf[935] ;
 wire \reg_module/gprf[936] ;
 wire \reg_module/gprf[937] ;
 wire \reg_module/gprf[938] ;
 wire \reg_module/gprf[939] ;
 wire \reg_module/gprf[93] ;
 wire \reg_module/gprf[940] ;
 wire \reg_module/gprf[941] ;
 wire \reg_module/gprf[942] ;
 wire \reg_module/gprf[943] ;
 wire \reg_module/gprf[944] ;
 wire \reg_module/gprf[945] ;
 wire \reg_module/gprf[946] ;
 wire \reg_module/gprf[947] ;
 wire \reg_module/gprf[948] ;
 wire \reg_module/gprf[949] ;
 wire \reg_module/gprf[94] ;
 wire \reg_module/gprf[950] ;
 wire \reg_module/gprf[951] ;
 wire \reg_module/gprf[952] ;
 wire \reg_module/gprf[953] ;
 wire \reg_module/gprf[954] ;
 wire \reg_module/gprf[955] ;
 wire \reg_module/gprf[956] ;
 wire \reg_module/gprf[957] ;
 wire \reg_module/gprf[958] ;
 wire \reg_module/gprf[959] ;
 wire \reg_module/gprf[95] ;
 wire \reg_module/gprf[960] ;
 wire \reg_module/gprf[961] ;
 wire \reg_module/gprf[962] ;
 wire \reg_module/gprf[963] ;
 wire \reg_module/gprf[964] ;
 wire \reg_module/gprf[965] ;
 wire \reg_module/gprf[966] ;
 wire \reg_module/gprf[967] ;
 wire \reg_module/gprf[968] ;
 wire \reg_module/gprf[969] ;
 wire \reg_module/gprf[96] ;
 wire \reg_module/gprf[970] ;
 wire \reg_module/gprf[971] ;
 wire \reg_module/gprf[972] ;
 wire \reg_module/gprf[973] ;
 wire \reg_module/gprf[974] ;
 wire \reg_module/gprf[975] ;
 wire \reg_module/gprf[976] ;
 wire \reg_module/gprf[977] ;
 wire \reg_module/gprf[978] ;
 wire \reg_module/gprf[979] ;
 wire \reg_module/gprf[97] ;
 wire \reg_module/gprf[980] ;
 wire \reg_module/gprf[981] ;
 wire \reg_module/gprf[982] ;
 wire \reg_module/gprf[983] ;
 wire \reg_module/gprf[984] ;
 wire \reg_module/gprf[985] ;
 wire \reg_module/gprf[986] ;
 wire \reg_module/gprf[987] ;
 wire \reg_module/gprf[988] ;
 wire \reg_module/gprf[989] ;
 wire \reg_module/gprf[98] ;
 wire \reg_module/gprf[990] ;
 wire \reg_module/gprf[991] ;
 wire \reg_module/gprf[992] ;
 wire \reg_module/gprf[993] ;
 wire \reg_module/gprf[994] ;
 wire \reg_module/gprf[995] ;
 wire \reg_module/gprf[996] ;
 wire \reg_module/gprf[997] ;
 wire \reg_module/gprf[998] ;
 wire \reg_module/gprf[999] ;
 wire \reg_module/gprf[99] ;
 wire \reg_module/gprf[9] ;
 wire \reg_module/rRs1[0] ;
 wire \reg_module/rRs1[1] ;
 wire \reg_module/rRs1[2] ;
 wire \reg_module/rRs1[3] ;
 wire \reg_module/rRs1[4] ;
 wire \reg_module/rRs2[0] ;
 wire \reg_module/rRs2[1] ;
 wire \reg_module/rRs2[2] ;
 wire \reg_module/rRs2[3] ;
 wire \reg_module/rRs2[4] ;
 wire \rpc/_000_ ;
 wire \rpc/_001_ ;
 wire \rpc/_002_ ;
 wire \rpc/_003_ ;
 wire \rpc/_004_ ;
 wire \rpc/_005_ ;
 wire \rpc/_006_ ;
 wire \rpc/_007_ ;
 wire \rpc/_008_ ;
 wire \rpc/_009_ ;
 wire \rpc/_010_ ;
 wire \rpc/_011_ ;
 wire \rpc/_012_ ;
 wire \rpc/_013_ ;
 wire \rpc/_014_ ;
 wire \rpc/_015_ ;
 wire \rpc/_016_ ;
 wire \rpc/_017_ ;
 wire \rpc/_018_ ;
 wire \rpc/_019_ ;
 wire \rpc/_020_ ;
 wire \rpc/_021_ ;
 wire \rpc/_022_ ;
 wire \rpc/_023_ ;
 wire \rpc/_024_ ;
 wire \rpc/_025_ ;
 wire \rpc/_026_ ;
 wire \rpc/_027_ ;
 wire \rpc/_028_ ;
 wire \rpc/_029_ ;
 wire \rpc/_030_ ;
 wire \rpc/_031_ ;
 wire \rpc/_032_ ;
 wire \rpc/_033_ ;
 wire \rpc/_034_ ;
 wire \rpc/_035_ ;
 wire \rpc/_036_ ;
 wire \rpc/_037_ ;
 wire \rpc/_038_ ;
 wire \rpc/_039_ ;
 wire \rpc/_040_ ;
 wire \rpc/_041_ ;
 wire \rpc/_042_ ;
 wire \rpc/_043_ ;
 wire \rpc/_044_ ;
 wire \rpc/_045_ ;
 wire \rpc/_046_ ;
 wire \rpc/_047_ ;
 wire \rpc/_048_ ;
 wire \rpc/_049_ ;
 wire \rpc/_050_ ;
 wire \rpc/_051_ ;
 wire \rpc/_052_ ;
 wire \rpc/_053_ ;
 wire \rpc/_054_ ;
 wire \rpc/_055_ ;
 wire \rpc/_056_ ;
 wire \rpc/_057_ ;
 wire \rpc/_058_ ;
 wire \rpc/_059_ ;
 wire \rpc/_060_ ;
 wire \rpc/_061_ ;
 wire \rpc/_062_ ;
 wire \rpc/_063_ ;
 wire \rpc/_064_ ;
 wire \rpc/_065_ ;
 wire \rpc/_066_ ;
 wire \rpc/_067_ ;
 wire \rpc/_068_ ;
 wire \rpc/_069_ ;
 wire \rpc/_070_ ;
 wire \rpc/_071_ ;
 wire \rpc/_072_ ;
 wire \rpc/_073_ ;
 wire \rpc/_074_ ;
 wire \rpc/_075_ ;
 wire \rpc/_076_ ;
 wire \rpc/_077_ ;
 wire \rpc/_078_ ;
 wire \rpc/_079_ ;
 wire \rpc/_080_ ;
 wire \rpc/_081_ ;
 wire \rpc/_082_ ;
 wire \rpc/_083_ ;
 wire \rpc/_084_ ;
 wire \rpc/_085_ ;
 wire \rpc/_086_ ;
 wire \rpc/_087_ ;
 wire \rpc/_088_ ;
 wire \rpc/_089_ ;
 wire \rpc/_090_ ;
 wire \rpc/_091_ ;
 wire \rpc/_092_ ;
 wire \rpc/_093_ ;
 wire \rpc/_094_ ;
 wire \rpc/_095_ ;
 wire \rpc/_096_ ;
 wire \rpc/_097_ ;
 wire \rpc/_098_ ;
 wire \rpc/_099_ ;
 wire \rpc/_100_ ;
 wire \rpc/_101_ ;
 wire \rpc/_102_ ;
 wire \rpc/_103_ ;
 wire \rpc/_104_ ;
 wire \rpc/_105_ ;
 wire \rpc/_106_ ;
 wire \rpc/_107_ ;
 wire \rpc/_108_ ;
 wire \rpc/_109_ ;
 wire \rpc/_110_ ;
 wire \rpc/_111_ ;
 wire \rpc/_112_ ;
 wire \rpc/_113_ ;
 wire \rpc/_114_ ;
 wire \rpc/_115_ ;
 wire \rpc/_116_ ;
 wire \rpc/_117_ ;
 wire \rpc/_118_ ;
 wire \rpc/_119_ ;
 wire \rpc/_120_ ;
 wire \rpc/_121_ ;
 wire \rpc/_122_ ;
 wire \rpc/_123_ ;
 wire \rpc/_124_ ;
 wire \rpc/_125_ ;
 wire \rpc/_126_ ;
 wire \rpc/_127_ ;
 wire \rpc/_128_ ;
 wire \rpc/_129_ ;
 wire \rpc/_130_ ;
 wire \rpc/_131_ ;
 wire \rpc/_132_ ;
 wire \rpc/_133_ ;
 wire \rpc/_134_ ;
 wire \rpc/_135_ ;
 wire \rpc/_136_ ;
 wire \rpc/_137_ ;
 wire \rpc/_138_ ;
 wire \rpc/_139_ ;
 wire \rpc/_140_ ;
 wire \rpc/_141_ ;
 wire \rpc/_142_ ;
 wire \rpc/_143_ ;
 wire \rpc/_144_ ;
 wire \rpc/_145_ ;
 wire \rpc/_146_ ;
 wire \rpc/_147_ ;
 wire \rpc/_148_ ;
 wire \rpc/_149_ ;
 wire \rpc/_150_ ;
 wire \rpc/_151_ ;
 wire \rpc/_152_ ;
 wire \rpc/_153_ ;
 wire \rpc/_154_ ;
 wire \rpc/_155_ ;
 wire \rpc/_156_ ;
 wire \rpc/_157_ ;
 wire \rpc/_158_ ;
 wire \rpc/_159_ ;
 wire \rpc/_160_ ;
 wire \rpc/_161_ ;
 wire \rpc/_162_ ;
 wire \rpc/_163_ ;
 wire \rpc/_164_ ;
 wire \rpc/_165_ ;
 wire \rpc/_166_ ;
 wire \rpc/_167_ ;
 wire \rpc/_168_ ;
 wire \rpc/_169_ ;
 wire \rpc/_170_ ;
 wire \rpc/_171_ ;
 wire \rpc/_172_ ;
 wire \rpc/_173_ ;
 wire \rpc/_174_ ;
 wire \rpc/_175_ ;
 wire \rpc/_176_ ;
 wire \rpc/_177_ ;
 wire \rpc/_178_ ;
 wire \rpc/_179_ ;
 wire \rpc/_180_ ;
 wire \rpc/_181_ ;
 wire \rpc/_182_ ;
 wire \rpc/_183_ ;
 wire \rpc/_184_ ;
 wire \rpc/_185_ ;
 wire \rpc/_186_ ;
 wire \rpc/_187_ ;
 wire \rpc/_188_ ;
 wire \rpc/_189_ ;
 wire \rpc/_190_ ;
 wire \rpc/_191_ ;
 wire \rpc/_192_ ;
 wire \rpc/_193_ ;
 wire \rpc/_194_ ;
 wire \rpc/_195_ ;
 wire \rpc/_196_ ;
 wire \rpc/_197_ ;
 wire \rpc/_198_ ;
 wire \rpc/_199_ ;
 wire \rpc/_200_ ;
 wire \rpc/_201_ ;
 wire \rpc/_202_ ;
 wire \rpc/_203_ ;
 wire \rpc/_204_ ;
 wire \rpc/_205_ ;
 wire \rpc/_206_ ;
 wire \rpc/_207_ ;
 wire \rpc/_208_ ;
 wire \rpc/_209_ ;
 wire \rpc/_210_ ;
 wire \rpc/_211_ ;
 wire \rpc/_212_ ;
 wire \rpc/_213_ ;
 wire \rpc/_214_ ;
 wire \rpc/_215_ ;
 wire \rpc/_216_ ;
 wire \rpc/_217_ ;
 wire \rpc/_218_ ;
 wire \rpc/_219_ ;
 wire \rpc/_220_ ;
 wire \rpc/_221_ ;
 wire \rpc/_222_ ;
 wire \rpc/_223_ ;
 wire \rpc/_224_ ;
 wire \rpc/_225_ ;
 wire \rpc/_226_ ;
 wire \rpc/_227_ ;
 wire \rpc/_228_ ;
 wire \rpc/_229_ ;
 wire \rpc/_230_ ;
 wire \rpc/_231_ ;
 wire \rpc/_232_ ;
 wire \rpc/_233_ ;
 wire \rpc/_234_ ;
 wire \rpc/_235_ ;
 wire \rpc/_236_ ;
 wire \rpc/_237_ ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1077;
 wire net1079;
 wire net1081;
 wire net1083;
 wire net1085;
 wire net1087;
 wire net1089;
 wire net1091;
 wire net1093;
 wire net1095;
 wire net1097;
 wire net1099;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_leaf_98_clk;
 wire clknet_leaf_99_clk;
 wire clknet_leaf_100_clk;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_102_clk;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_113_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_133_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_138_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_leaf_145_clk;
 wire clknet_leaf_146_clk;
 wire clknet_leaf_147_clk;
 wire clknet_leaf_148_clk;
 wire clknet_leaf_149_clk;
 wire clknet_leaf_150_clk;
 wire clknet_leaf_151_clk;
 wire clknet_leaf_152_clk;
 wire clknet_leaf_153_clk;
 wire clknet_leaf_154_clk;
 wire clknet_leaf_155_clk;
 wire clknet_leaf_156_clk;
 wire clknet_leaf_157_clk;
 wire clknet_leaf_158_clk;
 wire clknet_leaf_159_clk;
 wire clknet_leaf_160_clk;
 wire clknet_leaf_161_clk;
 wire clknet_leaf_162_clk;
 wire clknet_leaf_163_clk;
 wire clknet_leaf_164_clk;
 wire clknet_leaf_165_clk;
 wire clknet_leaf_166_clk;
 wire clknet_leaf_167_clk;
 wire clknet_leaf_168_clk;
 wire clknet_leaf_169_clk;
 wire clknet_leaf_170_clk;
 wire clknet_leaf_171_clk;
 wire clknet_leaf_172_clk;
 wire clknet_leaf_173_clk;
 wire clknet_leaf_174_clk;
 wire clknet_leaf_175_clk;
 wire clknet_leaf_176_clk;
 wire clknet_leaf_177_clk;
 wire clknet_leaf_178_clk;
 wire clknet_leaf_179_clk;
 wire clknet_leaf_180_clk;
 wire clknet_leaf_181_clk;
 wire clknet_leaf_182_clk;
 wire clknet_leaf_183_clk;
 wire clknet_leaf_184_clk;
 wire clknet_leaf_185_clk;
 wire clknet_leaf_186_clk;
 wire clknet_leaf_187_clk;
 wire clknet_leaf_188_clk;
 wire clknet_leaf_189_clk;
 wire clknet_leaf_190_clk;
 wire clknet_leaf_191_clk;
 wire clknet_leaf_192_clk;
 wire clknet_leaf_193_clk;
 wire clknet_leaf_194_clk;
 wire clknet_leaf_195_clk;
 wire clknet_leaf_196_clk;
 wire clknet_leaf_197_clk;
 wire clknet_leaf_198_clk;
 wire clknet_leaf_199_clk;
 wire clknet_leaf_200_clk;
 wire clknet_leaf_201_clk;
 wire clknet_leaf_202_clk;
 wire clknet_leaf_203_clk;
 wire clknet_leaf_204_clk;
 wire clknet_leaf_205_clk;
 wire clknet_leaf_206_clk;
 wire clknet_leaf_207_clk;
 wire clknet_leaf_208_clk;
 wire clknet_leaf_209_clk;
 wire clknet_leaf_210_clk;
 wire clknet_leaf_211_clk;
 wire clknet_leaf_212_clk;
 wire clknet_leaf_213_clk;
 wire clknet_leaf_214_clk;
 wire clknet_leaf_215_clk;
 wire clknet_leaf_216_clk;
 wire clknet_leaf_217_clk;
 wire clknet_leaf_218_clk;
 wire clknet_leaf_219_clk;
 wire clknet_leaf_220_clk;
 wire clknet_leaf_221_clk;
 wire clknet_leaf_222_clk;
 wire clknet_leaf_223_clk;
 wire clknet_0_clk;
 wire clknet_2_0_0_clk;
 wire clknet_2_1_0_clk;
 wire clknet_2_2_0_clk;
 wire clknet_2_3_0_clk;
 wire clknet_4_0__leaf_clk;
 wire clknet_4_1__leaf_clk;
 wire clknet_4_2__leaf_clk;
 wire clknet_4_3__leaf_clk;
 wire clknet_4_4__leaf_clk;
 wire clknet_4_5__leaf_clk;
 wire clknet_4_6__leaf_clk;
 wire clknet_4_7__leaf_clk;
 wire clknet_4_8__leaf_clk;
 wire clknet_4_9__leaf_clk;
 wire clknet_4_10__leaf_clk;
 wire clknet_4_11__leaf_clk;
 wire clknet_4_12__leaf_clk;
 wire clknet_4_13__leaf_clk;
 wire clknet_4_14__leaf_clk;
 wire clknet_4_15__leaf_clk;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;

 sky130_fd_sc_hd__inv_2 _0963_ (.A(\funct3[0] ),
    .Y(_0592_));
 sky130_fd_sc_hd__nor2_1 _0964_ (.A(\funct3[1] ),
    .B(_0592_),
    .Y(wRamHalfEn));
 sky130_fd_sc_hd__inv_2 _0965_ (.A(\funct3[1] ),
    .Y(_0593_));
 sky130_fd_sc_hd__nor2_2 _0966_ (.A(\funct3[0] ),
    .B(_0593_),
    .Y(wRamWordEn));
 sky130_fd_sc_hd__inv_2 _0967_ (.A(\rReg_d[1] ),
    .Y(_0594_));
 sky130_fd_sc_hd__inv_2 _0968_ (.A(\rReg_d[0] ),
    .Y(_0595_));
 sky130_fd_sc_hd__nand2_1 _0969_ (.A(_0595_),
    .B(\reg_s1[0] ),
    .Y(_0596_));
 sky130_fd_sc_hd__inv_2 _0970_ (.A(\reg_s1[0] ),
    .Y(_0597_));
 sky130_fd_sc_hd__nand2_1 _0971_ (.A(_0597_),
    .B(\rReg_d[0] ),
    .Y(_0598_));
 sky130_fd_sc_hd__o211ai_1 _0972_ (.A1(\reg_s1[1] ),
    .A2(_0594_),
    .B1(_0596_),
    .C1(_0598_),
    .Y(_0599_));
 sky130_fd_sc_hd__nor2_1 _0973_ (.A(\rReg_d[0] ),
    .B(\rReg_d[1] ),
    .Y(_0600_));
 sky130_fd_sc_hd__nor2_1 _0974_ (.A(\rReg_d[2] ),
    .B(\rReg_d[4] ),
    .Y(_0601_));
 sky130_fd_sc_hd__inv_4 _0975_ (.A(\rReg_d[3] ),
    .Y(_0602_));
 sky130_fd_sc_hd__and3_1 _0976_ (.A(_0600_),
    .B(_0601_),
    .C(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__nor2_1 _0977_ (.A(_0599_),
    .B(_0603_),
    .Y(_0604_));
 sky130_fd_sc_hd__xnor2_1 _0978_ (.A(\reg_s1[4] ),
    .B(\rReg_d[4] ),
    .Y(_0605_));
 sky130_fd_sc_hd__a21boi_1 _0979_ (.A1(_0602_),
    .A2(\reg_s1[3] ),
    .B1_N(rRegWrEn),
    .Y(_0606_));
 sky130_fd_sc_hd__nand2_1 _0980_ (.A(_0605_),
    .B(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__inv_2 _0981_ (.A(\reg_s1[3] ),
    .Y(_0608_));
 sky130_fd_sc_hd__nand2_1 _0982_ (.A(_0608_),
    .B(\rReg_d[3] ),
    .Y(_0609_));
 sky130_fd_sc_hd__nand2_1 _0983_ (.A(_0594_),
    .B(\reg_s1[1] ),
    .Y(_0610_));
 sky130_fd_sc_hd__nand2_1 _0984_ (.A(_0609_),
    .B(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__inv_2 _0985_ (.A(_0611_),
    .Y(_0612_));
 sky130_fd_sc_hd__xnor2_1 _0986_ (.A(\reg_s1[2] ),
    .B(\rReg_d[2] ),
    .Y(_0613_));
 sky130_fd_sc_hd__nand2_1 _0987_ (.A(_0612_),
    .B(_0613_),
    .Y(_0614_));
 sky130_fd_sc_hd__nor2_1 _0988_ (.A(_0607_),
    .B(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__nand2_4 _0989_ (.A(_0604_),
    .B(_0615_),
    .Y(_0616_));
 sky130_fd_sc_hd__inv_2 _0990_ (.A(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__buf_4 _0991_ (.A(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__clkbuf_2 _0992_ (.A(_0618_),
    .X(_0619_));
 sky130_fd_sc_hd__clkbuf_2 _0993_ (.A(_0619_),
    .X(_0620_));
 sky130_fd_sc_hd__inv_2 _0994_ (.A(\reg_s2[1] ),
    .Y(_0621_));
 sky130_fd_sc_hd__xnor2_1 _0995_ (.A(\rReg_d[2] ),
    .B(\reg_s2[2] ),
    .Y(_0622_));
 sky130_fd_sc_hd__o221a_1 _0996_ (.A1(\rReg_d[1] ),
    .A2(_0621_),
    .B1(_0602_),
    .B2(\reg_s2[3] ),
    .C1(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__xnor2_1 _0997_ (.A(\rReg_d[4] ),
    .B(\reg_s2[4] ),
    .Y(_0624_));
 sky130_fd_sc_hd__nand2_1 _0998_ (.A(_0602_),
    .B(\reg_s2[3] ),
    .Y(_0625_));
 sky130_fd_sc_hd__and4_1 _0999_ (.A(_0623_),
    .B(rRegWrEn),
    .C(_0624_),
    .D(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__nor2_1 _1000_ (.A(\reg_s2[0] ),
    .B(_0595_),
    .Y(_0627_));
 sky130_fd_sc_hd__inv_2 _1001_ (.A(\reg_s2[0] ),
    .Y(_0628_));
 sky130_fd_sc_hd__nor2_1 _1002_ (.A(\rReg_d[0] ),
    .B(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__a2111oi_1 _1003_ (.A1(\rReg_d[1] ),
    .A2(_0621_),
    .B1(_0627_),
    .C1(_0629_),
    .D1(_0603_),
    .Y(_0630_));
 sky130_fd_sc_hd__and2_2 _1004_ (.A(_0626_),
    .B(_0630_),
    .X(_0631_));
 sky130_fd_sc_hd__nor2_1 _1005_ (.A(rHazardStallRs2),
    .B(net1508),
    .Y(_0632_));
 sky130_fd_sc_hd__o2111a_1 _1006_ (.A1(_0620_),
    .A2(_0631_),
    .B1(net1073),
    .C1(net1114),
    .D1(net1509),
    .X(wStall1));
 sky130_fd_sc_hd__nor2_1 _1007_ (.A(\funct3[0] ),
    .B(\funct3[1] ),
    .Y(wRamByteEn));
 sky130_fd_sc_hd__or4_1 _1008_ (.A(\wAluOut[21] ),
    .B(\wAluOut[20] ),
    .C(\wAluOut[23] ),
    .D(\wAluOut[22] ),
    .X(_0633_));
 sky130_fd_sc_hd__or4_1 _1009_ (.A(\wAluOut[17] ),
    .B(\wAluOut[16] ),
    .C(\wAluOut[19] ),
    .D(\wAluOut[18] ),
    .X(_0634_));
 sky130_fd_sc_hd__or4_1 _1010_ (.A(\wAluOut[29] ),
    .B(\wAluOut[28] ),
    .C(\wAluOut[31] ),
    .D(\wAluOut[30] ),
    .X(_0635_));
 sky130_fd_sc_hd__or4_1 _1011_ (.A(\wAluOut[25] ),
    .B(\wAluOut[24] ),
    .C(\wAluOut[27] ),
    .D(\wAluOut[26] ),
    .X(_0636_));
 sky130_fd_sc_hd__or4_1 _1012_ (.A(_0633_),
    .B(_0634_),
    .C(_0635_),
    .D(_0636_),
    .X(_0637_));
 sky130_fd_sc_hd__or4_1 _1013_ (.A(\wAluOut[5] ),
    .B(\wAluOut[4] ),
    .C(\wAluOut[7] ),
    .D(\wAluOut[6] ),
    .X(_0638_));
 sky130_fd_sc_hd__or4_1 _1014_ (.A(\wAluOut[1] ),
    .B(\wAluOut[0] ),
    .C(\wAluOut[3] ),
    .D(\wAluOut[2] ),
    .X(_0639_));
 sky130_fd_sc_hd__or4_1 _1015_ (.A(\wAluOut[13] ),
    .B(\wAluOut[12] ),
    .C(\wAluOut[15] ),
    .D(\wAluOut[14] ),
    .X(_0640_));
 sky130_fd_sc_hd__or4_1 _1016_ (.A(\wAluOut[9] ),
    .B(\wAluOut[8] ),
    .C(\wAluOut[11] ),
    .D(\wAluOut[10] ),
    .X(_0641_));
 sky130_fd_sc_hd__or4_1 _1017_ (.A(_0638_),
    .B(_0639_),
    .C(_0640_),
    .D(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__nor2_1 _1018_ (.A(_0637_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__nand2_1 _1019_ (.A(wRamWordEn),
    .B(net67),
    .Y(_0644_));
 sky130_fd_sc_hd__o21bai_1 _1020_ (.A1(wAluFlag),
    .A2(_0643_),
    .B1_N(_0644_),
    .Y(_0645_));
 sky130_fd_sc_hd__nor2_1 _1021_ (.A(wAluFlag),
    .B(_0643_),
    .Y(_0646_));
 sky130_fd_sc_hd__and3_1 _1022_ (.A(\funct3[0] ),
    .B(\funct3[1] ),
    .C(net67),
    .X(_0647_));
 sky130_fd_sc_hd__a21o_1 _1023_ (.A1(net67),
    .A2(wRamHalfEn),
    .B1(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__nand2_1 _1024_ (.A(_0646_),
    .B(_0648_),
    .Y(_0649_));
 sky130_fd_sc_hd__nand2_1 _1025_ (.A(_0645_),
    .B(_0649_),
    .Y(_0650_));
 sky130_fd_sc_hd__inv_2 _1026_ (.A(wAluFlag),
    .Y(_0651_));
 sky130_fd_sc_hd__nand2_1 _1027_ (.A(_0643_),
    .B(_0651_),
    .Y(_0652_));
 sky130_fd_sc_hd__inv_2 _1028_ (.A(net67),
    .Y(_0653_));
 sky130_fd_sc_hd__and2_1 _1029_ (.A(wRamHalfEn),
    .B(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__nand2_1 _1030_ (.A(_0652_),
    .B(_0654_),
    .Y(_0655_));
 sky130_fd_sc_hd__and2_1 _1031_ (.A(wRamByteEn),
    .B(_0653_),
    .X(_0656_));
 sky130_fd_sc_hd__nand3_1 _1032_ (.A(_0643_),
    .B(_0651_),
    .C(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__or3b_1 _1033_ (.A(_0651_),
    .B(_0653_),
    .C_N(wRamByteEn),
    .X(_0658_));
 sky130_fd_sc_hd__nand3_1 _1034_ (.A(_0655_),
    .B(_0657_),
    .C(_0658_),
    .Y(_0659_));
 sky130_fd_sc_hd__nor2_1 _1035_ (.A(_0650_),
    .B(_0659_),
    .Y(_0660_));
 sky130_fd_sc_hd__inv_2 _1036_ (.A(_0660_),
    .Y(wCond));
 sky130_fd_sc_hd__inv_2 _1037_ (.A(net896),
    .Y(_0661_));
 sky130_fd_sc_hd__buf_1 _1038_ (.A(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__inv_2 _1039_ (.A(net919),
    .Y(_0663_));
 sky130_fd_sc_hd__buf_1 _1040_ (.A(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1041_ (.A(_0664_),
    .X(_0665_));
 sky130_fd_sc_hd__nand2_2 _1042_ (.A(_0662_),
    .B(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__nor2_4 _1043_ (.A(_0592_),
    .B(_0666_),
    .Y(\wFunct3_aluIn[0] ));
 sky130_fd_sc_hd__nor2_2 _1044_ (.A(_0593_),
    .B(_0666_),
    .Y(\wFunct3_aluIn[1] ));
 sky130_fd_sc_hd__nor2_2 _1045_ (.A(_0653_),
    .B(_0666_),
    .Y(\wFunct3_aluIn[2] ));
 sky130_fd_sc_hd__and3_1 _1046_ (.A(_0662_),
    .B(_0665_),
    .C(\funct7[0] ),
    .X(_0667_));
 sky130_fd_sc_hd__buf_1 _1047_ (.A(_0667_),
    .X(\wFunct7_aluIn[0] ));
 sky130_fd_sc_hd__and3_1 _1048_ (.A(_0662_),
    .B(_0665_),
    .C(\funct7[1] ),
    .X(_0668_));
 sky130_fd_sc_hd__buf_1 _1049_ (.A(_0668_),
    .X(\wFunct7_aluIn[1] ));
 sky130_fd_sc_hd__and3_1 _1050_ (.A(_0662_),
    .B(_0665_),
    .C(\funct7[2] ),
    .X(_0669_));
 sky130_fd_sc_hd__buf_1 _1051_ (.A(_0669_),
    .X(\wFunct7_aluIn[2] ));
 sky130_fd_sc_hd__and3_1 _1052_ (.A(_0662_),
    .B(_0665_),
    .C(\funct7[3] ),
    .X(_0670_));
 sky130_fd_sc_hd__buf_1 _1053_ (.A(_0670_),
    .X(\wFunct7_aluIn[3] ));
 sky130_fd_sc_hd__buf_1 _1054_ (.A(_0663_),
    .X(_0671_));
 sky130_fd_sc_hd__and3_1 _1055_ (.A(_0662_),
    .B(_0671_),
    .C(\funct7[4] ),
    .X(_0672_));
 sky130_fd_sc_hd__buf_1 _1056_ (.A(_0672_),
    .X(\wFunct7_aluIn[4] ));
 sky130_fd_sc_hd__a21o_1 _1057_ (.A1(_0665_),
    .A2(\funct7[5] ),
    .B1(net896),
    .X(\wFunct7_aluIn[5] ));
 sky130_fd_sc_hd__and3_1 _1058_ (.A(_0661_),
    .B(_0671_),
    .C(\funct7[6] ),
    .X(_0673_));
 sky130_fd_sc_hd__buf_1 _1059_ (.A(_0673_),
    .X(\wFunct7_aluIn[6] ));
 sky130_fd_sc_hd__mux2_1 _1060_ (.A0(\rWrDataWB[0] ),
    .A1(net2),
    .S(net999),
    .X(_0674_));
 sky130_fd_sc_hd__clkbuf_1 _1061_ (.A(_0674_),
    .X(\wRegWrData[0] ));
 sky130_fd_sc_hd__mux2_2 _1062_ (.A0(\rWrDataWB[1] ),
    .A1(net13),
    .S(net1001),
    .X(_0675_));
 sky130_fd_sc_hd__buf_1 _1063_ (.A(_0675_),
    .X(\wRegWrData[1] ));
 sky130_fd_sc_hd__mux2_2 _1064_ (.A0(\rWrDataWB[2] ),
    .A1(net24),
    .S(net1002),
    .X(_0676_));
 sky130_fd_sc_hd__buf_1 _1065_ (.A(_0676_),
    .X(\wRegWrData[2] ));
 sky130_fd_sc_hd__mux2_2 _1066_ (.A0(\rWrDataWB[3] ),
    .A1(net27),
    .S(net1001),
    .X(_0677_));
 sky130_fd_sc_hd__buf_1 _1067_ (.A(_0677_),
    .X(\wRegWrData[3] ));
 sky130_fd_sc_hd__mux2_2 _1068_ (.A0(\rWrDataWB[4] ),
    .A1(net28),
    .S(net1000),
    .X(_0678_));
 sky130_fd_sc_hd__clkbuf_4 _1069_ (.A(_0678_),
    .X(\wRegWrData[4] ));
 sky130_fd_sc_hd__mux2_2 _1070_ (.A0(\rWrDataWB[5] ),
    .A1(net29),
    .S(net1001),
    .X(_0679_));
 sky130_fd_sc_hd__clkbuf_2 _1071_ (.A(_0679_),
    .X(\wRegWrData[5] ));
 sky130_fd_sc_hd__mux2_2 _1072_ (.A0(\rWrDataWB[6] ),
    .A1(net30),
    .S(net1001),
    .X(_0680_));
 sky130_fd_sc_hd__clkbuf_4 _1073_ (.A(_0680_),
    .X(\wRegWrData[6] ));
 sky130_fd_sc_hd__mux2_2 _1074_ (.A0(\rWrDataWB[7] ),
    .A1(net31),
    .S(net1000),
    .X(_0681_));
 sky130_fd_sc_hd__clkbuf_2 _1075_ (.A(_0681_),
    .X(\wRegWrData[7] ));
 sky130_fd_sc_hd__mux2_1 _1076_ (.A0(\rWrDataWB[8] ),
    .A1(net32),
    .S(net1001),
    .X(_0682_));
 sky130_fd_sc_hd__buf_2 _1077_ (.A(_0682_),
    .X(\wRegWrData[8] ));
 sky130_fd_sc_hd__mux2_2 _1078_ (.A0(\rWrDataWB[9] ),
    .A1(net33),
    .S(net1000),
    .X(_0683_));
 sky130_fd_sc_hd__clkbuf_2 _1079_ (.A(_0683_),
    .X(\wRegWrData[9] ));
 sky130_fd_sc_hd__mux2_2 _1080_ (.A0(\rWrDataWB[10] ),
    .A1(net3),
    .S(net1000),
    .X(_0684_));
 sky130_fd_sc_hd__clkbuf_2 _1081_ (.A(_0684_),
    .X(\wRegWrData[10] ));
 sky130_fd_sc_hd__mux2_1 _1082_ (.A0(\rWrDataWB[11] ),
    .A1(net4),
    .S(net1000),
    .X(_0685_));
 sky130_fd_sc_hd__clkbuf_2 _1083_ (.A(_0685_),
    .X(\wRegWrData[11] ));
 sky130_fd_sc_hd__mux2_1 _1084_ (.A0(\rWrDataWB[12] ),
    .A1(net5),
    .S(net999),
    .X(_0686_));
 sky130_fd_sc_hd__buf_4 _1085_ (.A(_0686_),
    .X(\wRegWrData[12] ));
 sky130_fd_sc_hd__mux2_1 _1086_ (.A0(\rWrDataWB[13] ),
    .A1(net6),
    .S(net999),
    .X(_0687_));
 sky130_fd_sc_hd__buf_2 _1087_ (.A(_0687_),
    .X(\wRegWrData[13] ));
 sky130_fd_sc_hd__mux2_1 _1088_ (.A0(\rWrDataWB[14] ),
    .A1(net7),
    .S(net999),
    .X(_0688_));
 sky130_fd_sc_hd__clkbuf_2 _1089_ (.A(_0688_),
    .X(\wRegWrData[14] ));
 sky130_fd_sc_hd__mux2_1 _1090_ (.A0(\rWrDataWB[15] ),
    .A1(net8),
    .S(net1002),
    .X(_0689_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1091_ (.A(_0689_),
    .X(\wRegWrData[15] ));
 sky130_fd_sc_hd__mux2_1 _1092_ (.A0(\rWrDataWB[16] ),
    .A1(net9),
    .S(net1000),
    .X(_0690_));
 sky130_fd_sc_hd__buf_4 _1093_ (.A(_0690_),
    .X(\wRegWrData[16] ));
 sky130_fd_sc_hd__mux2_1 _1094_ (.A0(\rWrDataWB[17] ),
    .A1(net10),
    .S(net1001),
    .X(_0691_));
 sky130_fd_sc_hd__clkbuf_2 _1095_ (.A(_0691_),
    .X(\wRegWrData[17] ));
 sky130_fd_sc_hd__mux2_1 _1096_ (.A0(\rWrDataWB[18] ),
    .A1(net11),
    .S(net999),
    .X(_0692_));
 sky130_fd_sc_hd__buf_1 _1097_ (.A(_0692_),
    .X(\wRegWrData[18] ));
 sky130_fd_sc_hd__mux2_1 _1098_ (.A0(\rWrDataWB[19] ),
    .A1(net12),
    .S(net998),
    .X(_0693_));
 sky130_fd_sc_hd__buf_1 _1099_ (.A(_0693_),
    .X(\wRegWrData[19] ));
 sky130_fd_sc_hd__mux2_1 _1100_ (.A0(\rWrDataWB[20] ),
    .A1(net14),
    .S(net999),
    .X(_0694_));
 sky130_fd_sc_hd__buf_1 _1101_ (.A(_0694_),
    .X(\wRegWrData[20] ));
 sky130_fd_sc_hd__mux2_1 _1102_ (.A0(\rWrDataWB[21] ),
    .A1(net15),
    .S(net998),
    .X(_0695_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1103_ (.A(_0695_),
    .X(\wRegWrData[21] ));
 sky130_fd_sc_hd__mux2_1 _1104_ (.A0(\rWrDataWB[22] ),
    .A1(net16),
    .S(net997),
    .X(_0696_));
 sky130_fd_sc_hd__buf_1 _1105_ (.A(_0696_),
    .X(\wRegWrData[22] ));
 sky130_fd_sc_hd__mux2_1 _1106_ (.A0(\rWrDataWB[23] ),
    .A1(net17),
    .S(net1003),
    .X(_0697_));
 sky130_fd_sc_hd__clkbuf_2 _1107_ (.A(_0697_),
    .X(\wRegWrData[23] ));
 sky130_fd_sc_hd__mux2_1 _1108_ (.A0(\rWrDataWB[24] ),
    .A1(net18),
    .S(net996),
    .X(_0698_));
 sky130_fd_sc_hd__clkbuf_2 _1109_ (.A(_0698_),
    .X(\wRegWrData[24] ));
 sky130_fd_sc_hd__mux2_1 _1110_ (.A0(\rWrDataWB[25] ),
    .A1(net19),
    .S(net996),
    .X(_0699_));
 sky130_fd_sc_hd__clkbuf_1 _1111_ (.A(_0699_),
    .X(\wRegWrData[25] ));
 sky130_fd_sc_hd__mux2_1 _1112_ (.A0(\rWrDataWB[26] ),
    .A1(net20),
    .S(net997),
    .X(_0700_));
 sky130_fd_sc_hd__clkbuf_1 _1113_ (.A(_0700_),
    .X(\wRegWrData[26] ));
 sky130_fd_sc_hd__mux2_2 _1114_ (.A0(\rWrDataWB[27] ),
    .A1(net21),
    .S(net998),
    .X(_0701_));
 sky130_fd_sc_hd__buf_1 _1115_ (.A(_0701_),
    .X(\wRegWrData[27] ));
 sky130_fd_sc_hd__mux2_1 _1116_ (.A0(\rWrDataWB[28] ),
    .A1(net22),
    .S(net996),
    .X(_0702_));
 sky130_fd_sc_hd__buf_2 _1117_ (.A(_0702_),
    .X(\wRegWrData[28] ));
 sky130_fd_sc_hd__mux2_1 _1118_ (.A0(\rWrDataWB[29] ),
    .A1(net23),
    .S(net996),
    .X(_0703_));
 sky130_fd_sc_hd__clkbuf_1 _1119_ (.A(_0703_),
    .X(\wRegWrData[29] ));
 sky130_fd_sc_hd__mux2_1 _1120_ (.A0(\rWrDataWB[30] ),
    .A1(net25),
    .S(net997),
    .X(_0704_));
 sky130_fd_sc_hd__buf_2 _1121_ (.A(_0704_),
    .X(\wRegWrData[30] ));
 sky130_fd_sc_hd__mux2_1 _1122_ (.A0(\rWrDataWB[31] ),
    .A1(net26),
    .S(net996),
    .X(_0705_));
 sky130_fd_sc_hd__buf_1 _1123_ (.A(_0705_),
    .X(\wRegWrData[31] ));
 sky130_fd_sc_hd__nand2b_1 _1124_ (.A_N(\reg_s1[1] ),
    .B(net994),
    .Y(_0706_));
 sky130_fd_sc_hd__nand2_1 _1125_ (.A(_0597_),
    .B(net995),
    .Y(_0707_));
 sky130_fd_sc_hd__inv_2 _1126_ (.A(net995),
    .Y(_0708_));
 sky130_fd_sc_hd__nand2_1 _1127_ (.A(_0708_),
    .B(\reg_s1[0] ),
    .Y(_0709_));
 sky130_fd_sc_hd__nand3_1 _1128_ (.A(_0706_),
    .B(_0707_),
    .C(_0709_),
    .Y(_0710_));
 sky130_fd_sc_hd__nand2_1 _1129_ (.A(_0608_),
    .B(net972),
    .Y(_0711_));
 sky130_fd_sc_hd__inv_2 _1130_ (.A(\rReg_d2[1] ),
    .Y(_0712_));
 sky130_fd_sc_hd__nand2_1 _1131_ (.A(_0712_),
    .B(\reg_s1[1] ),
    .Y(_0713_));
 sky130_fd_sc_hd__nand2_1 _1132_ (.A(_0711_),
    .B(_0713_),
    .Y(_0714_));
 sky130_fd_sc_hd__inv_2 _1133_ (.A(_0714_),
    .Y(_0715_));
 sky130_fd_sc_hd__inv_2 _1134_ (.A(\reg_s1[2] ),
    .Y(_0716_));
 sky130_fd_sc_hd__inv_4 _1135_ (.A(net987),
    .Y(_0717_));
 sky130_fd_sc_hd__nand2_1 _1136_ (.A(_0716_),
    .B(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__nand2_1 _1137_ (.A(\reg_s1[2] ),
    .B(net987),
    .Y(_0719_));
 sky130_fd_sc_hd__nand2_1 _1138_ (.A(_0718_),
    .B(_0719_),
    .Y(_0720_));
 sky130_fd_sc_hd__nand2_1 _1139_ (.A(_0715_),
    .B(_0720_),
    .Y(_0721_));
 sky130_fd_sc_hd__nor2_2 _1140_ (.A(_0710_),
    .B(_0721_),
    .Y(_0722_));
 sky130_fd_sc_hd__nand2_1 _1141_ (.A(_0708_),
    .B(_0712_),
    .Y(_0723_));
 sky130_fd_sc_hd__inv_4 _1142_ (.A(net962),
    .Y(_0724_));
 sky130_fd_sc_hd__nand3b_1 _1143_ (.A_N(net972),
    .B(_0717_),
    .C(_0724_),
    .Y(_0725_));
 sky130_fd_sc_hd__nor2_1 _1144_ (.A(_0723_),
    .B(_0725_),
    .Y(_0726_));
 sky130_fd_sc_hd__inv_2 _1145_ (.A(net996),
    .Y(_0727_));
 sky130_fd_sc_hd__nand2_1 _1146_ (.A(_0727_),
    .B(rRegWrEn2),
    .Y(_0728_));
 sky130_fd_sc_hd__nor2_1 _1147_ (.A(net972),
    .B(_0608_),
    .Y(_0729_));
 sky130_fd_sc_hd__nor2_1 _1148_ (.A(_0728_),
    .B(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__inv_2 _1149_ (.A(\reg_s1[4] ),
    .Y(_0731_));
 sky130_fd_sc_hd__nand2_1 _1150_ (.A(_0731_),
    .B(_0724_),
    .Y(_0732_));
 sky130_fd_sc_hd__nand2_1 _1151_ (.A(\reg_s1[4] ),
    .B(net962),
    .Y(_0733_));
 sky130_fd_sc_hd__nand2_1 _1152_ (.A(_0732_),
    .B(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__nand2_1 _1153_ (.A(_0730_),
    .B(_0734_),
    .Y(_0735_));
 sky130_fd_sc_hd__nor2_2 _1154_ (.A(_0726_),
    .B(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__nand2_1 _1155_ (.A(_0722_),
    .B(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__buf_6 _1156_ (.A(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__buf_6 _1157_ (.A(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__nand2_1 _1158_ (.A(_0739_),
    .B(\wRs1Data[0] ),
    .Y(_0740_));
 sky130_fd_sc_hd__clkbuf_2 _1159_ (.A(_0722_),
    .X(_0741_));
 sky130_fd_sc_hd__clkbuf_2 _1160_ (.A(_0736_),
    .X(_0742_));
 sky130_fd_sc_hd__nand3_1 _1161_ (.A(_0741_),
    .B(_0742_),
    .C(\rWrDataWB[0] ),
    .Y(_0743_));
 sky130_fd_sc_hd__buf_6 _1162_ (.A(_0616_),
    .X(_0744_));
 sky130_fd_sc_hd__buf_6 _1163_ (.A(_0744_),
    .X(_0745_));
 sky130_fd_sc_hd__nand3_2 _1164_ (.A(_0740_),
    .B(_0743_),
    .C(_0745_),
    .Y(_0746_));
 sky130_fd_sc_hd__inv_2 _1165_ (.A(\rWrData[0] ),
    .Y(_0747_));
 sky130_fd_sc_hd__nand2_1 _1166_ (.A(_0618_),
    .B(_0747_),
    .Y(_0748_));
 sky130_fd_sc_hd__a21o_1 _1167_ (.A1(_0746_),
    .A2(_0748_),
    .B1(\imm12_i_s[0] ),
    .X(_0749_));
 sky130_fd_sc_hd__nand3_2 _1168_ (.A(_0746_),
    .B(\imm12_i_s[0] ),
    .C(_0748_),
    .Y(_0750_));
 sky130_fd_sc_hd__nor2_2 _1169_ (.A(op_memSt),
    .B(op_memLd),
    .Y(_0751_));
 sky130_fd_sc_hd__inv_2 _1170_ (.A(_0751_),
    .Y(_0752_));
 sky130_fd_sc_hd__clkbuf_2 _1171_ (.A(_0752_),
    .X(_0753_));
 sky130_fd_sc_hd__and3_1 _1172_ (.A(_0749_),
    .B(_0750_),
    .C(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__buf_1 _1173_ (.A(_0754_),
    .X(net71));
 sky130_fd_sc_hd__inv_2 _1174_ (.A(\wRs1Data[1] ),
    .Y(_0755_));
 sky130_fd_sc_hd__nand2_1 _1175_ (.A(_0738_),
    .B(_0755_),
    .Y(_0756_));
 sky130_fd_sc_hd__inv_2 _1176_ (.A(\rWrDataWB[1] ),
    .Y(_0757_));
 sky130_fd_sc_hd__nand3_1 _1177_ (.A(_0722_),
    .B(_0736_),
    .C(_0757_),
    .Y(_0758_));
 sky130_fd_sc_hd__nand3_2 _1178_ (.A(_0756_),
    .B(_0758_),
    .C(_0744_),
    .Y(_0759_));
 sky130_fd_sc_hd__clkbuf_2 _1179_ (.A(_0617_),
    .X(_0760_));
 sky130_fd_sc_hd__nand2_1 _1180_ (.A(_0760_),
    .B(\rWrData[1] ),
    .Y(_0761_));
 sky130_fd_sc_hd__inv_2 _1181_ (.A(\imm12_i_s[1] ),
    .Y(_0762_));
 sky130_fd_sc_hd__a21o_1 _1182_ (.A1(_0759_),
    .A2(_0761_),
    .B1(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__nand3_1 _1183_ (.A(_0759_),
    .B(_0762_),
    .C(_0761_),
    .Y(_0764_));
 sky130_fd_sc_hd__and2_1 _1184_ (.A(_0763_),
    .B(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__or2b_1 _1185_ (.A(_0765_),
    .B_N(_0750_),
    .X(_0766_));
 sky130_fd_sc_hd__or2b_1 _1186_ (.A(_0750_),
    .B_N(_0765_),
    .X(_0767_));
 sky130_fd_sc_hd__and3_1 _1187_ (.A(_0766_),
    .B(_0767_),
    .C(_0752_),
    .X(_0768_));
 sky130_fd_sc_hd__clkbuf_1 _1188_ (.A(_0768_),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 _1189_ (.A(_0751_),
    .X(_0769_));
 sky130_fd_sc_hd__buf_6 _1190_ (.A(_0737_),
    .X(_0770_));
 sky130_fd_sc_hd__nand2_1 _1191_ (.A(_0770_),
    .B(\wRs1Data[2] ),
    .Y(_0771_));
 sky130_fd_sc_hd__nand3_1 _1192_ (.A(_0741_),
    .B(_0742_),
    .C(\rWrDataWB[2] ),
    .Y(_0772_));
 sky130_fd_sc_hd__nand3_2 _1193_ (.A(_0771_),
    .B(_0772_),
    .C(_0744_),
    .Y(_0773_));
 sky130_fd_sc_hd__inv_2 _1194_ (.A(\rWrData[2] ),
    .Y(_0774_));
 sky130_fd_sc_hd__nand2_1 _1195_ (.A(_0760_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__nand2_1 _1196_ (.A(_0773_),
    .B(_0775_),
    .Y(_0776_));
 sky130_fd_sc_hd__inv_2 _1197_ (.A(\imm12_i_s[2] ),
    .Y(_0777_));
 sky130_fd_sc_hd__nand2_1 _1198_ (.A(_0776_),
    .B(_0777_),
    .Y(_0778_));
 sky130_fd_sc_hd__nand3_1 _1199_ (.A(_0773_),
    .B(\imm12_i_s[2] ),
    .C(_0775_),
    .Y(_0779_));
 sky130_fd_sc_hd__nand2_1 _1200_ (.A(_0778_),
    .B(_0779_),
    .Y(_0780_));
 sky130_fd_sc_hd__inv_2 _1201_ (.A(_0764_),
    .Y(_0781_));
 sky130_fd_sc_hd__o21ai_2 _1202_ (.A1(_0750_),
    .A2(_0781_),
    .B1(_0763_),
    .Y(_0782_));
 sky130_fd_sc_hd__xor2_1 _1203_ (.A(_0780_),
    .B(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__nor2_1 _1204_ (.A(_0769_),
    .B(_0783_),
    .Y(net93));
 sky130_fd_sc_hd__inv_2 _1205_ (.A(\wRs1Data[3] ),
    .Y(_0784_));
 sky130_fd_sc_hd__nand2_1 _1206_ (.A(_0770_),
    .B(_0784_),
    .Y(_0785_));
 sky130_fd_sc_hd__inv_2 _1207_ (.A(\rWrDataWB[3] ),
    .Y(_0786_));
 sky130_fd_sc_hd__nand3_1 _1208_ (.A(_0741_),
    .B(_0742_),
    .C(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hd__nand3_1 _1209_ (.A(_0785_),
    .B(_0787_),
    .C(_0745_),
    .Y(_0788_));
 sky130_fd_sc_hd__nand2_1 _1210_ (.A(_0760_),
    .B(\rWrData[3] ),
    .Y(_0789_));
 sky130_fd_sc_hd__nand2_1 _1211_ (.A(_0788_),
    .B(_0789_),
    .Y(_0790_));
 sky130_fd_sc_hd__nand2_1 _1212_ (.A(_0790_),
    .B(\imm12_i_s[3] ),
    .Y(_0791_));
 sky130_fd_sc_hd__nand3b_1 _1213_ (.A_N(\imm12_i_s[3] ),
    .B(_0788_),
    .C(_0789_),
    .Y(_0792_));
 sky130_fd_sc_hd__nand2_1 _1214_ (.A(_0791_),
    .B(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__buf_2 _1215_ (.A(_0752_),
    .X(_0794_));
 sky130_fd_sc_hd__nor2_1 _1216_ (.A(_0780_),
    .B(_0793_),
    .Y(_0795_));
 sky130_fd_sc_hd__nand2_1 _1217_ (.A(_0782_),
    .B(_0795_),
    .Y(_0796_));
 sky130_fd_sc_hd__inv_2 _1218_ (.A(_0779_),
    .Y(_0797_));
 sky130_fd_sc_hd__inv_2 _1219_ (.A(_0793_),
    .Y(_0798_));
 sky130_fd_sc_hd__a211o_1 _1220_ (.A1(_0782_),
    .A2(_0778_),
    .B1(_0797_),
    .C1(_0798_),
    .X(_0799_));
 sky130_fd_sc_hd__o2111a_1 _1221_ (.A1(_0779_),
    .A2(_0793_),
    .B1(_0794_),
    .C1(_0796_),
    .D1(_0799_),
    .X(net96));
 sky130_fd_sc_hd__a21boi_1 _1222_ (.A1(_0797_),
    .A2(_0792_),
    .B1_N(_0791_),
    .Y(_0800_));
 sky130_fd_sc_hd__nand2_1 _1223_ (.A(_0796_),
    .B(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__inv_2 _1224_ (.A(\wRs1Data[4] ),
    .Y(_0802_));
 sky130_fd_sc_hd__nand2_1 _1225_ (.A(_0738_),
    .B(_0802_),
    .Y(_0803_));
 sky130_fd_sc_hd__inv_2 _1226_ (.A(\rWrDataWB[4] ),
    .Y(_0804_));
 sky130_fd_sc_hd__nand3_1 _1227_ (.A(_0741_),
    .B(_0736_),
    .C(_0804_),
    .Y(_0805_));
 sky130_fd_sc_hd__nand2_1 _1228_ (.A(_0803_),
    .B(_0805_),
    .Y(_0806_));
 sky130_fd_sc_hd__nand2_1 _1229_ (.A(_0806_),
    .B(_0744_),
    .Y(_0807_));
 sky130_fd_sc_hd__inv_2 _1230_ (.A(\rWrData[4] ),
    .Y(_0808_));
 sky130_fd_sc_hd__nand2_1 _1231_ (.A(_0760_),
    .B(_0808_),
    .Y(_0809_));
 sky130_fd_sc_hd__nand3_2 _1232_ (.A(_0807_),
    .B(\imm12_i_s[4] ),
    .C(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__nand3_1 _1233_ (.A(_0803_),
    .B(_0805_),
    .C(_0745_),
    .Y(_0811_));
 sky130_fd_sc_hd__nand2_1 _1234_ (.A(_0760_),
    .B(\rWrData[4] ),
    .Y(_0812_));
 sky130_fd_sc_hd__nand3b_1 _1235_ (.A_N(\imm12_i_s[4] ),
    .B(_0811_),
    .C(_0812_),
    .Y(_0813_));
 sky130_fd_sc_hd__nand2_1 _1236_ (.A(_0810_),
    .B(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__inv_2 _1237_ (.A(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__clkbuf_2 _1238_ (.A(_0752_),
    .X(_0816_));
 sky130_fd_sc_hd__o21ai_1 _1239_ (.A1(_0815_),
    .A2(_0801_),
    .B1(_0816_),
    .Y(_0817_));
 sky130_fd_sc_hd__a21oi_2 _1240_ (.A1(_0801_),
    .A2(_0815_),
    .B1(_0817_),
    .Y(net97));
 sky130_fd_sc_hd__inv_2 _1241_ (.A(\wRs1Data[5] ),
    .Y(_0818_));
 sky130_fd_sc_hd__nand2_1 _1242_ (.A(_0739_),
    .B(_0818_),
    .Y(_0819_));
 sky130_fd_sc_hd__inv_2 _1243_ (.A(\rWrDataWB[5] ),
    .Y(_0820_));
 sky130_fd_sc_hd__nand3_1 _1244_ (.A(_0741_),
    .B(_0742_),
    .C(_0820_),
    .Y(_0821_));
 sky130_fd_sc_hd__buf_6 _1245_ (.A(_0744_),
    .X(_0822_));
 sky130_fd_sc_hd__nand3_2 _1246_ (.A(_0819_),
    .B(_0821_),
    .C(_0822_),
    .Y(_0823_));
 sky130_fd_sc_hd__nand2_1 _1247_ (.A(_0618_),
    .B(\rWrData[5] ),
    .Y(_0824_));
 sky130_fd_sc_hd__a21o_1 _1248_ (.A1(_0823_),
    .A2(_0824_),
    .B1(\imm12_i_s[5] ),
    .X(_0825_));
 sky130_fd_sc_hd__nand3_1 _1249_ (.A(_0823_),
    .B(\imm12_i_s[5] ),
    .C(_0824_),
    .Y(_0826_));
 sky130_fd_sc_hd__nand2_1 _1250_ (.A(_0825_),
    .B(_0826_),
    .Y(_0827_));
 sky130_fd_sc_hd__inv_2 _1251_ (.A(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__nand2_1 _1252_ (.A(_0828_),
    .B(_0810_),
    .Y(_0829_));
 sky130_fd_sc_hd__a21o_1 _1253_ (.A1(_0801_),
    .A2(_0815_),
    .B1(_0829_),
    .X(_0830_));
 sky130_fd_sc_hd__nand2_1 _1254_ (.A(_0827_),
    .B(_0815_),
    .Y(_0831_));
 sky130_fd_sc_hd__a21o_1 _1255_ (.A1(_0796_),
    .A2(_0800_),
    .B1(_0831_),
    .X(_0832_));
 sky130_fd_sc_hd__nor2_1 _1256_ (.A(_0810_),
    .B(_0828_),
    .Y(_0833_));
 sky130_fd_sc_hd__inv_2 _1257_ (.A(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__and4_1 _1258_ (.A(_0830_),
    .B(_0752_),
    .C(_0832_),
    .D(_0834_),
    .X(_0835_));
 sky130_fd_sc_hd__clkbuf_1 _1259_ (.A(_0835_),
    .X(net98));
 sky130_fd_sc_hd__inv_2 _1260_ (.A(\wRs1Data[6] ),
    .Y(_0836_));
 sky130_fd_sc_hd__nand2_1 _1261_ (.A(_0738_),
    .B(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__nand3b_1 _1262_ (.A_N(\rWrDataWB[6] ),
    .B(_0722_),
    .C(_0742_),
    .Y(_0838_));
 sky130_fd_sc_hd__nand3_1 _1263_ (.A(_0837_),
    .B(_0838_),
    .C(_0745_),
    .Y(_0839_));
 sky130_fd_sc_hd__nand2_1 _1264_ (.A(_0618_),
    .B(\rWrData[6] ),
    .Y(_0840_));
 sky130_fd_sc_hd__nand3b_1 _1265_ (.A_N(\imm12_i_s[6] ),
    .B(_0839_),
    .C(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__nand2_1 _1266_ (.A(_0837_),
    .B(_0838_),
    .Y(_0842_));
 sky130_fd_sc_hd__nand2_1 _1267_ (.A(_0842_),
    .B(_0745_),
    .Y(_0843_));
 sky130_fd_sc_hd__or2_1 _1268_ (.A(\rWrData[6] ),
    .B(_0616_),
    .X(_0844_));
 sky130_fd_sc_hd__nand3_1 _1269_ (.A(_0843_),
    .B(\imm12_i_s[6] ),
    .C(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__nand2_1 _1270_ (.A(_0841_),
    .B(_0845_),
    .Y(_0846_));
 sky130_fd_sc_hd__inv_2 _1271_ (.A(_0846_),
    .Y(_0847_));
 sky130_fd_sc_hd__inv_2 _1272_ (.A(\imm12_i_s[5] ),
    .Y(_0848_));
 sky130_fd_sc_hd__a21o_1 _1273_ (.A1(_0823_),
    .A2(_0824_),
    .B1(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__nand3_1 _1274_ (.A(_0832_),
    .B(_0849_),
    .C(_0834_),
    .Y(_0850_));
 sky130_fd_sc_hd__or2_1 _1275_ (.A(_0847_),
    .B(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__nand2_1 _1276_ (.A(_0850_),
    .B(_0847_),
    .Y(_0852_));
 sky130_fd_sc_hd__nand3_1 _1277_ (.A(_0851_),
    .B(_0794_),
    .C(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__inv_2 _1278_ (.A(_0853_),
    .Y(net99));
 sky130_fd_sc_hd__inv_2 _1279_ (.A(\rWrData[7] ),
    .Y(_0854_));
 sky130_fd_sc_hd__buf_6 _1280_ (.A(_0745_),
    .X(_0855_));
 sky130_fd_sc_hd__inv_2 _1281_ (.A(\wRs1Data[7] ),
    .Y(_0856_));
 sky130_fd_sc_hd__nand2_1 _1282_ (.A(_0739_),
    .B(_0856_),
    .Y(_0857_));
 sky130_fd_sc_hd__inv_2 _1283_ (.A(\rWrDataWB[7] ),
    .Y(_0858_));
 sky130_fd_sc_hd__nand3_1 _1284_ (.A(_0741_),
    .B(_0742_),
    .C(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__nand3_2 _1285_ (.A(_0857_),
    .B(_0859_),
    .C(_0822_),
    .Y(_0860_));
 sky130_fd_sc_hd__o21ai_1 _1286_ (.A1(_0854_),
    .A2(_0855_),
    .B1(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__nand2_1 _1287_ (.A(_0861_),
    .B(\imm12_i_s[7] ),
    .Y(_0862_));
 sky130_fd_sc_hd__inv_2 _1288_ (.A(\imm12_i_s[7] ),
    .Y(_0863_));
 sky130_fd_sc_hd__o211ai_2 _1289_ (.A1(_0854_),
    .A2(_0822_),
    .B1(_0863_),
    .C1(_0860_),
    .Y(_0864_));
 sky130_fd_sc_hd__nand2_1 _1290_ (.A(_0862_),
    .B(_0864_),
    .Y(_0865_));
 sky130_fd_sc_hd__and2_1 _1291_ (.A(_0852_),
    .B(_0845_),
    .X(_0866_));
 sky130_fd_sc_hd__nor2_1 _1292_ (.A(_0865_),
    .B(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__nand2_1 _1293_ (.A(_0866_),
    .B(_0865_),
    .Y(_0868_));
 sky130_fd_sc_hd__nor3b_1 _1294_ (.A(_0769_),
    .B(_0867_),
    .C_N(_0868_),
    .Y(net100));
 sky130_fd_sc_hd__nand2_1 _1295_ (.A(_0861_),
    .B(_0863_),
    .Y(_0869_));
 sky130_fd_sc_hd__buf_4 _1296_ (.A(_0822_),
    .X(_0870_));
 sky130_fd_sc_hd__o211ai_1 _1297_ (.A1(_0854_),
    .A2(_0870_),
    .B1(\imm12_i_s[7] ),
    .C1(_0860_),
    .Y(_0871_));
 sky130_fd_sc_hd__nand2_1 _1298_ (.A(_0869_),
    .B(_0871_),
    .Y(_0872_));
 sky130_fd_sc_hd__nand2_1 _1299_ (.A(_0847_),
    .B(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__nor2_1 _1300_ (.A(_0873_),
    .B(_0831_),
    .Y(_0874_));
 sky130_fd_sc_hd__nand2_1 _1301_ (.A(_0801_),
    .B(_0874_),
    .Y(_0875_));
 sky130_fd_sc_hd__nor2_1 _1302_ (.A(_0846_),
    .B(_0865_),
    .Y(_0876_));
 sky130_fd_sc_hd__nand3_1 _1303_ (.A(_0823_),
    .B(_0848_),
    .C(_0824_),
    .Y(_0877_));
 sky130_fd_sc_hd__inv_2 _1304_ (.A(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__o21ai_1 _1305_ (.A1(_0810_),
    .A2(_0878_),
    .B1(_0849_),
    .Y(_0879_));
 sky130_fd_sc_hd__inv_2 _1306_ (.A(_0864_),
    .Y(_0880_));
 sky130_fd_sc_hd__o21ai_1 _1307_ (.A1(_0845_),
    .A2(_0880_),
    .B1(_0862_),
    .Y(_0881_));
 sky130_fd_sc_hd__a21oi_1 _1308_ (.A1(_0876_),
    .A2(_0879_),
    .B1(_0881_),
    .Y(_0882_));
 sky130_fd_sc_hd__nand2_1 _1309_ (.A(_0875_),
    .B(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__inv_2 _1310_ (.A(\rWrDataWB[8] ),
    .Y(_0884_));
 sky130_fd_sc_hd__buf_6 _1311_ (.A(_0738_),
    .X(_0885_));
 sky130_fd_sc_hd__nor2_1 _1312_ (.A(_0884_),
    .B(_0885_),
    .Y(_0886_));
 sky130_fd_sc_hd__and2_1 _1313_ (.A(_0770_),
    .B(\wRs1Data[8] ),
    .X(_0887_));
 sky130_fd_sc_hd__o21ai_2 _1314_ (.A1(_0886_),
    .A2(_0887_),
    .B1(_0855_),
    .Y(_0888_));
 sky130_fd_sc_hd__clkbuf_2 _1315_ (.A(_0760_),
    .X(_0889_));
 sky130_fd_sc_hd__nand2_1 _1316_ (.A(_0889_),
    .B(\rWrData[8] ),
    .Y(_0890_));
 sky130_fd_sc_hd__nand2_1 _1317_ (.A(_0888_),
    .B(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__nand2_1 _1318_ (.A(_0891_),
    .B(\imm12_i_s[8] ),
    .Y(_0892_));
 sky130_fd_sc_hd__nand3b_1 _1319_ (.A_N(\imm12_i_s[8] ),
    .B(_0888_),
    .C(_0890_),
    .Y(_0893_));
 sky130_fd_sc_hd__nand2_1 _1320_ (.A(_0892_),
    .B(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__inv_2 _1321_ (.A(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__and2_1 _1322_ (.A(_0883_),
    .B(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__nor2_1 _1323_ (.A(_0769_),
    .B(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__o21ai_1 _1324_ (.A1(_0883_),
    .A2(_0895_),
    .B1(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__inv_2 _1325_ (.A(_0898_),
    .Y(net101));
 sky130_fd_sc_hd__buf_6 _1326_ (.A(_0822_),
    .X(_0899_));
 sky130_fd_sc_hd__inv_2 _1327_ (.A(\rWrDataWB[9] ),
    .Y(_0900_));
 sky130_fd_sc_hd__nor2_1 _1328_ (.A(_0900_),
    .B(_0885_),
    .Y(_0901_));
 sky130_fd_sc_hd__and2_1 _1329_ (.A(_0770_),
    .B(\wRs1Data[9] ),
    .X(_0902_));
 sky130_fd_sc_hd__nor2_1 _1330_ (.A(_0901_),
    .B(_0902_),
    .Y(_0903_));
 sky130_fd_sc_hd__nand2_1 _1331_ (.A(_0903_),
    .B(_0870_),
    .Y(_0904_));
 sky130_fd_sc_hd__o211ai_2 _1332_ (.A1(\rWrData[9] ),
    .A2(_0899_),
    .B1(\imm12_i_s[9] ),
    .C1(_0904_),
    .Y(_0905_));
 sky130_fd_sc_hd__o21ai_1 _1333_ (.A1(_0901_),
    .A2(_0902_),
    .B1(_0855_),
    .Y(_0906_));
 sky130_fd_sc_hd__inv_2 _1334_ (.A(\imm12_i_s[9] ),
    .Y(_0907_));
 sky130_fd_sc_hd__nand2_1 _1335_ (.A(_0889_),
    .B(\rWrData[9] ),
    .Y(_0908_));
 sky130_fd_sc_hd__nand3_1 _1336_ (.A(_0906_),
    .B(_0907_),
    .C(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__nand2_1 _1337_ (.A(_0905_),
    .B(_0909_),
    .Y(_0910_));
 sky130_fd_sc_hd__nor2_1 _1338_ (.A(_0894_),
    .B(_0910_),
    .Y(_0911_));
 sky130_fd_sc_hd__nand2_1 _1339_ (.A(_0883_),
    .B(_0911_),
    .Y(_0912_));
 sky130_fd_sc_hd__nand2_1 _1340_ (.A(_0910_),
    .B(_0892_),
    .Y(_0913_));
 sky130_fd_sc_hd__clkbuf_2 _1341_ (.A(_0752_),
    .X(_0914_));
 sky130_fd_sc_hd__o21a_1 _1342_ (.A1(_0913_),
    .A2(_0896_),
    .B1(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__o211a_1 _1343_ (.A1(_0892_),
    .A2(_0910_),
    .B1(_0912_),
    .C1(_0915_),
    .X(net102));
 sky130_fd_sc_hd__inv_2 _1344_ (.A(_0909_),
    .Y(_0916_));
 sky130_fd_sc_hd__o21ai_1 _1345_ (.A1(_0892_),
    .A2(_0916_),
    .B1(_0905_),
    .Y(_0917_));
 sky130_fd_sc_hd__inv_2 _1346_ (.A(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__inv_2 _1347_ (.A(\rWrDataWB[10] ),
    .Y(_0919_));
 sky130_fd_sc_hd__nor2_1 _1348_ (.A(_0919_),
    .B(_0885_),
    .Y(_0920_));
 sky130_fd_sc_hd__and2_1 _1349_ (.A(_0770_),
    .B(\wRs1Data[10] ),
    .X(_0921_));
 sky130_fd_sc_hd__o21ai_1 _1350_ (.A1(_0920_),
    .A2(_0921_),
    .B1(_0870_),
    .Y(_0922_));
 sky130_fd_sc_hd__clkbuf_2 _1351_ (.A(_0618_),
    .X(_0923_));
 sky130_fd_sc_hd__nand2_1 _1352_ (.A(_0923_),
    .B(\rWrData[10] ),
    .Y(_0924_));
 sky130_fd_sc_hd__nand3b_1 _1353_ (.A_N(\imm12_i_s[10] ),
    .B(_0922_),
    .C(_0924_),
    .Y(_0925_));
 sky130_fd_sc_hd__nor2_1 _1354_ (.A(_0920_),
    .B(_0921_),
    .Y(_0926_));
 sky130_fd_sc_hd__nand2_1 _1355_ (.A(_0926_),
    .B(_0870_),
    .Y(_0927_));
 sky130_fd_sc_hd__inv_2 _1356_ (.A(\rWrData[10] ),
    .Y(_0928_));
 sky130_fd_sc_hd__nand2_1 _1357_ (.A(_0923_),
    .B(_0928_),
    .Y(_0929_));
 sky130_fd_sc_hd__nand3_2 _1358_ (.A(_0927_),
    .B(\imm12_i_s[10] ),
    .C(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__nand2_1 _1359_ (.A(_0925_),
    .B(_0930_),
    .Y(_0931_));
 sky130_fd_sc_hd__nand2_1 _1360_ (.A(_0912_),
    .B(_0918_),
    .Y(_0932_));
 sky130_fd_sc_hd__inv_2 _1361_ (.A(_0931_),
    .Y(_0933_));
 sky130_fd_sc_hd__nand2_1 _1362_ (.A(_0932_),
    .B(_0933_),
    .Y(_0934_));
 sky130_fd_sc_hd__nand2_1 _1363_ (.A(_0934_),
    .B(_0753_),
    .Y(_0935_));
 sky130_fd_sc_hd__a31o_1 _1364_ (.A1(_0912_),
    .A2(_0918_),
    .A3(_0931_),
    .B1(_0935_),
    .X(_0936_));
 sky130_fd_sc_hd__inv_2 _1365_ (.A(_0936_),
    .Y(net72));
 sky130_fd_sc_hd__inv_2 _1366_ (.A(\rWrDataWB[11] ),
    .Y(_0937_));
 sky130_fd_sc_hd__clkbuf_2 _1367_ (.A(_0738_),
    .X(_0938_));
 sky130_fd_sc_hd__nand2_1 _1368_ (.A(_0739_),
    .B(\wRs1Data[11] ),
    .Y(_0939_));
 sky130_fd_sc_hd__o211ai_2 _1369_ (.A1(_0937_),
    .A2(_0938_),
    .B1(_0870_),
    .C1(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__o211ai_2 _1370_ (.A1(\rWrData[11] ),
    .A2(_0899_),
    .B1(\imm12_i_s[11] ),
    .C1(_0940_),
    .Y(_0941_));
 sky130_fd_sc_hd__o21ai_1 _1371_ (.A1(_0937_),
    .A2(_0938_),
    .B1(_0939_),
    .Y(_0942_));
 sky130_fd_sc_hd__nand2_1 _1372_ (.A(_0942_),
    .B(_0855_),
    .Y(_0943_));
 sky130_fd_sc_hd__inv_2 _1373_ (.A(\imm12_i_s[11] ),
    .Y(_0944_));
 sky130_fd_sc_hd__nand2_1 _1374_ (.A(_0889_),
    .B(\rWrData[11] ),
    .Y(_0945_));
 sky130_fd_sc_hd__nand3_1 _1375_ (.A(_0943_),
    .B(_0944_),
    .C(_0945_),
    .Y(_0946_));
 sky130_fd_sc_hd__nand2_1 _1376_ (.A(_0941_),
    .B(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__a21oi_1 _1377_ (.A1(_0934_),
    .A2(_0930_),
    .B1(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__a31o_1 _1378_ (.A1(_0934_),
    .A2(_0930_),
    .A3(_0947_),
    .B1(_0769_),
    .X(_0949_));
 sky130_fd_sc_hd__nor2_1 _1379_ (.A(_0948_),
    .B(_0949_),
    .Y(net73));
 sky130_fd_sc_hd__inv_2 _1380_ (.A(_0737_),
    .Y(_0950_));
 sky130_fd_sc_hd__clkbuf_2 _1381_ (.A(_0950_),
    .X(_0951_));
 sky130_fd_sc_hd__or2_1 _1382_ (.A(\rWrDataWB[12] ),
    .B(_0770_),
    .X(_0952_));
 sky130_fd_sc_hd__o21ai_1 _1383_ (.A1(\wRs1Data[12] ),
    .A2(_0951_),
    .B1(_0952_),
    .Y(_0953_));
 sky130_fd_sc_hd__or2_1 _1384_ (.A(\rWrData[12] ),
    .B(_0744_),
    .X(_0954_));
 sky130_fd_sc_hd__inv_2 _1385_ (.A(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__a21o_1 _1386_ (.A1(_0953_),
    .A2(_0855_),
    .B1(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__inv_2 _1387_ (.A(_0956_),
    .Y(_0957_));
 sky130_fd_sc_hd__nor2_1 _1388_ (.A(_0931_),
    .B(_0947_),
    .Y(_0958_));
 sky130_fd_sc_hd__and2_1 _1389_ (.A(_0911_),
    .B(_0958_),
    .X(_0959_));
 sky130_fd_sc_hd__nand2_1 _1390_ (.A(_0917_),
    .B(_0958_),
    .Y(_0960_));
 sky130_fd_sc_hd__inv_2 _1391_ (.A(_0946_),
    .Y(_0961_));
 sky130_fd_sc_hd__o21a_1 _1392_ (.A1(_0930_),
    .A2(_0961_),
    .B1(_0941_),
    .X(_0962_));
 sky130_fd_sc_hd__nand2_1 _1393_ (.A(_0960_),
    .B(_0962_),
    .Y(_0035_));
 sky130_fd_sc_hd__a21o_1 _1394_ (.A1(_0883_),
    .A2(_0959_),
    .B1(_0035_),
    .X(_0036_));
 sky130_fd_sc_hd__or2_1 _1395_ (.A(_0957_),
    .B(_0036_),
    .X(_0037_));
 sky130_fd_sc_hd__nand2_1 _1396_ (.A(_0036_),
    .B(_0957_),
    .Y(_0038_));
 sky130_fd_sc_hd__nand3_1 _1397_ (.A(_0037_),
    .B(_0794_),
    .C(_0038_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _1398_ (.A(_0039_),
    .Y(net74));
 sky130_fd_sc_hd__and2_1 _1399_ (.A(_0739_),
    .B(\wRs1Data[13] ),
    .X(_0040_));
 sky130_fd_sc_hd__a21o_1 _1400_ (.A1(_0951_),
    .A2(\rWrDataWB[13] ),
    .B1(_0618_),
    .X(_0041_));
 sky130_fd_sc_hd__o22ai_4 _1401_ (.A1(\rWrData[13] ),
    .A2(_0855_),
    .B1(_0040_),
    .B2(_0041_),
    .Y(_0042_));
 sky130_fd_sc_hd__nand2_1 _1402_ (.A(_0038_),
    .B(_0042_),
    .Y(_0043_));
 sky130_fd_sc_hd__nor2_1 _1403_ (.A(_0042_),
    .B(_0956_),
    .Y(_0044_));
 sky130_fd_sc_hd__nand2_1 _1404_ (.A(_0036_),
    .B(_0044_),
    .Y(_0045_));
 sky130_fd_sc_hd__and3_1 _1405_ (.A(_0043_),
    .B(_0914_),
    .C(_0045_),
    .X(_0046_));
 sky130_fd_sc_hd__clkbuf_1 _1406_ (.A(_0046_),
    .X(net75));
 sky130_fd_sc_hd__nor2_1 _1407_ (.A(\rWrDataWB[14] ),
    .B(_0885_),
    .Y(_0047_));
 sky130_fd_sc_hd__nor2_1 _1408_ (.A(\wRs1Data[14] ),
    .B(_0951_),
    .Y(_0048_));
 sky130_fd_sc_hd__nand2_1 _1409_ (.A(_0889_),
    .B(\rWrData[14] ),
    .Y(_0049_));
 sky130_fd_sc_hd__o31a_2 _1410_ (.A1(_0889_),
    .A2(_0047_),
    .A3(_0048_),
    .B1(_0049_),
    .X(_0050_));
 sky130_fd_sc_hd__and2_1 _1411_ (.A(_0045_),
    .B(_0050_),
    .X(_0051_));
 sky130_fd_sc_hd__or2_1 _1412_ (.A(_0050_),
    .B(_0045_),
    .X(_0052_));
 sky130_fd_sc_hd__nand2_1 _1413_ (.A(_0052_),
    .B(_0794_),
    .Y(_0053_));
 sky130_fd_sc_hd__nor2_1 _1414_ (.A(_0051_),
    .B(_0053_),
    .Y(net76));
 sky130_fd_sc_hd__and2_1 _1415_ (.A(_0885_),
    .B(\wRs1Data[15] ),
    .X(_0054_));
 sky130_fd_sc_hd__a21o_1 _1416_ (.A1(_0951_),
    .A2(net307),
    .B1(_0889_),
    .X(_0055_));
 sky130_fd_sc_hd__o22ai_4 _1417_ (.A1(\rWrData[15] ),
    .A2(_0870_),
    .B1(_0054_),
    .B2(_0055_),
    .Y(_0056_));
 sky130_fd_sc_hd__nor2_1 _1418_ (.A(_0056_),
    .B(_0050_),
    .Y(_0057_));
 sky130_fd_sc_hd__nand2_1 _1419_ (.A(_0057_),
    .B(_0044_),
    .Y(_0058_));
 sky130_fd_sc_hd__nand2_1 _1420_ (.A(_0911_),
    .B(_0958_),
    .Y(_0059_));
 sky130_fd_sc_hd__nor2_1 _1421_ (.A(_0058_),
    .B(_0059_),
    .Y(_0060_));
 sky130_fd_sc_hd__nand2_1 _1422_ (.A(_0883_),
    .B(_0060_),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _1423_ (.A(_0058_),
    .Y(_0062_));
 sky130_fd_sc_hd__nand2_1 _1424_ (.A(_0035_),
    .B(_0062_),
    .Y(_0063_));
 sky130_fd_sc_hd__nand2_2 _1425_ (.A(_0061_),
    .B(_0063_),
    .Y(_0064_));
 sky130_fd_sc_hd__buf_6 _1426_ (.A(_0064_),
    .X(_0065_));
 sky130_fd_sc_hd__or2_1 _1427_ (.A(_0769_),
    .B(_0065_),
    .X(_0066_));
 sky130_fd_sc_hd__a21oi_1 _1428_ (.A1(_0052_),
    .A2(_0056_),
    .B1(_0066_),
    .Y(net77));
 sky130_fd_sc_hd__inv_2 _1429_ (.A(\rWrData[16] ),
    .Y(_0067_));
 sky130_fd_sc_hd__clkbuf_4 _1430_ (.A(_0899_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1431_ (.A0(\rWrDataWB[16] ),
    .A1(\wRs1Data[16] ),
    .S(_0938_),
    .X(_0069_));
 sky130_fd_sc_hd__nand2_1 _1432_ (.A(_0069_),
    .B(_0068_),
    .Y(_0070_));
 sky130_fd_sc_hd__o21ai_2 _1433_ (.A1(_0067_),
    .A2(_0068_),
    .B1(_0070_),
    .Y(_0071_));
 sky130_fd_sc_hd__or2_1 _1434_ (.A(_0071_),
    .B(_0065_),
    .X(_0072_));
 sky130_fd_sc_hd__nand2_1 _1435_ (.A(_0064_),
    .B(_0071_),
    .Y(_0073_));
 sky130_fd_sc_hd__nand3_1 _1436_ (.A(_0072_),
    .B(_0794_),
    .C(_0073_),
    .Y(_0074_));
 sky130_fd_sc_hd__inv_2 _1437_ (.A(_0074_),
    .Y(net78));
 sky130_fd_sc_hd__clkbuf_2 _1438_ (.A(_0950_),
    .X(_0075_));
 sky130_fd_sc_hd__clkbuf_2 _1439_ (.A(_0885_),
    .X(_0076_));
 sky130_fd_sc_hd__or2_1 _1440_ (.A(\rWrDataWB[17] ),
    .B(_0076_),
    .X(_0077_));
 sky130_fd_sc_hd__o21ai_1 _1441_ (.A1(\wRs1Data[17] ),
    .A2(_0075_),
    .B1(_0077_),
    .Y(_0078_));
 sky130_fd_sc_hd__or2_1 _1442_ (.A(\rWrData[17] ),
    .B(_0822_),
    .X(_0079_));
 sky130_fd_sc_hd__inv_2 _1443_ (.A(_0079_),
    .Y(_0080_));
 sky130_fd_sc_hd__a21oi_2 _1444_ (.A1(_0078_),
    .A2(_0068_),
    .B1(_0080_),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _1445_ (.A(_0081_),
    .Y(_0082_));
 sky130_fd_sc_hd__or2_1 _1446_ (.A(_0082_),
    .B(_0073_),
    .X(_0083_));
 sky130_fd_sc_hd__nand2_1 _1447_ (.A(_0073_),
    .B(_0082_),
    .Y(_0084_));
 sky130_fd_sc_hd__and3_1 _1448_ (.A(_0083_),
    .B(_0753_),
    .C(_0084_),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_1 _1449_ (.A(_0085_),
    .X(net79));
 sky130_fd_sc_hd__inv_2 _1450_ (.A(\rWrData[18] ),
    .Y(_0086_));
 sky130_fd_sc_hd__buf_2 _1451_ (.A(_0899_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _1452_ (.A0(\rWrDataWB[18] ),
    .A1(\wRs1Data[18] ),
    .S(_0076_),
    .X(_0088_));
 sky130_fd_sc_hd__nand2_1 _1453_ (.A(_0088_),
    .B(_0087_),
    .Y(_0089_));
 sky130_fd_sc_hd__o21ai_2 _1454_ (.A1(_0086_),
    .A2(_0087_),
    .B1(_0089_),
    .Y(_0090_));
 sky130_fd_sc_hd__inv_2 _1455_ (.A(_0090_),
    .Y(_0091_));
 sky130_fd_sc_hd__nand2_1 _1456_ (.A(_0071_),
    .B(_0081_),
    .Y(_0092_));
 sky130_fd_sc_hd__nor2_1 _1457_ (.A(_0091_),
    .B(_0092_),
    .Y(_0093_));
 sky130_fd_sc_hd__nand2_1 _1458_ (.A(_0065_),
    .B(_0093_),
    .Y(_0094_));
 sky130_fd_sc_hd__nand2_1 _1459_ (.A(_0094_),
    .B(_0816_),
    .Y(_0095_));
 sky130_fd_sc_hd__a21oi_1 _1460_ (.A1(_0083_),
    .A2(_0091_),
    .B1(_0095_),
    .Y(net80));
 sky130_fd_sc_hd__clkbuf_2 _1461_ (.A(_0938_),
    .X(_0096_));
 sky130_fd_sc_hd__or2_1 _1462_ (.A(\wRs1Data[19] ),
    .B(_0075_),
    .X(_0097_));
 sky130_fd_sc_hd__o21ai_1 _1463_ (.A1(\rWrDataWB[19] ),
    .A2(_0096_),
    .B1(_0097_),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _1464_ (.A(\rWrData[19] ),
    .Y(_0099_));
 sky130_fd_sc_hd__nand2_1 _1465_ (.A(_0923_),
    .B(_0099_),
    .Y(_0100_));
 sky130_fd_sc_hd__inv_2 _1466_ (.A(_0100_),
    .Y(_0101_));
 sky130_fd_sc_hd__a21oi_2 _1467_ (.A1(_0098_),
    .A2(_0068_),
    .B1(_0101_),
    .Y(_0102_));
 sky130_fd_sc_hd__a21o_1 _1468_ (.A1(_0065_),
    .A2(_0093_),
    .B1(_0102_),
    .X(_0103_));
 sky130_fd_sc_hd__nand2_1 _1469_ (.A(_0090_),
    .B(_0102_),
    .Y(_0104_));
 sky130_fd_sc_hd__nor2_1 _1470_ (.A(_0092_),
    .B(_0104_),
    .Y(_0105_));
 sky130_fd_sc_hd__nand2_1 _1471_ (.A(_0064_),
    .B(_0105_),
    .Y(_0106_));
 sky130_fd_sc_hd__and3_1 _1472_ (.A(_0103_),
    .B(_0753_),
    .C(_0106_),
    .X(_0107_));
 sky130_fd_sc_hd__clkbuf_1 _1473_ (.A(_0107_),
    .X(net81));
 sky130_fd_sc_hd__and2_1 _1474_ (.A(_0938_),
    .B(\wRs1Data[20] ),
    .X(_0108_));
 sky130_fd_sc_hd__a211o_1 _1475_ (.A1(_0075_),
    .A2(\rWrDataWB[20] ),
    .B1(_0923_),
    .C1(_0108_),
    .X(_0109_));
 sky130_fd_sc_hd__o21ai_4 _1476_ (.A1(\rWrData[20] ),
    .A2(_0068_),
    .B1(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__or2_1 _1477_ (.A(_0110_),
    .B(_0106_),
    .X(_0111_));
 sky130_fd_sc_hd__nand2_1 _1478_ (.A(_0106_),
    .B(_0110_),
    .Y(_0112_));
 sky130_fd_sc_hd__and3_1 _1479_ (.A(_0111_),
    .B(_0753_),
    .C(_0112_),
    .X(_0113_));
 sky130_fd_sc_hd__clkbuf_1 _1480_ (.A(_0113_),
    .X(net83));
 sky130_fd_sc_hd__a21o_1 _1481_ (.A1(_0075_),
    .A2(net301),
    .B1(_0923_),
    .X(_0114_));
 sky130_fd_sc_hd__a21o_1 _1482_ (.A1(\wRs1Data[21] ),
    .A2(_0096_),
    .B1(_0114_),
    .X(_0115_));
 sky130_fd_sc_hd__o21ai_4 _1483_ (.A1(\rWrData[21] ),
    .A2(_0068_),
    .B1(_0115_),
    .Y(_0116_));
 sky130_fd_sc_hd__nor2_1 _1484_ (.A(_0116_),
    .B(_0110_),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _1485_ (.A(_0117_),
    .Y(_0118_));
 sky130_fd_sc_hd__or2_1 _1486_ (.A(_0118_),
    .B(_0106_),
    .X(_0119_));
 sky130_fd_sc_hd__nand2_1 _1487_ (.A(_0119_),
    .B(_0914_),
    .Y(_0120_));
 sky130_fd_sc_hd__a21oi_1 _1488_ (.A1(_0111_),
    .A2(_0116_),
    .B1(_0120_),
    .Y(net84));
 sky130_fd_sc_hd__clkbuf_2 _1489_ (.A(_0951_),
    .X(_0121_));
 sky130_fd_sc_hd__and2_1 _1490_ (.A(_0076_),
    .B(\wRs1Data[22] ),
    .X(_0122_));
 sky130_fd_sc_hd__a211o_1 _1491_ (.A1(_0121_),
    .A2(\rWrDataWB[22] ),
    .B1(_0619_),
    .C1(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__o21ai_4 _1492_ (.A1(\rWrData[22] ),
    .A2(_0087_),
    .B1(_0123_),
    .Y(_0124_));
 sky130_fd_sc_hd__or2_1 _1493_ (.A(_0124_),
    .B(_0118_),
    .X(_0125_));
 sky130_fd_sc_hd__or2_1 _1494_ (.A(_0125_),
    .B(_0106_),
    .X(_0126_));
 sky130_fd_sc_hd__nand2_1 _1495_ (.A(_0126_),
    .B(_0914_),
    .Y(_0127_));
 sky130_fd_sc_hd__a21oi_1 _1496_ (.A1(_0119_),
    .A2(_0124_),
    .B1(_0127_),
    .Y(net85));
 sky130_fd_sc_hd__and2_1 _1497_ (.A(_0739_),
    .B(\wRs1Data[23] ),
    .X(_0128_));
 sky130_fd_sc_hd__a21o_1 _1498_ (.A1(\rWrDataWB[23] ),
    .A2(_0951_),
    .B1(_0128_),
    .X(_0129_));
 sky130_fd_sc_hd__nand2_1 _1499_ (.A(_0923_),
    .B(\rWrData[23] ),
    .Y(_0130_));
 sky130_fd_sc_hd__a21bo_1 _1500_ (.A1(_0129_),
    .A2(_0899_),
    .B1_N(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__inv_2 _1501_ (.A(_0131_),
    .Y(_0132_));
 sky130_fd_sc_hd__nand3_1 _1502_ (.A(_0093_),
    .B(_0102_),
    .C(_0131_),
    .Y(_0133_));
 sky130_fd_sc_hd__nor2_1 _1503_ (.A(_0133_),
    .B(_0125_),
    .Y(_0134_));
 sky130_fd_sc_hd__nand2_1 _1504_ (.A(_0134_),
    .B(_0065_),
    .Y(_0135_));
 sky130_fd_sc_hd__nand2_1 _1505_ (.A(_0135_),
    .B(_0914_),
    .Y(_0136_));
 sky130_fd_sc_hd__a21oi_2 _1506_ (.A1(_0126_),
    .A2(_0132_),
    .B1(_0136_),
    .Y(net86));
 sky130_fd_sc_hd__nand2_1 _1507_ (.A(_0121_),
    .B(\rWrDataWB[24] ),
    .Y(_0137_));
 sky130_fd_sc_hd__nand2_1 _1508_ (.A(_0096_),
    .B(\wRs1Data[24] ),
    .Y(_0138_));
 sky130_fd_sc_hd__nand2_1 _1509_ (.A(_0137_),
    .B(_0138_),
    .Y(_0139_));
 sky130_fd_sc_hd__nand2_1 _1510_ (.A(_0619_),
    .B(\rWrData[24] ),
    .Y(_0140_));
 sky130_fd_sc_hd__a21bo_2 _1511_ (.A1(_0139_),
    .A2(_0087_),
    .B1_N(_0140_),
    .X(_0141_));
 sky130_fd_sc_hd__inv_2 _1512_ (.A(_0141_),
    .Y(_0142_));
 sky130_fd_sc_hd__nand2_1 _1513_ (.A(_0135_),
    .B(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__nor2_1 _1514_ (.A(_0110_),
    .B(_0132_),
    .Y(_0144_));
 sky130_fd_sc_hd__nor2_1 _1515_ (.A(_0116_),
    .B(_0124_),
    .Y(_0145_));
 sky130_fd_sc_hd__nand3_1 _1516_ (.A(_0105_),
    .B(_0144_),
    .C(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__inv_2 _1517_ (.A(_0146_),
    .Y(_0147_));
 sky130_fd_sc_hd__nand3_1 _1518_ (.A(_0064_),
    .B(_0141_),
    .C(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__and3_1 _1519_ (.A(_0143_),
    .B(_0753_),
    .C(_0148_),
    .X(_0149_));
 sky130_fd_sc_hd__clkbuf_1 _1520_ (.A(_0149_),
    .X(net87));
 sky130_fd_sc_hd__and2_1 _1521_ (.A(_0076_),
    .B(\wRs1Data[25] ),
    .X(_0150_));
 sky130_fd_sc_hd__a21o_1 _1522_ (.A1(\rWrDataWB[25] ),
    .A2(_0121_),
    .B1(_0150_),
    .X(_0151_));
 sky130_fd_sc_hd__nand2_1 _1523_ (.A(_0619_),
    .B(\rWrData[25] ),
    .Y(_0152_));
 sky130_fd_sc_hd__a21bo_1 _1524_ (.A1(_0151_),
    .A2(_0087_),
    .B1_N(_0152_),
    .X(_0153_));
 sky130_fd_sc_hd__inv_2 _1525_ (.A(_0153_),
    .Y(_0154_));
 sky130_fd_sc_hd__nor2_1 _1526_ (.A(_0154_),
    .B(_0148_),
    .Y(_0155_));
 sky130_fd_sc_hd__a21o_1 _1527_ (.A1(_0148_),
    .A2(_0154_),
    .B1(_0769_),
    .X(_0156_));
 sky130_fd_sc_hd__nor2_2 _1528_ (.A(_0155_),
    .B(_0156_),
    .Y(net88));
 sky130_fd_sc_hd__and2_1 _1529_ (.A(_0076_),
    .B(\wRs1Data[26] ),
    .X(_0157_));
 sky130_fd_sc_hd__a211o_1 _1530_ (.A1(_0075_),
    .A2(\rWrDataWB[26] ),
    .B1(_0619_),
    .C1(_0157_),
    .X(_0158_));
 sky130_fd_sc_hd__o21ai_2 _1531_ (.A1(\rWrData[26] ),
    .A2(_0087_),
    .B1(_0158_),
    .Y(_0159_));
 sky130_fd_sc_hd__o21ai_1 _1532_ (.A1(_0154_),
    .A2(_0148_),
    .B1(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__inv_2 _1533_ (.A(_0160_),
    .Y(_0161_));
 sky130_fd_sc_hd__inv_2 _1534_ (.A(_0159_),
    .Y(_0162_));
 sky130_fd_sc_hd__nand2_1 _1535_ (.A(_0155_),
    .B(_0162_),
    .Y(_0163_));
 sky130_fd_sc_hd__nand2_1 _1536_ (.A(_0163_),
    .B(_0794_),
    .Y(_0164_));
 sky130_fd_sc_hd__nor2_1 _1537_ (.A(_0161_),
    .B(_0164_),
    .Y(net89));
 sky130_fd_sc_hd__or2_1 _1538_ (.A(\rWrDataWB[27] ),
    .B(_0938_),
    .X(_0165_));
 sky130_fd_sc_hd__o21ai_1 _1539_ (.A1(\wRs1Data[27] ),
    .A2(_0075_),
    .B1(_0165_),
    .Y(_0166_));
 sky130_fd_sc_hd__inv_2 _1540_ (.A(\rWrData[27] ),
    .Y(_0167_));
 sky130_fd_sc_hd__mux2_2 _1541_ (.A0(_0166_),
    .A1(_0167_),
    .S(_0619_),
    .X(_0168_));
 sky130_fd_sc_hd__inv_2 _1542_ (.A(_0168_),
    .Y(_0169_));
 sky130_fd_sc_hd__and4_1 _1543_ (.A(_0162_),
    .B(_0169_),
    .C(_0141_),
    .D(_0153_),
    .X(_0170_));
 sky130_fd_sc_hd__nand3_1 _1544_ (.A(_0134_),
    .B(_0065_),
    .C(_0170_),
    .Y(_0171_));
 sky130_fd_sc_hd__nand2_1 _1545_ (.A(_0171_),
    .B(_0914_),
    .Y(_0172_));
 sky130_fd_sc_hd__a21oi_1 _1546_ (.A1(_0163_),
    .A2(_0168_),
    .B1(_0172_),
    .Y(net90));
 sky130_fd_sc_hd__nand3_2 _1547_ (.A(_0064_),
    .B(_0147_),
    .C(_0170_),
    .Y(_0173_));
 sky130_fd_sc_hd__buf_2 _1548_ (.A(_0899_),
    .X(_0174_));
 sky130_fd_sc_hd__and2_1 _1549_ (.A(_0096_),
    .B(\wRs1Data[28] ),
    .X(_0175_));
 sky130_fd_sc_hd__a21o_1 _1550_ (.A1(_0121_),
    .A2(\wRegWrData[28] ),
    .B1(_0620_),
    .X(_0176_));
 sky130_fd_sc_hd__o22ai_4 _1551_ (.A1(\rWrData[28] ),
    .A2(_0174_),
    .B1(_0175_),
    .B2(_0176_),
    .Y(_0177_));
 sky130_fd_sc_hd__o21ai_1 _1552_ (.A1(_0177_),
    .A2(_0171_),
    .B1(_0816_),
    .Y(_0178_));
 sky130_fd_sc_hd__a21oi_1 _1553_ (.A1(_0173_),
    .A2(_0177_),
    .B1(_0178_),
    .Y(net91));
 sky130_fd_sc_hd__mux2_1 _1554_ (.A0(\rWrDataWB[29] ),
    .A1(\wRs1Data[29] ),
    .S(_0076_),
    .X(_0179_));
 sky130_fd_sc_hd__nand2_1 _1555_ (.A(_0620_),
    .B(\rWrData[29] ),
    .Y(_0180_));
 sky130_fd_sc_hd__a21bo_1 _1556_ (.A1(_0179_),
    .A2(_0174_),
    .B1_N(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__inv_2 _1557_ (.A(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__or2_1 _1558_ (.A(_0177_),
    .B(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__o21ai_1 _1559_ (.A1(_0183_),
    .A2(_0171_),
    .B1(_0816_),
    .Y(_0184_));
 sky130_fd_sc_hd__o21a_1 _1560_ (.A1(_0177_),
    .A2(_0173_),
    .B1(_0182_),
    .X(_0185_));
 sky130_fd_sc_hd__nor2_2 _1561_ (.A(_0184_),
    .B(_0185_),
    .Y(net92));
 sky130_fd_sc_hd__and2_1 _1562_ (.A(_0096_),
    .B(\wRs1Data[30] ),
    .X(_0186_));
 sky130_fd_sc_hd__a211o_1 _1563_ (.A1(_0121_),
    .A2(\rWrDataWB[30] ),
    .B1(_0620_),
    .C1(_0186_),
    .X(_0187_));
 sky130_fd_sc_hd__o21a_2 _1564_ (.A1(\rWrData[30] ),
    .A2(_0174_),
    .B1(_0187_),
    .X(_0188_));
 sky130_fd_sc_hd__nor2_1 _1565_ (.A(_0183_),
    .B(_0173_),
    .Y(_0189_));
 sky130_fd_sc_hd__nor2_1 _1566_ (.A(_0188_),
    .B(_0189_),
    .Y(_0190_));
 sky130_fd_sc_hd__nand2_1 _1567_ (.A(_0189_),
    .B(_0188_),
    .Y(_0191_));
 sky130_fd_sc_hd__nand2_1 _1568_ (.A(_0191_),
    .B(_0816_),
    .Y(_0192_));
 sky130_fd_sc_hd__nor2_1 _1569_ (.A(_0190_),
    .B(_0192_),
    .Y(net94));
 sky130_fd_sc_hd__and2_1 _1570_ (.A(_0096_),
    .B(\wRs1Data[31] ),
    .X(_0193_));
 sky130_fd_sc_hd__a211o_1 _1571_ (.A1(_0121_),
    .A2(\rWrDataWB[31] ),
    .B1(_0620_),
    .C1(_0193_),
    .X(_0194_));
 sky130_fd_sc_hd__o21a_2 _1572_ (.A1(\rWrData[31] ),
    .A2(_0174_),
    .B1(_0194_),
    .X(_0195_));
 sky130_fd_sc_hd__inv_2 _1573_ (.A(_0188_),
    .Y(_0196_));
 sky130_fd_sc_hd__nor3_1 _1574_ (.A(_0183_),
    .B(_0196_),
    .C(_0173_),
    .Y(_0197_));
 sky130_fd_sc_hd__nor2_1 _1575_ (.A(_0195_),
    .B(_0197_),
    .Y(_0198_));
 sky130_fd_sc_hd__nand3_1 _1576_ (.A(_0189_),
    .B(_0188_),
    .C(_0195_),
    .Y(_0199_));
 sky130_fd_sc_hd__nand2_1 _1577_ (.A(_0199_),
    .B(_0816_),
    .Y(_0200_));
 sky130_fd_sc_hd__nor2_1 _1578_ (.A(_0198_),
    .B(_0200_),
    .Y(net95));
 sky130_fd_sc_hd__inv_2 _1579_ (.A(_0631_),
    .Y(_0201_));
 sky130_fd_sc_hd__clkbuf_2 _1580_ (.A(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__xor2_1 _1581_ (.A(\reg_s2[3] ),
    .B(net972),
    .X(_0203_));
 sky130_fd_sc_hd__or2_1 _1582_ (.A(\reg_s2[4] ),
    .B(\rReg_d2[4] ),
    .X(_0204_));
 sky130_fd_sc_hd__nand2_1 _1583_ (.A(\reg_s2[4] ),
    .B(\rReg_d2[4] ),
    .Y(_0205_));
 sky130_fd_sc_hd__nor2_1 _1584_ (.A(\reg_s2[2] ),
    .B(_0717_),
    .Y(_0206_));
 sky130_fd_sc_hd__a221o_1 _1585_ (.A1(_0621_),
    .A2(\rReg_d2[1] ),
    .B1(_0204_),
    .B2(_0205_),
    .C1(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__a2111oi_2 _1586_ (.A1(\reg_s2[2] ),
    .A2(_0717_),
    .B1(_0728_),
    .C1(_0203_),
    .D1(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__nor2_1 _1587_ (.A(\rReg_d2[0] ),
    .B(_0628_),
    .Y(_0209_));
 sky130_fd_sc_hd__a21o_1 _1588_ (.A1(\reg_s2[1] ),
    .A2(_0712_),
    .B1(_0209_),
    .X(_0210_));
 sky130_fd_sc_hd__a211oi_4 _1589_ (.A1(_0628_),
    .A2(\rReg_d2[0] ),
    .B1(_0726_),
    .C1(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__nand2_1 _1590_ (.A(net286),
    .B(_0211_),
    .Y(_0212_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1591_ (.A(_0212_),
    .X(_0213_));
 sky130_fd_sc_hd__and2_1 _1592_ (.A(_0213_),
    .B(\wRs2Data[0] ),
    .X(_0214_));
 sky130_fd_sc_hd__clkbuf_2 _1593_ (.A(net286),
    .X(_0215_));
 sky130_fd_sc_hd__clkbuf_2 _1594_ (.A(_0211_),
    .X(_0216_));
 sky130_fd_sc_hd__clkbuf_2 _1595_ (.A(_0631_),
    .X(_0217_));
 sky130_fd_sc_hd__a31o_1 _1596_ (.A1(_0215_),
    .A2(net319),
    .A3(_0216_),
    .B1(_0217_),
    .X(_0218_));
 sky130_fd_sc_hd__o22a_2 _1597_ (.A1(\rWrData[0] ),
    .A2(_0202_),
    .B1(_0214_),
    .B2(_0218_),
    .X(net103));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1598_ (.A(_0212_),
    .X(_0219_));
 sky130_fd_sc_hd__and2_1 _1599_ (.A(_0219_),
    .B(\wRs2Data[1] ),
    .X(_0220_));
 sky130_fd_sc_hd__buf_2 _1600_ (.A(_0212_),
    .X(_0221_));
 sky130_fd_sc_hd__clkbuf_2 _1601_ (.A(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1602_ (.A(_0201_),
    .X(_0223_));
 sky130_fd_sc_hd__o21ai_1 _1603_ (.A1(_0757_),
    .A2(_0222_),
    .B1(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__o22a_2 _1604_ (.A1(\rWrData[1] ),
    .A2(_0202_),
    .B1(_0220_),
    .B2(_0224_),
    .X(net114));
 sky130_fd_sc_hd__buf_2 _1605_ (.A(_0201_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_1 _1606_ (.A0(\rWrDataWB[2] ),
    .A1(\wRs2Data[2] ),
    .S(_0221_),
    .X(_0226_));
 sky130_fd_sc_hd__clkbuf_2 _1607_ (.A(_0201_),
    .X(_0227_));
 sky130_fd_sc_hd__nand2_1 _1608_ (.A(_0226_),
    .B(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__o21ai_4 _1609_ (.A1(_0774_),
    .A2(_0225_),
    .B1(_0228_),
    .Y(net125));
 sky130_fd_sc_hd__and2_1 _1610_ (.A(_0219_),
    .B(\wRs2Data[3] ),
    .X(_0229_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1611_ (.A(_0212_),
    .X(_0230_));
 sky130_fd_sc_hd__o21ai_1 _1612_ (.A1(_0786_),
    .A2(_0230_),
    .B1(_0223_),
    .Y(_0231_));
 sky130_fd_sc_hd__o22a_1 _1613_ (.A1(\rWrData[3] ),
    .A2(_0202_),
    .B1(_0229_),
    .B2(_0231_),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_4 _1614_ (.A(_0201_),
    .X(_0232_));
 sky130_fd_sc_hd__inv_2 _1615_ (.A(_0219_),
    .Y(_0233_));
 sky130_fd_sc_hd__buf_2 _1616_ (.A(_0631_),
    .X(_0234_));
 sky130_fd_sc_hd__nor2_1 _1617_ (.A(\wRs2Data[4] ),
    .B(_0233_),
    .Y(_0235_));
 sky130_fd_sc_hd__a211o_1 _1618_ (.A1(_0804_),
    .A2(_0233_),
    .B1(_0234_),
    .C1(_0235_),
    .X(_0236_));
 sky130_fd_sc_hd__o21ai_2 _1619_ (.A1(_0808_),
    .A2(_0232_),
    .B1(_0236_),
    .Y(net129));
 sky130_fd_sc_hd__and2_1 _1620_ (.A(_0219_),
    .B(\wRs2Data[5] ),
    .X(_0237_));
 sky130_fd_sc_hd__o21ai_1 _1621_ (.A1(_0820_),
    .A2(_0230_),
    .B1(_0223_),
    .Y(_0238_));
 sky130_fd_sc_hd__o22a_2 _1622_ (.A1(\rWrData[5] ),
    .A2(_0202_),
    .B1(_0237_),
    .B2(_0238_),
    .X(net130));
 sky130_fd_sc_hd__buf_4 _1623_ (.A(_0223_),
    .X(_0239_));
 sky130_fd_sc_hd__a31o_1 _1624_ (.A1(_0215_),
    .A2(\rWrDataWB[6] ),
    .A3(_0216_),
    .B1(_0217_),
    .X(_0240_));
 sky130_fd_sc_hd__a21o_1 _1625_ (.A1(\wRs2Data[6] ),
    .A2(_0222_),
    .B1(_0240_),
    .X(_0241_));
 sky130_fd_sc_hd__o21ai_4 _1626_ (.A1(\rWrData[6] ),
    .A2(_0239_),
    .B1(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__inv_2 _1627_ (.A(_0242_),
    .Y(net131));
 sky130_fd_sc_hd__nor2_1 _1628_ (.A(\wRs2Data[7] ),
    .B(_0233_),
    .Y(_0243_));
 sky130_fd_sc_hd__a211o_1 _1629_ (.A1(_0858_),
    .A2(_0233_),
    .B1(_0234_),
    .C1(_0243_),
    .X(_0244_));
 sky130_fd_sc_hd__o21ai_2 _1630_ (.A1(_0854_),
    .A2(_0232_),
    .B1(_0244_),
    .Y(net132));
 sky130_fd_sc_hd__and2_1 _1631_ (.A(_0219_),
    .B(\wRs2Data[8] ),
    .X(_0245_));
 sky130_fd_sc_hd__o21ai_1 _1632_ (.A1(_0884_),
    .A2(_0230_),
    .B1(_0223_),
    .Y(_0246_));
 sky130_fd_sc_hd__o22a_1 _1633_ (.A1(\rWrData[8] ),
    .A2(_0202_),
    .B1(_0245_),
    .B2(_0246_),
    .X(net133));
 sky130_fd_sc_hd__and2_1 _1634_ (.A(_0219_),
    .B(\wRs2Data[9] ),
    .X(_0247_));
 sky130_fd_sc_hd__o21ai_1 _1635_ (.A1(_0900_),
    .A2(_0230_),
    .B1(_0223_),
    .Y(_0248_));
 sky130_fd_sc_hd__o22a_1 _1636_ (.A1(\rWrData[9] ),
    .A2(_0202_),
    .B1(_0247_),
    .B2(_0248_),
    .X(net134));
 sky130_fd_sc_hd__nor2_1 _1637_ (.A(\wRs2Data[10] ),
    .B(_0233_),
    .Y(_0249_));
 sky130_fd_sc_hd__a211o_1 _1638_ (.A1(_0919_),
    .A2(_0233_),
    .B1(_0234_),
    .C1(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__o21ai_2 _1639_ (.A1(_0928_),
    .A2(_0232_),
    .B1(_0250_),
    .Y(net104));
 sky130_fd_sc_hd__mux2_1 _1640_ (.A0(\rWrDataWB[11] ),
    .A1(\wRs2Data[11] ),
    .S(_0221_),
    .X(_0251_));
 sky130_fd_sc_hd__nand2_1 _1641_ (.A(_0251_),
    .B(_0239_),
    .Y(_0252_));
 sky130_fd_sc_hd__nand2_1 _1642_ (.A(_0234_),
    .B(\rWrData[11] ),
    .Y(_0253_));
 sky130_fd_sc_hd__nand2_2 _1643_ (.A(_0252_),
    .B(_0253_),
    .Y(net105));
 sky130_fd_sc_hd__a31o_1 _1644_ (.A1(_0215_),
    .A2(\rWrDataWB[12] ),
    .A3(_0216_),
    .B1(_0217_),
    .X(_0254_));
 sky130_fd_sc_hd__a21o_1 _1645_ (.A1(\wRs2Data[12] ),
    .A2(_0222_),
    .B1(_0254_),
    .X(_0255_));
 sky130_fd_sc_hd__o21ai_4 _1646_ (.A1(\rWrData[12] ),
    .A2(_0239_),
    .B1(_0255_),
    .Y(_0256_));
 sky130_fd_sc_hd__inv_2 _1647_ (.A(_0256_),
    .Y(net106));
 sky130_fd_sc_hd__a31o_1 _1648_ (.A1(_0215_),
    .A2(\rWrDataWB[13] ),
    .A3(_0216_),
    .B1(_0217_),
    .X(_0257_));
 sky130_fd_sc_hd__a21o_1 _1649_ (.A1(\wRs2Data[13] ),
    .A2(_0222_),
    .B1(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__o21ai_4 _1650_ (.A1(\rWrData[13] ),
    .A2(_0239_),
    .B1(_0258_),
    .Y(_0259_));
 sky130_fd_sc_hd__inv_2 _1651_ (.A(_0259_),
    .Y(net107));
 sky130_fd_sc_hd__and2_1 _1652_ (.A(_0230_),
    .B(\wRs2Data[14] ),
    .X(_0260_));
 sky130_fd_sc_hd__clkbuf_2 _1653_ (.A(net286),
    .X(_0261_));
 sky130_fd_sc_hd__clkbuf_2 _1654_ (.A(_0211_),
    .X(_0262_));
 sky130_fd_sc_hd__a31o_1 _1655_ (.A1(_0261_),
    .A2(net308),
    .A3(_0262_),
    .B1(_0234_),
    .X(_0263_));
 sky130_fd_sc_hd__o22a_2 _1656_ (.A1(\rWrData[14] ),
    .A2(_0227_),
    .B1(_0260_),
    .B2(_0263_),
    .X(net108));
 sky130_fd_sc_hd__and2_1 _1657_ (.A(_0230_),
    .B(\wRs2Data[15] ),
    .X(_0264_));
 sky130_fd_sc_hd__clkbuf_2 _1658_ (.A(_0631_),
    .X(_0265_));
 sky130_fd_sc_hd__a31o_1 _1659_ (.A1(_0261_),
    .A2(net307),
    .A3(_0262_),
    .B1(_0265_),
    .X(_0266_));
 sky130_fd_sc_hd__o22a_2 _1660_ (.A1(\rWrData[15] ),
    .A2(_0227_),
    .B1(_0264_),
    .B2(_0266_),
    .X(net109));
 sky130_fd_sc_hd__mux2_1 _1661_ (.A0(\rWrDataWB[16] ),
    .A1(\wRs2Data[16] ),
    .S(_0221_),
    .X(_0267_));
 sky130_fd_sc_hd__nand2_1 _1662_ (.A(_0267_),
    .B(_0227_),
    .Y(_0268_));
 sky130_fd_sc_hd__o21ai_2 _1663_ (.A1(_0067_),
    .A2(_0232_),
    .B1(_0268_),
    .Y(net110));
 sky130_fd_sc_hd__a31o_1 _1664_ (.A1(_0215_),
    .A2(\rWrDataWB[17] ),
    .A3(_0216_),
    .B1(_0217_),
    .X(_0269_));
 sky130_fd_sc_hd__a21o_1 _1665_ (.A1(\wRs2Data[17] ),
    .A2(_0222_),
    .B1(_0269_),
    .X(_0270_));
 sky130_fd_sc_hd__o21ai_4 _1666_ (.A1(\rWrData[17] ),
    .A2(_0239_),
    .B1(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__inv_2 _1667_ (.A(_0271_),
    .Y(net111));
 sky130_fd_sc_hd__mux2_1 _1668_ (.A0(\rWrDataWB[18] ),
    .A1(\wRs2Data[18] ),
    .S(_0221_),
    .X(_0272_));
 sky130_fd_sc_hd__nand2_1 _1669_ (.A(_0272_),
    .B(_0227_),
    .Y(_0273_));
 sky130_fd_sc_hd__o21ai_4 _1670_ (.A1(_0086_),
    .A2(_0232_),
    .B1(_0273_),
    .Y(net112));
 sky130_fd_sc_hd__clkbuf_2 _1671_ (.A(_0201_),
    .X(_0274_));
 sky130_fd_sc_hd__buf_1 _1672_ (.A(_0212_),
    .X(_0275_));
 sky130_fd_sc_hd__and2_1 _1673_ (.A(_0275_),
    .B(\wRs2Data[19] ),
    .X(_0276_));
 sky130_fd_sc_hd__a31o_1 _1674_ (.A1(_0261_),
    .A2(net303),
    .A3(_0262_),
    .B1(_0265_),
    .X(_0277_));
 sky130_fd_sc_hd__o22a_2 _1675_ (.A1(\rWrData[19] ),
    .A2(_0274_),
    .B1(_0276_),
    .B2(_0277_),
    .X(net113));
 sky130_fd_sc_hd__and2_1 _1676_ (.A(_0275_),
    .B(\wRs2Data[20] ),
    .X(_0278_));
 sky130_fd_sc_hd__a31o_1 _1677_ (.A1(_0261_),
    .A2(net302),
    .A3(_0262_),
    .B1(_0265_),
    .X(_0279_));
 sky130_fd_sc_hd__o22a_2 _1678_ (.A1(\rWrData[20] ),
    .A2(_0274_),
    .B1(_0278_),
    .B2(_0279_),
    .X(net115));
 sky130_fd_sc_hd__a31o_1 _1679_ (.A1(net286),
    .A2(\rWrDataWB[21] ),
    .A3(_0211_),
    .B1(_0217_),
    .X(_0280_));
 sky130_fd_sc_hd__a21o_1 _1680_ (.A1(\wRs2Data[21] ),
    .A2(_0222_),
    .B1(_0280_),
    .X(_0281_));
 sky130_fd_sc_hd__o21ai_4 _1681_ (.A1(\rWrData[21] ),
    .A2(_0239_),
    .B1(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__inv_2 _1682_ (.A(_0282_),
    .Y(net116));
 sky130_fd_sc_hd__and2_1 _1683_ (.A(_0275_),
    .B(\wRs2Data[22] ),
    .X(_0283_));
 sky130_fd_sc_hd__a31o_1 _1684_ (.A1(_0261_),
    .A2(net300),
    .A3(_0262_),
    .B1(_0265_),
    .X(_0284_));
 sky130_fd_sc_hd__o22a_2 _1685_ (.A1(\rWrData[22] ),
    .A2(_0274_),
    .B1(_0283_),
    .B2(_0284_),
    .X(net117));
 sky130_fd_sc_hd__and2_1 _1686_ (.A(_0275_),
    .B(\wRs2Data[23] ),
    .X(_0285_));
 sky130_fd_sc_hd__a31o_1 _1687_ (.A1(_0261_),
    .A2(\wRegWrData[23] ),
    .A3(_0262_),
    .B1(_0265_),
    .X(_0286_));
 sky130_fd_sc_hd__o22a_2 _1688_ (.A1(\rWrData[23] ),
    .A2(_0274_),
    .B1(_0285_),
    .B2(_0286_),
    .X(net118));
 sky130_fd_sc_hd__and2_1 _1689_ (.A(_0275_),
    .B(\wRs2Data[24] ),
    .X(_0287_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1690_ (.A(_0208_),
    .X(_0288_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1691_ (.A(_0211_),
    .X(_0289_));
 sky130_fd_sc_hd__a31o_1 _1692_ (.A1(_0288_),
    .A2(\wRegWrData[24] ),
    .A3(_0289_),
    .B1(_0265_),
    .X(_0290_));
 sky130_fd_sc_hd__o22a_2 _1693_ (.A1(\rWrData[24] ),
    .A2(_0274_),
    .B1(_0287_),
    .B2(_0290_),
    .X(net119));
 sky130_fd_sc_hd__and2_1 _1694_ (.A(_0275_),
    .B(\wRs2Data[25] ),
    .X(_0291_));
 sky130_fd_sc_hd__clkbuf_2 _1695_ (.A(_0631_),
    .X(_0292_));
 sky130_fd_sc_hd__a31o_1 _1696_ (.A1(_0288_),
    .A2(net297),
    .A3(_0289_),
    .B1(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__o22a_2 _1697_ (.A1(\rWrData[25] ),
    .A2(_0274_),
    .B1(_0291_),
    .B2(_0293_),
    .X(net120));
 sky130_fd_sc_hd__and2_1 _1698_ (.A(_0213_),
    .B(\wRs2Data[26] ),
    .X(_0294_));
 sky130_fd_sc_hd__a31o_1 _1699_ (.A1(_0288_),
    .A2(net295),
    .A3(_0289_),
    .B1(_0292_),
    .X(_0295_));
 sky130_fd_sc_hd__o22a_2 _1700_ (.A1(\rWrData[26] ),
    .A2(_0225_),
    .B1(_0294_),
    .B2(_0295_),
    .X(net121));
 sky130_fd_sc_hd__mux2_1 _1701_ (.A0(\rWrDataWB[27] ),
    .A1(\wRs2Data[27] ),
    .S(_0221_),
    .X(_0296_));
 sky130_fd_sc_hd__nand2_1 _1702_ (.A(_0296_),
    .B(_0227_),
    .Y(_0297_));
 sky130_fd_sc_hd__o21ai_4 _1703_ (.A1(_0167_),
    .A2(_0232_),
    .B1(_0297_),
    .Y(net122));
 sky130_fd_sc_hd__and2_1 _1704_ (.A(_0213_),
    .B(\wRs2Data[28] ),
    .X(_0298_));
 sky130_fd_sc_hd__a31o_1 _1705_ (.A1(_0288_),
    .A2(\wRegWrData[28] ),
    .A3(_0289_),
    .B1(_0292_),
    .X(_0299_));
 sky130_fd_sc_hd__o22a_2 _1706_ (.A1(\rWrData[28] ),
    .A2(_0225_),
    .B1(_0298_),
    .B2(_0299_),
    .X(net123));
 sky130_fd_sc_hd__and2_1 _1707_ (.A(_0213_),
    .B(\wRs2Data[29] ),
    .X(_0300_));
 sky130_fd_sc_hd__a31o_1 _1708_ (.A1(_0288_),
    .A2(net291),
    .A3(_0289_),
    .B1(_0292_),
    .X(_0301_));
 sky130_fd_sc_hd__o22a_2 _1709_ (.A1(\rWrData[29] ),
    .A2(_0225_),
    .B1(_0300_),
    .B2(_0301_),
    .X(net124));
 sky130_fd_sc_hd__and2_1 _1710_ (.A(_0213_),
    .B(\wRs2Data[30] ),
    .X(_0302_));
 sky130_fd_sc_hd__a31o_1 _1711_ (.A1(_0288_),
    .A2(\wRegWrData[30] ),
    .A3(_0289_),
    .B1(_0292_),
    .X(_0303_));
 sky130_fd_sc_hd__o22a_2 _1712_ (.A1(\rWrData[30] ),
    .A2(_0225_),
    .B1(_0302_),
    .B2(_0303_),
    .X(net126));
 sky130_fd_sc_hd__and2_1 _1713_ (.A(_0213_),
    .B(\wRs2Data[31] ),
    .X(_0304_));
 sky130_fd_sc_hd__a31o_1 _1714_ (.A1(_0215_),
    .A2(net288),
    .A3(_0216_),
    .B1(_0292_),
    .X(_0305_));
 sky130_fd_sc_hd__o22a_2 _1715_ (.A1(\rWrData[31] ),
    .A2(_0225_),
    .B1(_0304_),
    .B2(_0305_),
    .X(net127));
 sky130_fd_sc_hd__nor2_1 _1716_ (.A(net901),
    .B(net321),
    .Y(_0306_));
 sky130_fd_sc_hd__inv_2 _1717_ (.A(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__buf_1 _1718_ (.A(_0307_),
    .X(_0308_));
 sky130_fd_sc_hd__inv_2 _1719_ (.A(net925),
    .Y(_0309_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1720_ (.A(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__and3_1 _1721_ (.A(_0308_),
    .B(\wPcReturn[0] ),
    .C(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__a21o_1 _1722_ (.A1(net1076),
    .A2(net927),
    .B1(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__nor2_2 _1723_ (.A(op_intRegImm),
    .B(op_consShf),
    .Y(_0313_));
 sky130_fd_sc_hd__or3b_1 _1724_ (.A(net907),
    .B(op_intRegReg),
    .C_N(_0313_),
    .X(_0314_));
 sky130_fd_sc_hd__clkbuf_2 _1725_ (.A(_0314_),
    .X(_0315_));
 sky130_fd_sc_hd__clkbuf_4 _1726_ (.A(_0315_),
    .X(_0316_));
 sky130_fd_sc_hd__mux2_1 _1727_ (.A0(_0312_),
    .A1(\wAluOut[0] ),
    .S(_0316_),
    .X(_0317_));
 sky130_fd_sc_hd__clkbuf_1 _1728_ (.A(_0317_),
    .X(_0002_));
 sky130_fd_sc_hd__buf_1 _1729_ (.A(_0310_),
    .X(_0318_));
 sky130_fd_sc_hd__and3_1 _1730_ (.A(_0308_),
    .B(_0318_),
    .C(\wPcReturn[1] ),
    .X(_0319_));
 sky130_fd_sc_hd__a21o_1 _1731_ (.A1(net927),
    .A2(net1078),
    .B1(_0319_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_1 _1732_ (.A0(_0320_),
    .A1(\wAluOut[1] ),
    .S(_0316_),
    .X(_0321_));
 sky130_fd_sc_hd__clkbuf_1 _1733_ (.A(_0321_),
    .X(_0013_));
 sky130_fd_sc_hd__buf_1 _1734_ (.A(_0310_),
    .X(_0322_));
 sky130_fd_sc_hd__and2_1 _1735_ (.A(_0322_),
    .B(\wPcReturn[2] ),
    .X(_0323_));
 sky130_fd_sc_hd__buf_2 _1736_ (.A(_0307_),
    .X(_0324_));
 sky130_fd_sc_hd__a22o_1 _1737_ (.A1(net923),
    .A2(net1080),
    .B1(_0323_),
    .B2(_0324_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_1 _1738_ (.A0(_0325_),
    .A1(\wAluOut[2] ),
    .S(_0316_),
    .X(_0326_));
 sky130_fd_sc_hd__clkbuf_1 _1739_ (.A(_0326_),
    .X(_0024_));
 sky130_fd_sc_hd__and3_1 _1740_ (.A(_0308_),
    .B(_0318_),
    .C(\wPcReturn[3] ),
    .X(_0327_));
 sky130_fd_sc_hd__a21o_1 _1741_ (.A1(net927),
    .A2(net1082),
    .B1(_0327_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _1742_ (.A0(_0328_),
    .A1(\wAluOut[3] ),
    .S(_0316_),
    .X(_0329_));
 sky130_fd_sc_hd__clkbuf_1 _1743_ (.A(_0329_),
    .X(_0027_));
 sky130_fd_sc_hd__and2_1 _1744_ (.A(_0322_),
    .B(\wPcReturn[4] ),
    .X(_0330_));
 sky130_fd_sc_hd__a22o_1 _1745_ (.A1(net923),
    .A2(net1084),
    .B1(_0330_),
    .B2(_0324_),
    .X(_0331_));
 sky130_fd_sc_hd__mux2_1 _1746_ (.A0(_0331_),
    .A1(\wAluOut[4] ),
    .S(_0316_),
    .X(_0332_));
 sky130_fd_sc_hd__clkbuf_1 _1747_ (.A(_0332_),
    .X(_0028_));
 sky130_fd_sc_hd__buf_1 _1748_ (.A(_0310_),
    .X(_0333_));
 sky130_fd_sc_hd__and3_1 _1749_ (.A(_0308_),
    .B(_0333_),
    .C(\wPcReturn[5] ),
    .X(_0334_));
 sky130_fd_sc_hd__a21o_1 _1750_ (.A1(net923),
    .A2(net1086),
    .B1(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__clkbuf_2 _1751_ (.A(_0315_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_1 _1752_ (.A0(_0335_),
    .A1(\wAluOut[5] ),
    .S(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__clkbuf_1 _1753_ (.A(_0337_),
    .X(_0029_));
 sky130_fd_sc_hd__and2_1 _1754_ (.A(_0322_),
    .B(\wPcReturn[6] ),
    .X(_0338_));
 sky130_fd_sc_hd__a22o_1 _1755_ (.A1(net923),
    .A2(net1088),
    .B1(_0338_),
    .B2(_0324_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_1 _1756_ (.A0(_0339_),
    .A1(\wAluOut[6] ),
    .S(_0336_),
    .X(_0340_));
 sky130_fd_sc_hd__clkbuf_1 _1757_ (.A(_0340_),
    .X(_0030_));
 sky130_fd_sc_hd__and2_1 _1758_ (.A(_0322_),
    .B(\wPcReturn[7] ),
    .X(_0341_));
 sky130_fd_sc_hd__a22o_1 _1759_ (.A1(net923),
    .A2(net1090),
    .B1(_0341_),
    .B2(_0324_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_1 _1760_ (.A0(_0342_),
    .A1(\wAluOut[7] ),
    .S(_0336_),
    .X(_0343_));
 sky130_fd_sc_hd__clkbuf_1 _1761_ (.A(_0343_),
    .X(_0031_));
 sky130_fd_sc_hd__and2_1 _1762_ (.A(_0322_),
    .B(\wPcReturn[8] ),
    .X(_0344_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1763_ (.A(_0307_),
    .X(_0345_));
 sky130_fd_sc_hd__clkbuf_2 _1764_ (.A(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__a22o_1 _1765_ (.A1(net924),
    .A2(net1092),
    .B1(_0344_),
    .B2(_0346_),
    .X(_0347_));
 sky130_fd_sc_hd__mux2_1 _1766_ (.A0(_0347_),
    .A1(\wAluOut[8] ),
    .S(_0336_),
    .X(_0348_));
 sky130_fd_sc_hd__clkbuf_1 _1767_ (.A(_0348_),
    .X(_0032_));
 sky130_fd_sc_hd__and3_1 _1768_ (.A(_0308_),
    .B(_0333_),
    .C(\wPcReturn[9] ),
    .X(_0349_));
 sky130_fd_sc_hd__a21o_1 _1769_ (.A1(net924),
    .A2(net1094),
    .B1(_0349_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _1770_ (.A0(_0350_),
    .A1(\wAluOut[9] ),
    .S(_0336_),
    .X(_0351_));
 sky130_fd_sc_hd__clkbuf_1 _1771_ (.A(_0351_),
    .X(_0033_));
 sky130_fd_sc_hd__and2_1 _1772_ (.A(_0322_),
    .B(\wPcReturn[10] ),
    .X(_0352_));
 sky130_fd_sc_hd__a22o_1 _1773_ (.A1(net923),
    .A2(net1096),
    .B1(_0352_),
    .B2(_0346_),
    .X(_0353_));
 sky130_fd_sc_hd__mux2_1 _1774_ (.A0(_0353_),
    .A1(\wAluOut[10] ),
    .S(_0336_),
    .X(_0354_));
 sky130_fd_sc_hd__clkbuf_1 _1775_ (.A(_0354_),
    .X(_0003_));
 sky130_fd_sc_hd__buf_1 _1776_ (.A(_0310_),
    .X(_0355_));
 sky130_fd_sc_hd__and2_1 _1777_ (.A(_0355_),
    .B(\wPcReturn[11] ),
    .X(_0356_));
 sky130_fd_sc_hd__a22o_1 _1778_ (.A1(net922),
    .A2(net1098),
    .B1(_0356_),
    .B2(_0346_),
    .X(_0357_));
 sky130_fd_sc_hd__clkbuf_2 _1779_ (.A(_0315_),
    .X(_0358_));
 sky130_fd_sc_hd__mux2_1 _1780_ (.A0(_0357_),
    .A1(\wAluOut[11] ),
    .S(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__clkbuf_1 _1781_ (.A(_0359_),
    .X(_0004_));
 sky130_fd_sc_hd__and2_1 _1782_ (.A(_0355_),
    .B(\wPcReturn[12] ),
    .X(_0360_));
 sky130_fd_sc_hd__a22o_1 _1783_ (.A1(net922),
    .A2(\imm32_u[12] ),
    .B1(_0360_),
    .B2(_0346_),
    .X(_0361_));
 sky130_fd_sc_hd__mux2_1 _1784_ (.A0(_0361_),
    .A1(\wAluOut[12] ),
    .S(_0358_),
    .X(_0362_));
 sky130_fd_sc_hd__clkbuf_1 _1785_ (.A(_0362_),
    .X(_0005_));
 sky130_fd_sc_hd__and3_1 _1786_ (.A(_0308_),
    .B(_0333_),
    .C(\wPcReturn[13] ),
    .X(_0363_));
 sky130_fd_sc_hd__a21o_1 _1787_ (.A1(net922),
    .A2(\imm32_u[13] ),
    .B1(_0363_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_1 _1788_ (.A0(_0364_),
    .A1(\wAluOut[13] ),
    .S(_0358_),
    .X(_0365_));
 sky130_fd_sc_hd__clkbuf_1 _1789_ (.A(_0365_),
    .X(_0006_));
 sky130_fd_sc_hd__buf_1 _1790_ (.A(_0307_),
    .X(_0366_));
 sky130_fd_sc_hd__and3_1 _1791_ (.A(_0366_),
    .B(_0333_),
    .C(\wPcReturn[14] ),
    .X(_0367_));
 sky130_fd_sc_hd__a21o_1 _1792_ (.A1(net924),
    .A2(\imm32_u[14] ),
    .B1(_0367_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_1 _1793_ (.A0(_0368_),
    .A1(\wAluOut[14] ),
    .S(_0358_),
    .X(_0369_));
 sky130_fd_sc_hd__clkbuf_1 _1794_ (.A(_0369_),
    .X(_0007_));
 sky130_fd_sc_hd__and2_1 _1795_ (.A(_0355_),
    .B(\wPcReturn[15] ),
    .X(_0370_));
 sky130_fd_sc_hd__a22o_1 _1796_ (.A1(net924),
    .A2(\imm32_u[15] ),
    .B1(_0370_),
    .B2(_0346_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_1 _1797_ (.A0(_0371_),
    .A1(\wAluOut[15] ),
    .S(_0358_),
    .X(_0372_));
 sky130_fd_sc_hd__clkbuf_1 _1798_ (.A(_0372_),
    .X(_0008_));
 sky130_fd_sc_hd__and2_1 _1799_ (.A(_0355_),
    .B(\wPcReturn[16] ),
    .X(_0373_));
 sky130_fd_sc_hd__a22o_1 _1800_ (.A1(net922),
    .A2(\imm32_u[16] ),
    .B1(_0373_),
    .B2(_0346_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_1 _1801_ (.A0(_0374_),
    .A1(\wAluOut[16] ),
    .S(_0358_),
    .X(_0375_));
 sky130_fd_sc_hd__clkbuf_1 _1802_ (.A(_0375_),
    .X(_0009_));
 sky130_fd_sc_hd__and3_1 _1803_ (.A(_0366_),
    .B(_0333_),
    .C(\wPcReturn[17] ),
    .X(_0376_));
 sky130_fd_sc_hd__a21o_1 _1804_ (.A1(net922),
    .A2(\imm32_u[17] ),
    .B1(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__clkbuf_2 _1805_ (.A(_0314_),
    .X(_0378_));
 sky130_fd_sc_hd__mux2_1 _1806_ (.A0(_0377_),
    .A1(\wAluOut[17] ),
    .S(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__clkbuf_1 _1807_ (.A(_0379_),
    .X(_0010_));
 sky130_fd_sc_hd__and3_1 _1808_ (.A(_0366_),
    .B(_0333_),
    .C(\wPcReturn[18] ),
    .X(_0380_));
 sky130_fd_sc_hd__a21o_1 _1809_ (.A1(net922),
    .A2(\imm32_u[18] ),
    .B1(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__mux2_1 _1810_ (.A0(_0381_),
    .A1(\wAluOut[18] ),
    .S(_0378_),
    .X(_0382_));
 sky130_fd_sc_hd__clkbuf_1 _1811_ (.A(_0382_),
    .X(_0011_));
 sky130_fd_sc_hd__and2_1 _1812_ (.A(_0355_),
    .B(\wPcReturn[19] ),
    .X(_0383_));
 sky130_fd_sc_hd__clkbuf_2 _1813_ (.A(_0345_),
    .X(_0384_));
 sky130_fd_sc_hd__a22o_1 _1814_ (.A1(net926),
    .A2(\imm32_u[19] ),
    .B1(_0383_),
    .B2(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _1815_ (.A0(_0385_),
    .A1(\wAluOut[19] ),
    .S(_0378_),
    .X(_0386_));
 sky130_fd_sc_hd__clkbuf_1 _1816_ (.A(_0386_),
    .X(_0012_));
 sky130_fd_sc_hd__and2_1 _1817_ (.A(_0355_),
    .B(\wPcReturn[20] ),
    .X(_0387_));
 sky130_fd_sc_hd__a22o_1 _1818_ (.A1(net926),
    .A2(\imm32_u[20] ),
    .B1(_0387_),
    .B2(_0384_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _1819_ (.A0(_0388_),
    .A1(\wAluOut[20] ),
    .S(_0378_),
    .X(_0389_));
 sky130_fd_sc_hd__clkbuf_1 _1820_ (.A(_0389_),
    .X(_0014_));
 sky130_fd_sc_hd__buf_1 _1821_ (.A(_0309_),
    .X(_0390_));
 sky130_fd_sc_hd__and3_1 _1822_ (.A(_0366_),
    .B(_0390_),
    .C(\wPcReturn[21] ),
    .X(_0391_));
 sky130_fd_sc_hd__a21o_1 _1823_ (.A1(net926),
    .A2(\imm32_u[21] ),
    .B1(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_1 _1824_ (.A0(_0392_),
    .A1(\wAluOut[21] ),
    .S(_0378_),
    .X(_0393_));
 sky130_fd_sc_hd__clkbuf_1 _1825_ (.A(_0393_),
    .X(_0015_));
 sky130_fd_sc_hd__and2_1 _1826_ (.A(_0318_),
    .B(\wPcReturn[22] ),
    .X(_0394_));
 sky130_fd_sc_hd__a22o_1 _1827_ (.A1(net926),
    .A2(\imm32_u[22] ),
    .B1(_0394_),
    .B2(_0384_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_1 _1828_ (.A0(_0395_),
    .A1(\wAluOut[22] ),
    .S(_0378_),
    .X(_0396_));
 sky130_fd_sc_hd__clkbuf_1 _1829_ (.A(_0396_),
    .X(_0016_));
 sky130_fd_sc_hd__and2_1 _1830_ (.A(_0318_),
    .B(\wPcReturn[23] ),
    .X(_0397_));
 sky130_fd_sc_hd__a22o_1 _1831_ (.A1(net928),
    .A2(\imm32_u[23] ),
    .B1(_0397_),
    .B2(_0384_),
    .X(_0398_));
 sky130_fd_sc_hd__clkbuf_2 _1832_ (.A(_0314_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_1 _1833_ (.A0(_0398_),
    .A1(\wAluOut[23] ),
    .S(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__clkbuf_1 _1834_ (.A(_0400_),
    .X(_0017_));
 sky130_fd_sc_hd__and2_1 _1835_ (.A(_0318_),
    .B(\wPcReturn[24] ),
    .X(_0401_));
 sky130_fd_sc_hd__a22o_1 _1836_ (.A1(net928),
    .A2(\imm32_u[24] ),
    .B1(_0401_),
    .B2(_0384_),
    .X(_0402_));
 sky130_fd_sc_hd__mux2_1 _1837_ (.A0(_0402_),
    .A1(\wAluOut[24] ),
    .S(_0399_),
    .X(_0403_));
 sky130_fd_sc_hd__clkbuf_1 _1838_ (.A(_0403_),
    .X(_0018_));
 sky130_fd_sc_hd__and3_1 _1839_ (.A(_0366_),
    .B(_0390_),
    .C(\wPcReturn[25] ),
    .X(_0404_));
 sky130_fd_sc_hd__a21o_1 _1840_ (.A1(net925),
    .A2(\imm32_u[25] ),
    .B1(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__mux2_1 _1841_ (.A0(_0405_),
    .A1(\wAluOut[25] ),
    .S(_0399_),
    .X(_0406_));
 sky130_fd_sc_hd__clkbuf_1 _1842_ (.A(_0406_),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _1843_ (.A(_0318_),
    .B(\wPcReturn[26] ),
    .X(_0407_));
 sky130_fd_sc_hd__a22o_1 _1844_ (.A1(net926),
    .A2(\imm32_u[26] ),
    .B1(_0407_),
    .B2(_0384_),
    .X(_0408_));
 sky130_fd_sc_hd__mux2_1 _1845_ (.A0(_0408_),
    .A1(\wAluOut[26] ),
    .S(_0399_),
    .X(_0409_));
 sky130_fd_sc_hd__clkbuf_1 _1846_ (.A(_0409_),
    .X(_0020_));
 sky130_fd_sc_hd__and3_1 _1847_ (.A(_0366_),
    .B(_0390_),
    .C(\wPcReturn[27] ),
    .X(_0410_));
 sky130_fd_sc_hd__a21o_1 _1848_ (.A1(net927),
    .A2(\imm32_u[27] ),
    .B1(_0410_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _1849_ (.A0(_0411_),
    .A1(\wAluOut[27] ),
    .S(_0399_),
    .X(_0412_));
 sky130_fd_sc_hd__buf_1 _1850_ (.A(_0412_),
    .X(_0021_));
 sky130_fd_sc_hd__and3_1 _1851_ (.A(_0345_),
    .B(_0390_),
    .C(\wPcReturn[28] ),
    .X(_0413_));
 sky130_fd_sc_hd__a21o_1 _1852_ (.A1(net925),
    .A2(\imm32_u[28] ),
    .B1(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_1 _1853_ (.A0(_0414_),
    .A1(\wAluOut[28] ),
    .S(_0399_),
    .X(_0415_));
 sky130_fd_sc_hd__buf_1 _1854_ (.A(_0415_),
    .X(_0022_));
 sky130_fd_sc_hd__and3_1 _1855_ (.A(_0345_),
    .B(_0390_),
    .C(\wPcReturn[29] ),
    .X(_0416_));
 sky130_fd_sc_hd__a21o_1 _1856_ (.A1(net925),
    .A2(\imm32_u[29] ),
    .B1(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _1857_ (.A0(_0417_),
    .A1(\wAluOut[29] ),
    .S(_0315_),
    .X(_0418_));
 sky130_fd_sc_hd__buf_1 _1858_ (.A(_0418_),
    .X(_0023_));
 sky130_fd_sc_hd__and3_1 _1859_ (.A(_0345_),
    .B(_0390_),
    .C(\wPcReturn[30] ),
    .X(_0419_));
 sky130_fd_sc_hd__a21o_1 _1860_ (.A1(net925),
    .A2(\imm32_u[30] ),
    .B1(_0419_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_1 _1861_ (.A0(_0420_),
    .A1(\wAluOut[30] ),
    .S(_0315_),
    .X(_0421_));
 sky130_fd_sc_hd__buf_1 _1862_ (.A(_0421_),
    .X(_0025_));
 sky130_fd_sc_hd__and3_1 _1863_ (.A(_0345_),
    .B(_0310_),
    .C(\wPcReturn[31] ),
    .X(_0422_));
 sky130_fd_sc_hd__a21o_1 _1864_ (.A1(net925),
    .A2(\imm32_u[31] ),
    .B1(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__mux2_1 _1865_ (.A0(_0423_),
    .A1(\wAluOut[31] ),
    .S(_0315_),
    .X(_0424_));
 sky130_fd_sc_hd__buf_1 _1866_ (.A(_0424_),
    .X(_0026_));
 sky130_fd_sc_hd__nor2_4 _1867_ (.A(net896),
    .B(r_type),
    .Y(_0425_));
 sky130_fd_sc_hd__inv_2 _1868_ (.A(_0425_),
    .Y(_0426_));
 sky130_fd_sc_hd__clkbuf_2 _1869_ (.A(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__clkbuf_2 _1870_ (.A(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__clkbuf_2 _1871_ (.A(_0426_),
    .X(_0429_));
 sky130_fd_sc_hd__inv_2 _1872_ (.A(net901),
    .Y(_0430_));
 sky130_fd_sc_hd__nand2_1 _1873_ (.A(_0313_),
    .B(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__clkbuf_2 _1874_ (.A(_0431_),
    .X(_0432_));
 sky130_fd_sc_hd__clkbuf_2 _1875_ (.A(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__nand2_1 _1876_ (.A(_0433_),
    .B(\imm12_i_s[0] ),
    .Y(_0434_));
 sky130_fd_sc_hd__nand2_2 _1877_ (.A(net918),
    .B(net1077),
    .Y(_0435_));
 sky130_fd_sc_hd__nor2_1 _1878_ (.A(_0426_),
    .B(_0431_),
    .Y(_0436_));
 sky130_fd_sc_hd__inv_2 _1879_ (.A(_0436_),
    .Y(_0437_));
 sky130_fd_sc_hd__buf_1 _1880_ (.A(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__clkbuf_2 _1881_ (.A(_0438_),
    .X(_0439_));
 sky130_fd_sc_hd__o22a_1 _1882_ (.A1(_0429_),
    .A2(_0434_),
    .B1(_0435_),
    .B2(_0439_),
    .X(_0440_));
 sky130_fd_sc_hd__a21bo_1 _1883_ (.A1(net103),
    .A2(_0428_),
    .B1_N(_0440_),
    .X(\wAluB[0] ));
 sky130_fd_sc_hd__nand2_1 _1884_ (.A(_0432_),
    .B(\imm12_i_s[1] ),
    .Y(_0441_));
 sky130_fd_sc_hd__nand2_2 _1885_ (.A(net920),
    .B(net1079),
    .Y(_0442_));
 sky130_fd_sc_hd__o22a_1 _1886_ (.A1(_0429_),
    .A2(_0441_),
    .B1(_0442_),
    .B2(_0439_),
    .X(_0443_));
 sky130_fd_sc_hd__a21bo_1 _1887_ (.A1(net114),
    .A2(_0428_),
    .B1_N(_0443_),
    .X(\wAluB[1] ));
 sky130_fd_sc_hd__clkbuf_2 _1888_ (.A(_0426_),
    .X(_0444_));
 sky130_fd_sc_hd__clkbuf_2 _1889_ (.A(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__nand2_1 _1890_ (.A(net125),
    .B(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__nand2_1 _1891_ (.A(_0433_),
    .B(\imm12_i_s[2] ),
    .Y(_0447_));
 sky130_fd_sc_hd__nand2_2 _1892_ (.A(net910),
    .B(net1081),
    .Y(_0448_));
 sky130_fd_sc_hd__clkbuf_2 _1893_ (.A(_0438_),
    .X(_0449_));
 sky130_fd_sc_hd__o22a_1 _1894_ (.A1(_0427_),
    .A2(_0447_),
    .B1(_0448_),
    .B2(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__nand2_2 _1895_ (.A(_0446_),
    .B(_0450_),
    .Y(\wAluB[2] ));
 sky130_fd_sc_hd__nand2_1 _1896_ (.A(_0432_),
    .B(\imm12_i_s[3] ),
    .Y(_0451_));
 sky130_fd_sc_hd__nand2_2 _1897_ (.A(net919),
    .B(net1083),
    .Y(_0452_));
 sky130_fd_sc_hd__o22a_1 _1898_ (.A1(_0429_),
    .A2(_0451_),
    .B1(_0452_),
    .B2(_0439_),
    .X(_0453_));
 sky130_fd_sc_hd__a21bo_1 _1899_ (.A1(net128),
    .A2(_0428_),
    .B1_N(_0453_),
    .X(\wAluB[3] ));
 sky130_fd_sc_hd__nand2_1 _1900_ (.A(net129),
    .B(_0445_),
    .Y(_0454_));
 sky130_fd_sc_hd__nand2_1 _1901_ (.A(_0433_),
    .B(\imm12_i_s[4] ),
    .Y(_0455_));
 sky130_fd_sc_hd__nand2_2 _1902_ (.A(net910),
    .B(net1085),
    .Y(_0456_));
 sky130_fd_sc_hd__o22a_1 _1903_ (.A1(_0427_),
    .A2(_0455_),
    .B1(_0456_),
    .B2(_0449_),
    .X(_0457_));
 sky130_fd_sc_hd__nand2_1 _1904_ (.A(_0454_),
    .B(_0457_),
    .Y(\wAluB[4] ));
 sky130_fd_sc_hd__nand2_1 _1905_ (.A(_0432_),
    .B(\imm12_i_s[5] ),
    .Y(_0458_));
 sky130_fd_sc_hd__nand2_2 _1906_ (.A(net913),
    .B(net1087),
    .Y(_0459_));
 sky130_fd_sc_hd__clkbuf_2 _1907_ (.A(_0437_),
    .X(_0460_));
 sky130_fd_sc_hd__o22a_1 _1908_ (.A1(_0429_),
    .A2(_0458_),
    .B1(_0459_),
    .B2(_0460_),
    .X(_0461_));
 sky130_fd_sc_hd__a21bo_2 _1909_ (.A1(net130),
    .A2(_0444_),
    .B1_N(_0461_),
    .X(\wAluB[5] ));
 sky130_fd_sc_hd__nand2_1 _1910_ (.A(_0433_),
    .B(\imm12_i_s[6] ),
    .Y(_0462_));
 sky130_fd_sc_hd__nand2_2 _1911_ (.A(net910),
    .B(net1089),
    .Y(_0463_));
 sky130_fd_sc_hd__clkbuf_2 _1912_ (.A(_0438_),
    .X(_0464_));
 sky130_fd_sc_hd__o22a_1 _1913_ (.A1(_0444_),
    .A2(_0462_),
    .B1(_0463_),
    .B2(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__o21ai_4 _1914_ (.A1(_0425_),
    .A2(_0242_),
    .B1(_0465_),
    .Y(\wAluB[6] ));
 sky130_fd_sc_hd__nand2_1 _1915_ (.A(net132),
    .B(_0445_),
    .Y(_0466_));
 sky130_fd_sc_hd__nand2_1 _1916_ (.A(_0433_),
    .B(\imm12_i_s[7] ),
    .Y(_0467_));
 sky130_fd_sc_hd__nand2_2 _1917_ (.A(net909),
    .B(net1091),
    .Y(_0468_));
 sky130_fd_sc_hd__clkbuf_2 _1918_ (.A(_0438_),
    .X(_0469_));
 sky130_fd_sc_hd__o22a_1 _1919_ (.A1(_0427_),
    .A2(_0467_),
    .B1(_0468_),
    .B2(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__nand2_2 _1920_ (.A(_0466_),
    .B(_0470_),
    .Y(\wAluB[7] ));
 sky130_fd_sc_hd__nand2_1 _1921_ (.A(_0432_),
    .B(\imm12_i_s[8] ),
    .Y(_0471_));
 sky130_fd_sc_hd__nand2_2 _1922_ (.A(net912),
    .B(net1093),
    .Y(_0472_));
 sky130_fd_sc_hd__o22a_1 _1923_ (.A1(_0429_),
    .A2(_0471_),
    .B1(_0472_),
    .B2(_0460_),
    .X(_0473_));
 sky130_fd_sc_hd__a21bo_2 _1924_ (.A1(net133),
    .A2(_0444_),
    .B1_N(_0473_),
    .X(\wAluB[8] ));
 sky130_fd_sc_hd__nand2_1 _1925_ (.A(_0432_),
    .B(\imm12_i_s[9] ),
    .Y(_0474_));
 sky130_fd_sc_hd__nand2_2 _1926_ (.A(net913),
    .B(net1095),
    .Y(_0475_));
 sky130_fd_sc_hd__o22a_1 _1927_ (.A1(_0429_),
    .A2(_0474_),
    .B1(_0475_),
    .B2(_0460_),
    .X(_0476_));
 sky130_fd_sc_hd__a21bo_2 _1928_ (.A1(net134),
    .A2(_0444_),
    .B1_N(_0476_),
    .X(\wAluB[9] ));
 sky130_fd_sc_hd__nand2_1 _1929_ (.A(net104),
    .B(_0445_),
    .Y(_0477_));
 sky130_fd_sc_hd__nand2_1 _1930_ (.A(_0433_),
    .B(\imm12_i_s[10] ),
    .Y(_0478_));
 sky130_fd_sc_hd__nand2_2 _1931_ (.A(net909),
    .B(net1097),
    .Y(_0479_));
 sky130_fd_sc_hd__o22a_1 _1932_ (.A1(_0427_),
    .A2(_0478_),
    .B1(_0479_),
    .B2(_0469_),
    .X(_0480_));
 sky130_fd_sc_hd__nand2_1 _1933_ (.A(_0477_),
    .B(_0480_),
    .Y(\wAluB[10] ));
 sky130_fd_sc_hd__nand2_1 _1934_ (.A(net105),
    .B(_0445_),
    .Y(_0481_));
 sky130_fd_sc_hd__nand2_2 _1935_ (.A(net907),
    .B(net1099),
    .Y(_0482_));
 sky130_fd_sc_hd__or3b_1 _1936_ (.A(_0944_),
    .B(_0426_),
    .C_N(_0431_),
    .X(_0483_));
 sky130_fd_sc_hd__clkbuf_2 _1937_ (.A(_0483_),
    .X(_0484_));
 sky130_fd_sc_hd__clkbuf_2 _1938_ (.A(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__o21a_1 _1939_ (.A1(_0482_),
    .A2(_0469_),
    .B1(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__nand2_1 _1940_ (.A(_0481_),
    .B(_0486_),
    .Y(\wAluB[11] ));
 sky130_fd_sc_hd__nand2_1 _1941_ (.A(net907),
    .B(\imm32_u[12] ),
    .Y(_0487_));
 sky130_fd_sc_hd__o21a_1 _1942_ (.A1(_0487_),
    .A2(_0449_),
    .B1(_0485_),
    .X(_0488_));
 sky130_fd_sc_hd__o21ai_2 _1943_ (.A1(_0425_),
    .A2(_0256_),
    .B1(_0488_),
    .Y(\wAluB[12] ));
 sky130_fd_sc_hd__nand2_1 _1944_ (.A(net907),
    .B(\imm32_u[13] ),
    .Y(_0489_));
 sky130_fd_sc_hd__o21a_1 _1945_ (.A1(_0489_),
    .A2(_0449_),
    .B1(_0485_),
    .X(_0490_));
 sky130_fd_sc_hd__o21ai_2 _1946_ (.A1(_0425_),
    .A2(_0259_),
    .B1(_0490_),
    .Y(\wAluB[13] ));
 sky130_fd_sc_hd__clkbuf_2 _1947_ (.A(_0444_),
    .X(_0491_));
 sky130_fd_sc_hd__buf_2 _1948_ (.A(_0460_),
    .X(_0492_));
 sky130_fd_sc_hd__nand2_1 _1949_ (.A(net907),
    .B(\imm32_u[14] ),
    .Y(_0493_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _1950_ (.A(_0484_),
    .X(_0494_));
 sky130_fd_sc_hd__o21ai_1 _1951_ (.A1(_0492_),
    .A2(_0493_),
    .B1(_0494_),
    .Y(_0495_));
 sky130_fd_sc_hd__a21o_1 _1952_ (.A1(net108),
    .A2(_0491_),
    .B1(_0495_),
    .X(\wAluB[14] ));
 sky130_fd_sc_hd__nand2_1 _1953_ (.A(net907),
    .B(\imm32_u[15] ),
    .Y(_0496_));
 sky130_fd_sc_hd__o21ai_1 _1954_ (.A1(_0492_),
    .A2(_0496_),
    .B1(_0494_),
    .Y(_0497_));
 sky130_fd_sc_hd__a21o_1 _1955_ (.A1(net109),
    .A2(_0491_),
    .B1(_0497_),
    .X(\wAluB[15] ));
 sky130_fd_sc_hd__nand2_1 _1956_ (.A(net110),
    .B(_0445_),
    .Y(_0498_));
 sky130_fd_sc_hd__nand2_1 _1957_ (.A(net908),
    .B(\imm32_u[16] ),
    .Y(_0499_));
 sky130_fd_sc_hd__o21a_1 _1958_ (.A1(_0499_),
    .A2(_0469_),
    .B1(_0484_),
    .X(_0500_));
 sky130_fd_sc_hd__nand2_1 _1959_ (.A(_0498_),
    .B(_0500_),
    .Y(\wAluB[16] ));
 sky130_fd_sc_hd__nand2_1 _1960_ (.A(net908),
    .B(\imm32_u[17] ),
    .Y(_0501_));
 sky130_fd_sc_hd__o21a_1 _1961_ (.A1(_0501_),
    .A2(_0449_),
    .B1(_0485_),
    .X(_0502_));
 sky130_fd_sc_hd__o21ai_2 _1962_ (.A1(_0425_),
    .A2(_0271_),
    .B1(_0502_),
    .Y(\wAluB[17] ));
 sky130_fd_sc_hd__nand2_1 _1963_ (.A(net112),
    .B(_0491_),
    .Y(_0503_));
 sky130_fd_sc_hd__nand2_1 _1964_ (.A(net911),
    .B(\imm32_u[18] ),
    .Y(_0504_));
 sky130_fd_sc_hd__o21a_1 _1965_ (.A1(_0504_),
    .A2(_0469_),
    .B1(_0484_),
    .X(_0505_));
 sky130_fd_sc_hd__nand2_2 _1966_ (.A(_0503_),
    .B(_0505_),
    .Y(\wAluB[18] ));
 sky130_fd_sc_hd__clkbuf_2 _1967_ (.A(_0460_),
    .X(_0506_));
 sky130_fd_sc_hd__nand2_1 _1968_ (.A(net917),
    .B(\imm32_u[19] ),
    .Y(_0507_));
 sky130_fd_sc_hd__o21ai_1 _1969_ (.A1(_0506_),
    .A2(_0507_),
    .B1(_0494_),
    .Y(_0508_));
 sky130_fd_sc_hd__a21o_1 _1970_ (.A1(net113),
    .A2(_0491_),
    .B1(_0508_),
    .X(\wAluB[19] ));
 sky130_fd_sc_hd__nand2_1 _1971_ (.A(net917),
    .B(\imm32_u[20] ),
    .Y(_0509_));
 sky130_fd_sc_hd__o21ai_1 _1972_ (.A1(_0506_),
    .A2(_0509_),
    .B1(_0494_),
    .Y(_0510_));
 sky130_fd_sc_hd__a21o_1 _1973_ (.A1(net115),
    .A2(_0491_),
    .B1(_0510_),
    .X(\wAluB[20] ));
 sky130_fd_sc_hd__nand2_1 _1974_ (.A(net908),
    .B(\imm32_u[21] ),
    .Y(_0511_));
 sky130_fd_sc_hd__o21a_1 _1975_ (.A1(_0511_),
    .A2(_0449_),
    .B1(_0485_),
    .X(_0512_));
 sky130_fd_sc_hd__o21ai_2 _1976_ (.A1(_0425_),
    .A2(_0282_),
    .B1(_0512_),
    .Y(\wAluB[21] ));
 sky130_fd_sc_hd__clkbuf_2 _1977_ (.A(_0427_),
    .X(_0513_));
 sky130_fd_sc_hd__nand2_1 _1978_ (.A(net917),
    .B(\imm32_u[22] ),
    .Y(_0514_));
 sky130_fd_sc_hd__o21ai_1 _1979_ (.A1(_0506_),
    .A2(_0514_),
    .B1(_0494_),
    .Y(_0515_));
 sky130_fd_sc_hd__a21o_1 _1980_ (.A1(net117),
    .A2(_0513_),
    .B1(_0515_),
    .X(\wAluB[22] ));
 sky130_fd_sc_hd__nand2_1 _1981_ (.A(net917),
    .B(\imm32_u[23] ),
    .Y(_0516_));
 sky130_fd_sc_hd__o21ai_1 _1982_ (.A1(_0506_),
    .A2(_0516_),
    .B1(_0494_),
    .Y(_0517_));
 sky130_fd_sc_hd__a21o_1 _1983_ (.A1(net118),
    .A2(_0513_),
    .B1(_0517_),
    .X(\wAluB[23] ));
 sky130_fd_sc_hd__nand2_1 _1984_ (.A(net915),
    .B(\imm32_u[24] ),
    .Y(_0518_));
 sky130_fd_sc_hd__buf_1 _1985_ (.A(_0484_),
    .X(_0519_));
 sky130_fd_sc_hd__o21ai_1 _1986_ (.A1(_0506_),
    .A2(_0518_),
    .B1(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__a21o_1 _1987_ (.A1(net119),
    .A2(_0513_),
    .B1(_0520_),
    .X(\wAluB[24] ));
 sky130_fd_sc_hd__nand2_1 _1988_ (.A(net916),
    .B(\imm32_u[25] ),
    .Y(_0521_));
 sky130_fd_sc_hd__o21ai_1 _1989_ (.A1(_0506_),
    .A2(_0521_),
    .B1(_0519_),
    .Y(_0522_));
 sky130_fd_sc_hd__a21o_1 _1990_ (.A1(net120),
    .A2(_0513_),
    .B1(_0522_),
    .X(\wAluB[25] ));
 sky130_fd_sc_hd__nand2_1 _1991_ (.A(net915),
    .B(\imm32_u[26] ),
    .Y(_0523_));
 sky130_fd_sc_hd__o21ai_1 _1992_ (.A1(_0464_),
    .A2(_0523_),
    .B1(_0519_),
    .Y(_0524_));
 sky130_fd_sc_hd__a21o_1 _1993_ (.A1(net121),
    .A2(_0513_),
    .B1(_0524_),
    .X(\wAluB[26] ));
 sky130_fd_sc_hd__nand2_1 _1994_ (.A(net122),
    .B(_0491_),
    .Y(_0525_));
 sky130_fd_sc_hd__nand2_1 _1995_ (.A(net919),
    .B(\imm32_u[27] ),
    .Y(_0526_));
 sky130_fd_sc_hd__o21a_1 _1996_ (.A1(_0526_),
    .A2(_0469_),
    .B1(_0484_),
    .X(_0527_));
 sky130_fd_sc_hd__nand2_2 _1997_ (.A(_0525_),
    .B(_0527_),
    .Y(\wAluB[27] ));
 sky130_fd_sc_hd__nand2_1 _1998_ (.A(net916),
    .B(\imm32_u[28] ),
    .Y(_0528_));
 sky130_fd_sc_hd__o21ai_1 _1999_ (.A1(_0464_),
    .A2(_0528_),
    .B1(_0519_),
    .Y(_0529_));
 sky130_fd_sc_hd__a21o_2 _2000_ (.A1(net123),
    .A2(_0513_),
    .B1(_0529_),
    .X(\wAluB[28] ));
 sky130_fd_sc_hd__nand2_1 _2001_ (.A(net915),
    .B(\imm32_u[29] ),
    .Y(_0530_));
 sky130_fd_sc_hd__o21ai_1 _2002_ (.A1(_0464_),
    .A2(_0530_),
    .B1(_0519_),
    .Y(_0531_));
 sky130_fd_sc_hd__a21o_2 _2003_ (.A1(net124),
    .A2(_0428_),
    .B1(_0531_),
    .X(\wAluB[29] ));
 sky130_fd_sc_hd__nand2_1 _2004_ (.A(net915),
    .B(\imm32_u[30] ),
    .Y(_0532_));
 sky130_fd_sc_hd__o21ai_1 _2005_ (.A1(_0464_),
    .A2(_0532_),
    .B1(_0519_),
    .Y(_0533_));
 sky130_fd_sc_hd__a21o_2 _2006_ (.A1(net126),
    .A2(_0428_),
    .B1(_0533_),
    .X(\wAluB[30] ));
 sky130_fd_sc_hd__nand2_1 _2007_ (.A(net917),
    .B(\imm32_u[31] ),
    .Y(_0534_));
 sky130_fd_sc_hd__o21ai_1 _2008_ (.A1(_0464_),
    .A2(_0534_),
    .B1(_0485_),
    .Y(_0535_));
 sky130_fd_sc_hd__a21o_2 _2009_ (.A1(net127),
    .A2(_0428_),
    .B1(_0535_),
    .X(\wAluB[31] ));
 sky130_fd_sc_hd__buf_2 _2010_ (.A(_0439_),
    .X(_0536_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2011_ (.A(_0436_),
    .X(_0537_));
 sky130_fd_sc_hd__and3_1 _2012_ (.A(_0537_),
    .B(net918),
    .C(net135),
    .X(_0538_));
 sky130_fd_sc_hd__a31o_4 _2013_ (.A1(_0746_),
    .A2(_0748_),
    .A3(_0536_),
    .B1(_0538_),
    .X(\wAluA[0] ));
 sky130_fd_sc_hd__buf_2 _2014_ (.A(_0436_),
    .X(_0539_));
 sky130_fd_sc_hd__a21o_1 _2015_ (.A1(_0759_),
    .A2(_0761_),
    .B1(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__or3b_1 _2016_ (.A(_0664_),
    .B(_0438_),
    .C_N(net146),
    .X(_0541_));
 sky130_fd_sc_hd__nand2_2 _2017_ (.A(_0540_),
    .B(_0541_),
    .Y(\wAluA[1] ));
 sky130_fd_sc_hd__and3_1 _2018_ (.A(_0537_),
    .B(net911),
    .C(net379),
    .X(_0542_));
 sky130_fd_sc_hd__a31o_2 _2019_ (.A1(_0773_),
    .A2(_0775_),
    .A3(_0536_),
    .B1(_0542_),
    .X(\wAluA[2] ));
 sky130_fd_sc_hd__clkbuf_2 _2020_ (.A(_0439_),
    .X(_0543_));
 sky130_fd_sc_hd__and3_1 _2021_ (.A(_0539_),
    .B(net919),
    .C(net377),
    .X(_0544_));
 sky130_fd_sc_hd__a21o_2 _2022_ (.A1(_0790_),
    .A2(_0543_),
    .B1(_0544_),
    .X(\wAluA[3] ));
 sky130_fd_sc_hd__and3_1 _2023_ (.A(_0537_),
    .B(net910),
    .C(net376),
    .X(_0545_));
 sky130_fd_sc_hd__a31o_4 _2024_ (.A1(_0807_),
    .A2(_0809_),
    .A3(_0536_),
    .B1(_0545_),
    .X(\wAluA[4] ));
 sky130_fd_sc_hd__a21o_1 _2025_ (.A1(_0823_),
    .A2(_0824_),
    .B1(_0539_),
    .X(_0546_));
 sky130_fd_sc_hd__or3b_2 _2026_ (.A(_0664_),
    .B(_0438_),
    .C_N(net375),
    .X(_0547_));
 sky130_fd_sc_hd__nand2_4 _2027_ (.A(_0546_),
    .B(_0547_),
    .Y(\wAluA[5] ));
 sky130_fd_sc_hd__and3_1 _2028_ (.A(_0537_),
    .B(net909),
    .C(net374),
    .X(_0548_));
 sky130_fd_sc_hd__a31o_4 _2029_ (.A1(_0843_),
    .A2(_0844_),
    .A3(_0492_),
    .B1(_0548_),
    .X(\wAluA[6] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 _2030_ (.A(_0436_),
    .X(_0549_));
 sky130_fd_sc_hd__buf_1 _2031_ (.A(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__and3_1 _2032_ (.A(_0550_),
    .B(net911),
    .C(net372),
    .X(_0551_));
 sky130_fd_sc_hd__a21o_1 _2033_ (.A1(_0861_),
    .A2(_0543_),
    .B1(_0551_),
    .X(\wAluA[7] ));
 sky130_fd_sc_hd__and3_1 _2034_ (.A(_0550_),
    .B(net912),
    .C(net371),
    .X(_0552_));
 sky130_fd_sc_hd__a21o_2 _2035_ (.A1(_0891_),
    .A2(_0543_),
    .B1(_0552_),
    .X(\wAluA[8] ));
 sky130_fd_sc_hd__or2_1 _2036_ (.A(\rWrData[9] ),
    .B(_0174_),
    .X(_0553_));
 sky130_fd_sc_hd__and3_1 _2037_ (.A(_0549_),
    .B(net909),
    .C(net370),
    .X(_0554_));
 sky130_fd_sc_hd__a31o_4 _2038_ (.A1(_0904_),
    .A2(_0553_),
    .A3(_0492_),
    .B1(_0554_),
    .X(\wAluA[9] ));
 sky130_fd_sc_hd__and3_1 _2039_ (.A(_0549_),
    .B(net909),
    .C(net369),
    .X(_0555_));
 sky130_fd_sc_hd__a31o_2 _2040_ (.A1(_0927_),
    .A2(_0929_),
    .A3(_0492_),
    .B1(_0555_),
    .X(\wAluA[10] ));
 sky130_fd_sc_hd__or2_1 _2041_ (.A(\rWrData[11] ),
    .B(_0174_),
    .X(_0556_));
 sky130_fd_sc_hd__and3_1 _2042_ (.A(_0549_),
    .B(net909),
    .C(net367),
    .X(_0557_));
 sky130_fd_sc_hd__a31o_1 _2043_ (.A1(_0940_),
    .A2(_0556_),
    .A3(_0492_),
    .B1(_0557_),
    .X(\wAluA[11] ));
 sky130_fd_sc_hd__and3_1 _2044_ (.A(_0550_),
    .B(net911),
    .C(net365),
    .X(_0558_));
 sky130_fd_sc_hd__a21o_2 _2045_ (.A1(_0957_),
    .A2(_0543_),
    .B1(_0558_),
    .X(\wAluA[12] ));
 sky130_fd_sc_hd__buf_4 _2046_ (.A(_0549_),
    .X(_0559_));
 sky130_fd_sc_hd__or3b_2 _2047_ (.A(_0671_),
    .B(_0460_),
    .C_N(net139),
    .X(_0560_));
 sky130_fd_sc_hd__o21ai_4 _2048_ (.A1(_0559_),
    .A2(_0042_),
    .B1(_0560_),
    .Y(\wAluA[13] ));
 sky130_fd_sc_hd__buf_1 _2049_ (.A(_0437_),
    .X(_0561_));
 sky130_fd_sc_hd__or3b_2 _2050_ (.A(_0671_),
    .B(_0561_),
    .C_N(net361),
    .X(_0562_));
 sky130_fd_sc_hd__o21ai_4 _2051_ (.A1(_0559_),
    .A2(_0050_),
    .B1(_0562_),
    .Y(\wAluA[14] ));
 sky130_fd_sc_hd__or3b_2 _2052_ (.A(_0671_),
    .B(_0561_),
    .C_N(net359),
    .X(_0563_));
 sky130_fd_sc_hd__o21ai_4 _2053_ (.A1(_0559_),
    .A2(_0056_),
    .B1(_0563_),
    .Y(\wAluA[15] ));
 sky130_fd_sc_hd__and3_1 _2054_ (.A(_0550_),
    .B(net911),
    .C(net356),
    .X(_0564_));
 sky130_fd_sc_hd__a21o_1 _2055_ (.A1(_0071_),
    .A2(_0543_),
    .B1(_0564_),
    .X(\wAluA[16] ));
 sky130_fd_sc_hd__and3_1 _2056_ (.A(_0550_),
    .B(net911),
    .C(net353),
    .X(_0565_));
 sky130_fd_sc_hd__a21o_1 _2057_ (.A1(_0081_),
    .A2(_0543_),
    .B1(_0565_),
    .X(\wAluA[17] ));
 sky130_fd_sc_hd__nor2_1 _2058_ (.A(_0539_),
    .B(_0091_),
    .Y(_0566_));
 sky130_fd_sc_hd__a31o_2 _2059_ (.A1(net920),
    .A2(net144),
    .A3(_0539_),
    .B1(_0566_),
    .X(\wAluA[18] ));
 sky130_fd_sc_hd__clkbuf_2 _2060_ (.A(_0439_),
    .X(_0567_));
 sky130_fd_sc_hd__and3_1 _2061_ (.A(_0550_),
    .B(net919),
    .C(net349),
    .X(_0568_));
 sky130_fd_sc_hd__a21o_2 _2062_ (.A1(_0102_),
    .A2(_0567_),
    .B1(_0568_),
    .X(\wAluA[19] ));
 sky130_fd_sc_hd__or3b_1 _2063_ (.A(_0671_),
    .B(_0561_),
    .C_N(net147),
    .X(_0569_));
 sky130_fd_sc_hd__o21ai_4 _2064_ (.A1(_0559_),
    .A2(_0110_),
    .B1(_0569_),
    .Y(\wAluA[20] ));
 sky130_fd_sc_hd__or3b_1 _2065_ (.A(_0664_),
    .B(_0561_),
    .C_N(net345),
    .X(_0570_));
 sky130_fd_sc_hd__o21ai_4 _2066_ (.A1(_0559_),
    .A2(_0116_),
    .B1(_0570_),
    .Y(\wAluA[21] ));
 sky130_fd_sc_hd__or3b_1 _2067_ (.A(_0664_),
    .B(_0561_),
    .C_N(net344),
    .X(_0571_));
 sky130_fd_sc_hd__o21ai_2 _2068_ (.A1(_0559_),
    .A2(_0124_),
    .B1(_0571_),
    .Y(\wAluA[22] ));
 sky130_fd_sc_hd__buf_1 _2069_ (.A(_0549_),
    .X(_0572_));
 sky130_fd_sc_hd__and3_1 _2070_ (.A(_0572_),
    .B(net918),
    .C(net342),
    .X(_0573_));
 sky130_fd_sc_hd__a21o_2 _2071_ (.A1(_0131_),
    .A2(_0567_),
    .B1(_0573_),
    .X(\wAluA[23] ));
 sky130_fd_sc_hd__and3_1 _2072_ (.A(_0572_),
    .B(net915),
    .C(net341),
    .X(_0574_));
 sky130_fd_sc_hd__a21o_2 _2073_ (.A1(_0141_),
    .A2(_0567_),
    .B1(_0574_),
    .X(\wAluA[24] ));
 sky130_fd_sc_hd__and3_1 _2074_ (.A(_0572_),
    .B(net915),
    .C(net152),
    .X(_0575_));
 sky130_fd_sc_hd__a21o_2 _2075_ (.A1(_0153_),
    .A2(_0567_),
    .B1(_0575_),
    .X(\wAluA[25] ));
 sky130_fd_sc_hd__and3_1 _2076_ (.A(_0572_),
    .B(net916),
    .C(net338),
    .X(_0576_));
 sky130_fd_sc_hd__a21o_2 _2077_ (.A1(_0162_),
    .A2(_0567_),
    .B1(_0576_),
    .X(\wAluA[26] ));
 sky130_fd_sc_hd__and3_1 _2078_ (.A(_0572_),
    .B(net916),
    .C(net154),
    .X(_0577_));
 sky130_fd_sc_hd__a21o_2 _2079_ (.A1(_0169_),
    .A2(_0567_),
    .B1(_0577_),
    .X(\wAluA[27] ));
 sky130_fd_sc_hd__or3b_1 _2080_ (.A(_0664_),
    .B(_0561_),
    .C_N(net155),
    .X(_0578_));
 sky130_fd_sc_hd__o21ai_4 _2081_ (.A1(_0539_),
    .A2(_0177_),
    .B1(_0578_),
    .Y(\wAluA[28] ));
 sky130_fd_sc_hd__and3_1 _2082_ (.A(_0572_),
    .B(net918),
    .C(net332),
    .X(_0579_));
 sky130_fd_sc_hd__a21o_2 _2083_ (.A1(_0181_),
    .A2(_0536_),
    .B1(_0579_),
    .X(\wAluA[29] ));
 sky130_fd_sc_hd__and3_1 _2084_ (.A(_0537_),
    .B(net918),
    .C(net331),
    .X(_0580_));
 sky130_fd_sc_hd__a21o_2 _2085_ (.A1(_0188_),
    .A2(_0536_),
    .B1(_0580_),
    .X(\wAluA[30] ));
 sky130_fd_sc_hd__and3_1 _2086_ (.A(_0537_),
    .B(net918),
    .C(net159),
    .X(_0581_));
 sky130_fd_sc_hd__a21o_2 _2087_ (.A1(_0195_),
    .A2(_0536_),
    .B1(_0581_),
    .X(\wAluA[31] ));
 sky130_fd_sc_hd__or3_1 _2088_ (.A(_0593_),
    .B(_0653_),
    .C(_0661_),
    .X(_0582_));
 sky130_fd_sc_hd__buf_1 _2089_ (.A(_0582_),
    .X(wAluSextEn));
 sky130_fd_sc_hd__or2_1 _2090_ (.A(rStall2),
    .B(wStall1),
    .X(_0583_));
 sky130_fd_sc_hd__clkbuf_1 _2091_ (.A(_0583_),
    .X(wStall));
 sky130_fd_sc_hd__and2_1 _2092_ (.A(net269),
    .B(_0620_),
    .X(_0584_));
 sky130_fd_sc_hd__clkbuf_1 _2093_ (.A(_0584_),
    .X(_0000_));
 sky130_fd_sc_hd__and2_1 _2094_ (.A(net269),
    .B(_0234_),
    .X(_0585_));
 sky130_fd_sc_hd__clkbuf_1 _2095_ (.A(_0585_),
    .X(_0001_));
 sky130_fd_sc_hd__nand2_1 _2096_ (.A(_0660_),
    .B(net896),
    .Y(_0586_));
 sky130_fd_sc_hd__o21a_1 _2097_ (.A1(net896),
    .A2(_0324_),
    .B1(net1073),
    .X(_0587_));
 sky130_fd_sc_hd__nand2_1 _2098_ (.A(_0586_),
    .B(_0587_),
    .Y(_0588_));
 sky130_fd_sc_hd__inv_2 _2099_ (.A(_0588_),
    .Y(wJmp));
 sky130_fd_sc_hd__nor2_1 _2100_ (.A(net961),
    .B(rJumping2),
    .Y(_0589_));
 sky130_fd_sc_hd__nand2_1 _2101_ (.A(_0588_),
    .B(_0589_),
    .Y(wJumping));
 sky130_fd_sc_hd__nand2_1 _2102_ (.A(op_memSt),
    .B(net1019),
    .Y(_0590_));
 sky130_fd_sc_hd__inv_2 _2103_ (.A(_0590_),
    .Y(net168));
 sky130_fd_sc_hd__nand2_1 _2104_ (.A(op_memLd),
    .B(net1027),
    .Y(_0591_));
 sky130_fd_sc_hd__inv_2 _2105_ (.A(_0591_),
    .Y(net167));
 sky130_fd_sc_hd__o41a_1 _2106_ (.A1(op_memLd),
    .A2(net928),
    .A3(_0324_),
    .A4(_0316_),
    .B1(net1029),
    .X(_0034_));
 sky130_fd_sc_hd__dfxtp_1 _2107_ (.CLK(clknet_leaf_60_clk),
    .D(net1201),
    .Q(rOp_memLd));
 sky130_fd_sc_hd__dfxtp_1 _2108_ (.CLK(clknet_leaf_60_clk),
    .D(net1114),
    .Q(rOp_memLd2));
 sky130_fd_sc_hd__dfxtp_2 _2109_ (.CLK(clknet_leaf_65_clk),
    .D(net1185),
    .Q(rRegWrEn2));
 sky130_fd_sc_hd__dfxtp_1 _2110_ (.CLK(clknet_leaf_92_clk),
    .D(_0002_),
    .Q(\rWrData[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2111_ (.CLK(clknet_4_7__leaf_clk),
    .D(_0013_),
    .Q(\rWrData[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2112_ (.CLK(clknet_leaf_90_clk),
    .D(_0024_),
    .Q(\rWrData[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2113_ (.CLK(clknet_leaf_91_clk),
    .D(_0027_),
    .Q(\rWrData[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2114_ (.CLK(clknet_leaf_90_clk),
    .D(_0028_),
    .Q(\rWrData[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2115_ (.CLK(clknet_leaf_90_clk),
    .D(_0029_),
    .Q(\rWrData[5] ));
 sky130_fd_sc_hd__dfxtp_2 _2116_ (.CLK(clknet_leaf_88_clk),
    .D(_0030_),
    .Q(\rWrData[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2117_ (.CLK(clknet_leaf_90_clk),
    .D(_0031_),
    .Q(\rWrData[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2118_ (.CLK(clknet_leaf_89_clk),
    .D(_0032_),
    .Q(\rWrData[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2119_ (.CLK(clknet_leaf_90_clk),
    .D(_0033_),
    .Q(\rWrData[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2120_ (.CLK(clknet_leaf_85_clk),
    .D(_0003_),
    .Q(\rWrData[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2121_ (.CLK(clknet_leaf_88_clk),
    .D(_0004_),
    .Q(\rWrData[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2122_ (.CLK(clknet_leaf_87_clk),
    .D(_0005_),
    .Q(\rWrData[12] ));
 sky130_fd_sc_hd__dfxtp_2 _2123_ (.CLK(clknet_leaf_87_clk),
    .D(_0006_),
    .Q(\rWrData[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2124_ (.CLK(clknet_leaf_88_clk),
    .D(_0007_),
    .Q(\rWrData[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2125_ (.CLK(clknet_leaf_88_clk),
    .D(_0008_),
    .Q(\rWrData[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2126_ (.CLK(clknet_leaf_86_clk),
    .D(_0009_),
    .Q(\rWrData[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2127_ (.CLK(clknet_leaf_91_clk),
    .D(_0010_),
    .Q(\rWrData[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2128_ (.CLK(clknet_leaf_87_clk),
    .D(_0011_),
    .Q(\rWrData[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2129_ (.CLK(clknet_leaf_59_clk),
    .D(_0012_),
    .Q(\rWrData[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2130_ (.CLK(clknet_leaf_91_clk),
    .D(_0014_),
    .Q(\rWrData[20] ));
 sky130_fd_sc_hd__dfxtp_2 _2131_ (.CLK(clknet_leaf_59_clk),
    .D(_0015_),
    .Q(\rWrData[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2132_ (.CLK(clknet_leaf_55_clk),
    .D(_0016_),
    .Q(\rWrData[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2133_ (.CLK(clknet_leaf_58_clk),
    .D(_0017_),
    .Q(\rWrData[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2134_ (.CLK(clknet_leaf_59_clk),
    .D(_0018_),
    .Q(\rWrData[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2135_ (.CLK(clknet_leaf_92_clk),
    .D(_0019_),
    .Q(\rWrData[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2136_ (.CLK(clknet_leaf_55_clk),
    .D(_0020_),
    .Q(\rWrData[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2137_ (.CLK(clknet_leaf_59_clk),
    .D(_0021_),
    .Q(\rWrData[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2138_ (.CLK(clknet_leaf_59_clk),
    .D(_0022_),
    .Q(\rWrData[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2139_ (.CLK(clknet_leaf_59_clk),
    .D(_0023_),
    .Q(\rWrData[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2140_ (.CLK(clknet_leaf_59_clk),
    .D(_0025_),
    .Q(\rWrData[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2141_ (.CLK(clknet_leaf_59_clk),
    .D(_0026_),
    .Q(\rWrData[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2142_ (.CLK(clknet_leaf_86_clk),
    .D(net1161),
    .Q(\rWrDataWB[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2143_ (.CLK(clknet_leaf_79_clk),
    .D(net1100),
    .Q(\rWrDataWB[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2144_ (.CLK(clknet_leaf_84_clk),
    .D(net1155),
    .Q(\rWrDataWB[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2145_ (.CLK(clknet_leaf_86_clk),
    .D(net1158),
    .Q(\rWrDataWB[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2146_ (.CLK(clknet_leaf_84_clk),
    .D(net1169),
    .Q(\rWrDataWB[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2147_ (.CLK(clknet_leaf_84_clk),
    .D(net1175),
    .Q(\rWrDataWB[5] ));
 sky130_fd_sc_hd__dfxtp_1 _2148_ (.CLK(clknet_leaf_84_clk),
    .D(net1192),
    .Q(\rWrDataWB[6] ));
 sky130_fd_sc_hd__dfxtp_1 _2149_ (.CLK(clknet_4_13__leaf_clk),
    .D(\rWrData[7] ),
    .Q(\rWrDataWB[7] ));
 sky130_fd_sc_hd__dfxtp_1 _2150_ (.CLK(clknet_leaf_80_clk),
    .D(net1164),
    .Q(\rWrDataWB[8] ));
 sky130_fd_sc_hd__dfxtp_1 _2151_ (.CLK(clknet_leaf_84_clk),
    .D(net1214),
    .Q(\rWrDataWB[9] ));
 sky130_fd_sc_hd__dfxtp_1 _2152_ (.CLK(clknet_leaf_84_clk),
    .D(net1163),
    .Q(\rWrDataWB[10] ));
 sky130_fd_sc_hd__dfxtp_1 _2153_ (.CLK(clknet_leaf_85_clk),
    .D(net1179),
    .Q(\rWrDataWB[11] ));
 sky130_fd_sc_hd__dfxtp_1 _2154_ (.CLK(clknet_leaf_79_clk),
    .D(net1187),
    .Q(\rWrDataWB[12] ));
 sky130_fd_sc_hd__dfxtp_1 _2155_ (.CLK(clknet_leaf_86_clk),
    .D(net1166),
    .Q(\rWrDataWB[13] ));
 sky130_fd_sc_hd__dfxtp_1 _2156_ (.CLK(clknet_leaf_85_clk),
    .D(net1150),
    .Q(\rWrDataWB[14] ));
 sky130_fd_sc_hd__dfxtp_1 _2157_ (.CLK(clknet_leaf_84_clk),
    .D(net1225),
    .Q(\rWrDataWB[15] ));
 sky130_fd_sc_hd__dfxtp_1 _2158_ (.CLK(clknet_leaf_85_clk),
    .D(net1137),
    .Q(\rWrDataWB[16] ));
 sky130_fd_sc_hd__dfxtp_1 _2159_ (.CLK(clknet_leaf_86_clk),
    .D(net1190),
    .Q(\rWrDataWB[17] ));
 sky130_fd_sc_hd__dfxtp_1 _2160_ (.CLK(clknet_leaf_86_clk),
    .D(net1136),
    .Q(\rWrDataWB[18] ));
 sky130_fd_sc_hd__dfxtp_1 _2161_ (.CLK(clknet_leaf_87_clk),
    .D(net1156),
    .Q(\rWrDataWB[19] ));
 sky130_fd_sc_hd__dfxtp_1 _2162_ (.CLK(clknet_leaf_86_clk),
    .D(net1188),
    .Q(\rWrDataWB[20] ));
 sky130_fd_sc_hd__dfxtp_1 _2163_ (.CLK(clknet_leaf_87_clk),
    .D(net1181),
    .Q(\rWrDataWB[21] ));
 sky130_fd_sc_hd__dfxtp_1 _2164_ (.CLK(clknet_leaf_59_clk),
    .D(net1177),
    .Q(\rWrDataWB[22] ));
 sky130_fd_sc_hd__dfxtp_1 _2165_ (.CLK(clknet_leaf_87_clk),
    .D(net1154),
    .Q(\rWrDataWB[23] ));
 sky130_fd_sc_hd__dfxtp_1 _2166_ (.CLK(clknet_leaf_59_clk),
    .D(net1146),
    .Q(\rWrDataWB[24] ));
 sky130_fd_sc_hd__dfxtp_1 _2167_ (.CLK(clknet_leaf_59_clk),
    .D(net1159),
    .Q(\rWrDataWB[25] ));
 sky130_fd_sc_hd__dfxtp_1 _2168_ (.CLK(clknet_leaf_87_clk),
    .D(net1186),
    .Q(\rWrDataWB[26] ));
 sky130_fd_sc_hd__dfxtp_1 _2169_ (.CLK(clknet_leaf_87_clk),
    .D(net1133),
    .Q(\rWrDataWB[27] ));
 sky130_fd_sc_hd__dfxtp_1 _2170_ (.CLK(clknet_leaf_60_clk),
    .D(net1176),
    .Q(\rWrDataWB[28] ));
 sky130_fd_sc_hd__dfxtp_1 _2171_ (.CLK(clknet_leaf_59_clk),
    .D(net1145),
    .Q(\rWrDataWB[29] ));
 sky130_fd_sc_hd__dfxtp_1 _2172_ (.CLK(clknet_leaf_59_clk),
    .D(net1140),
    .Q(\rWrDataWB[30] ));
 sky130_fd_sc_hd__dfxtp_1 _2173_ (.CLK(clknet_leaf_59_clk),
    .D(net1142),
    .Q(\rWrDataWB[31] ));
 sky130_fd_sc_hd__dfxtp_1 _2174_ (.CLK(clknet_leaf_64_clk),
    .D(\reg_d[0] ),
    .Q(\rReg_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2175_ (.CLK(clknet_leaf_64_clk),
    .D(\reg_d[1] ),
    .Q(\rReg_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2176_ (.CLK(clknet_leaf_64_clk),
    .D(\reg_d[2] ),
    .Q(\rReg_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2177_ (.CLK(clknet_leaf_63_clk),
    .D(\reg_d[3] ),
    .Q(\rReg_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2178_ (.CLK(clknet_leaf_63_clk),
    .D(\reg_d[4] ),
    .Q(\rReg_d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2179_ (.CLK(clknet_leaf_65_clk),
    .D(net1971),
    .Q(\rReg_d2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _2180_ (.CLK(clknet_leaf_65_clk),
    .D(net1853),
    .Q(\rReg_d2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _2181_ (.CLK(clknet_leaf_65_clk),
    .D(net1722),
    .Q(\rReg_d2[2] ));
 sky130_fd_sc_hd__dfxtp_1 _2182_ (.CLK(clknet_leaf_64_clk),
    .D(net1165),
    .Q(\rReg_d2[3] ));
 sky130_fd_sc_hd__dfxtp_1 _2183_ (.CLK(clknet_leaf_63_clk),
    .D(net1167),
    .Q(\rReg_d2[4] ));
 sky130_fd_sc_hd__dfxtp_1 _2184_ (.CLK(clknet_leaf_62_clk),
    .D(wJmp),
    .Q(rJumping1));
 sky130_fd_sc_hd__dfxtp_1 _2185_ (.CLK(clknet_leaf_45_clk),
    .D(net961),
    .Q(rJumping2));
 sky130_fd_sc_hd__dfxtp_1 _2186_ (.CLK(clknet_leaf_60_clk),
    .D(wCond),
    .Q(rCond));
 sky130_fd_sc_hd__dfxtp_1 _2187_ (.CLK(clknet_leaf_67_clk),
    .D(wStall1),
    .Q(rStall2));
 sky130_fd_sc_hd__dfxtp_1 _2188_ (.CLK(clknet_leaf_60_clk),
    .D(_0000_),
    .Q(rHazardStallRs1));
 sky130_fd_sc_hd__dfxtp_1 _2189_ (.CLK(clknet_leaf_60_clk),
    .D(_0001_),
    .Q(rHazardStallRs2));
 sky130_fd_sc_hd__dfxtp_1 _2190_ (.CLK(clknet_leaf_67_clk),
    .D(_0034_),
    .Q(rRegWrEn));
 sky130_fd_sc_hd__clkbuf_1 _2191_ (.A(wRamWordEn),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _2192_ (.A(wRamHalfEn),
    .X(net69));
 sky130_fd_sc_hd__buf_1 _2193_ (.A(wRamByteEn),
    .X(net70));
 sky130_fd_sc_hd__nand2_2 \alu/_1341_  (.A(\wAluA[0] ),
    .B(net226),
    .Y(\alu/_0057_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1342_  (.A(\alu/_0057_ ),
    .Y(\alu/_0068_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1343_  (.A(\wAluA[0] ),
    .B(net225),
    .Y(\alu/_0079_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1344_  (.A(net191),
    .Y(\alu/_0089_ ));
 sky130_fd_sc_hd__inv_4 \alu/_1345_  (.A(net210),
    .Y(\alu/_0100_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1346_  (.A(\alu/_0089_ ),
    .B(\alu/_0100_ ),
    .Y(\alu/_0111_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1347_  (.A(net191),
    .B(net211),
    .Y(\alu/_0121_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1348_  (.A(\alu/_0111_ ),
    .B(\alu/_0121_ ),
    .Y(\alu/_0132_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1349_  (.A(\wAluA[3] ),
    .Y(\alu/_0143_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1350_  (.A(\alu/_0143_ ),
    .B(net197),
    .Y(\alu/_0153_ ));
 sky130_fd_sc_hd__inv_4 \alu/_1351_  (.A(net196),
    .Y(\alu/_0164_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1352_  (.A(\alu/_0164_ ),
    .B(\wAluA[3] ),
    .Y(\alu/_0174_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1353_  (.A(\alu/_0153_ ),
    .B(\alu/_0174_ ),
    .Y(\alu/_0185_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1354_  (.A(\wAluA[2] ),
    .Y(\alu/_0196_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1355_  (.A(\alu/_0196_ ),
    .B(net176),
    .Y(\alu/_0206_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1356_  (.A(net179),
    .Y(\alu/_0217_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1357_  (.A(\alu/_0217_ ),
    .B(\wAluA[2] ),
    .Y(\alu/_0227_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1358_  (.A(\alu/_0206_ ),
    .B(\alu/_0227_ ),
    .Y(\alu/_0238_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1359_  (.A(\alu/_0185_ ),
    .B(\alu/_0238_ ),
    .Y(\alu/_0249_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_1360_  (.A1(\alu/_0068_ ),
    .A2(\alu/_0079_ ),
    .B1(\alu/_0132_ ),
    .C1(\alu/_0249_ ),
    .X(\alu/_0259_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1361_  (.A(\wAluB[9] ),
    .Y(\alu/_0270_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1362_  (.A(\alu/_0270_ ),
    .B(\wAluA[9] ),
    .Y(\alu/_0281_ ));
 sky130_fd_sc_hd__inv_4 \alu/_1363_  (.A(\wAluA[9] ),
    .Y(\alu/_0291_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1364_  (.A(\alu/_0291_ ),
    .B(\wAluB[9] ),
    .Y(\alu/_0302_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1365_  (.A(\alu/_0281_ ),
    .B(\alu/_0302_ ),
    .Y(\alu/_0313_ ));
 sky130_fd_sc_hd__nand2b_1 \alu/_1366_  (.A_N(net194),
    .B(\wAluB[8] ),
    .Y(\alu/_0323_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1367_  (.A(\wAluB[8] ),
    .Y(\alu/_0334_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1368_  (.A(\alu/_0334_ ),
    .B(net194),
    .Y(\alu/_0344_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1369_  (.A(\alu/_0323_ ),
    .B(\alu/_0344_ ),
    .Y(\alu/_0355_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1370_  (.A(\alu/_0313_ ),
    .B(\alu/_0355_ ),
    .Y(\alu/_0366_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1371_  (.A(\wAluB[11] ),
    .Y(\alu/_0376_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1372_  (.A(\alu/_0376_ ),
    .B(net237),
    .Y(\alu/_0387_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1373_  (.A(net237),
    .Y(\alu/_0397_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1374_  (.A(\alu/_0397_ ),
    .B(\wAluB[11] ),
    .Y(\alu/_0408_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1375_  (.A(\alu/_0387_ ),
    .B(\alu/_0408_ ),
    .Y(\alu/_0419_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1376_  (.A(\wAluA[10] ),
    .Y(\alu/_0429_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1377_  (.A(\alu/_0429_ ),
    .B(\wAluB[10] ),
    .Y(\alu/_0440_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1378_  (.A(\wAluB[10] ),
    .Y(\alu/_0450_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1379_  (.A(\alu/_0450_ ),
    .B(\wAluA[10] ),
    .Y(\alu/_0461_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1380_  (.A(\alu/_0440_ ),
    .B(\alu/_0461_ ),
    .Y(\alu/_0472_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1381_  (.A(\alu/_0419_ ),
    .B(\alu/_0472_ ),
    .Y(\alu/_0482_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1382_  (.A(\alu/_0366_ ),
    .B(\alu/_0482_ ),
    .Y(\alu/_0493_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1383_  (.A(\wAluA[13] ),
    .Y(\alu/_0502_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1384_  (.A(\alu/_0502_ ),
    .B(\wAluB[13] ),
    .Y(\alu/_0503_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1385_  (.A(\wAluB[13] ),
    .Y(\alu/_0504_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1386_  (.A(\alu/_0504_ ),
    .B(\wAluA[13] ),
    .Y(\alu/_0505_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1387_  (.A(\alu/_0503_ ),
    .B(\alu/_0505_ ),
    .Y(\alu/_0506_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1388_  (.A(\wAluA[12] ),
    .Y(\alu/_0507_ ));
 sky130_fd_sc_hd__inv_4 \alu/_1389_  (.A(\wAluB[12] ),
    .Y(\alu/_0508_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1390_  (.A(\alu/_0507_ ),
    .B(\alu/_0508_ ),
    .Y(\alu/_0509_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1391_  (.A(\wAluA[12] ),
    .B(\wAluB[12] ),
    .Y(\alu/_0510_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1392_  (.A(\alu/_0509_ ),
    .B(\alu/_0510_ ),
    .Y(\alu/_0511_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1393_  (.A(\alu/_0511_ ),
    .Y(\alu/_0512_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1394_  (.A(\alu/_0506_ ),
    .B(\alu/_0512_ ),
    .Y(\alu/_0513_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1395_  (.A(\wAluB[15] ),
    .Y(\alu/_0514_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1396_  (.A(\alu/_0514_ ),
    .B(\wAluA[15] ),
    .Y(\alu/_0515_ ));
 sky130_fd_sc_hd__inv_4 \alu/_1397_  (.A(\wAluA[15] ),
    .Y(\alu/_0516_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1398_  (.A(\alu/_0516_ ),
    .B(\wAluB[15] ),
    .Y(\alu/_0517_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1399_  (.A(\alu/_0515_ ),
    .B(\alu/_0517_ ),
    .Y(\alu/_0518_ ));
 sky130_fd_sc_hd__buf_6 \alu/_1400_  (.A(\alu/_0518_ ),
    .X(\alu/_0519_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1401_  (.A(\wAluA[14] ),
    .Y(\alu/_0520_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1402_  (.A(\alu/_0520_ ),
    .B(\wAluB[14] ),
    .Y(\alu/_0521_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1403_  (.A(\wAluB[14] ),
    .Y(\alu/_0522_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1404_  (.A(\alu/_0522_ ),
    .B(\wAluA[14] ),
    .Y(\alu/_0523_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1405_  (.A(\alu/_0521_ ),
    .B(\alu/_0523_ ),
    .Y(\alu/_0524_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1406_  (.A(\alu/_0519_ ),
    .B(\alu/_0524_ ),
    .Y(\alu/_0525_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1407_  (.A(\alu/_0513_ ),
    .B(\alu/_0525_ ),
    .Y(\alu/_0526_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1408_  (.A(\alu/_0493_ ),
    .B(\alu/_0526_ ),
    .Y(\alu/_0527_ ));
 sky130_fd_sc_hd__inv_4 \alu/_1409_  (.A(\wAluA[6] ),
    .Y(\alu/_0528_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1410_  (.A(\alu/_0528_ ),
    .B(\wAluB[6] ),
    .Y(\alu/_0529_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1411_  (.A(\wAluB[6] ),
    .Y(\alu/_0530_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1412_  (.A(\alu/_0530_ ),
    .B(\wAluA[6] ),
    .Y(\alu/_0531_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1413_  (.A(\alu/_0529_ ),
    .B(\alu/_0531_ ),
    .Y(\alu/_0532_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1414_  (.A(net190),
    .Y(\alu/_0533_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1415_  (.A(\alu/_0533_ ),
    .B(\wAluB[7] ),
    .Y(\alu/_0534_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1416_  (.A(\wAluB[7] ),
    .Y(\alu/_0535_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1417_  (.A(\alu/_0535_ ),
    .B(net190),
    .Y(\alu/_0536_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1418_  (.A(\alu/_0534_ ),
    .B(\alu/_0536_ ),
    .Y(\alu/_0537_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1419_  (.A(\alu/_0532_ ),
    .B(\alu/_0537_ ),
    .Y(\alu/_0538_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1420_  (.A(\alu/_0538_ ),
    .Y(\alu/_0539_ ));
 sky130_fd_sc_hd__inv_6 \alu/_1421_  (.A(\wAluA[5] ),
    .Y(\alu/_0540_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1422_  (.A(\wAluB[5] ),
    .B(\alu/_0540_ ),
    .Y(\alu/_0541_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1423_  (.A(\alu/_0541_ ),
    .Y(\alu/_0542_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1424_  (.A(\alu/_0540_ ),
    .B(\wAluB[5] ),
    .Y(\alu/_0543_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1425_  (.A(\alu/_0542_ ),
    .B(\alu/_0543_ ),
    .Y(\alu/_0544_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1426_  (.A(\alu/_0544_ ),
    .Y(\alu/_0545_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1427_  (.A(\wAluA[4] ),
    .Y(\alu/_0546_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1428_  (.A(\alu/_0546_ ),
    .B(net173),
    .Y(\alu/_0547_ ));
 sky130_fd_sc_hd__inv_4 \alu/_1429_  (.A(net169),
    .Y(\alu/_0548_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1430_  (.A(\alu/_0548_ ),
    .B(\wAluA[4] ),
    .Y(\alu/_0549_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1431_  (.A(\alu/_0547_ ),
    .B(\alu/_0549_ ),
    .Y(\alu/_0550_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1432_  (.A(\alu/_0550_ ),
    .Y(\alu/_0551_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1433_  (.A(\alu/_0545_ ),
    .B(\alu/_0551_ ),
    .Y(\alu/_0552_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1434_  (.A(\alu/_0539_ ),
    .B(\alu/_0552_ ),
    .Y(\alu/_0553_ ));
 sky130_fd_sc_hd__and3_1 \alu/_1435_  (.A(\alu/_0259_ ),
    .B(\alu/_0527_ ),
    .C(\alu/_0553_ ),
    .X(\alu/_0554_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1436_  (.A(\wAluA[25] ),
    .Y(\alu/_0555_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1437_  (.A(\wAluB[25] ),
    .Y(\alu/_0556_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1438_  (.A(\alu/_0555_ ),
    .B(\alu/_0556_ ),
    .Y(\alu/_0557_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1439_  (.A(\wAluA[25] ),
    .B(\wAluB[25] ),
    .Y(\alu/_0558_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1440_  (.A(\alu/_0557_ ),
    .B(\alu/_0558_ ),
    .Y(\alu/_0559_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1441_  (.A(\alu/_0559_ ),
    .Y(\alu/_0560_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1442_  (.A(\wAluA[24] ),
    .Y(\alu/_0561_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1443_  (.A(\wAluB[24] ),
    .B(\alu/_0561_ ),
    .X(\alu/_0562_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1444_  (.A(\alu/_0561_ ),
    .B(\wAluB[24] ),
    .Y(\alu/_0563_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1445_  (.A(\alu/_0562_ ),
    .B(\alu/_0563_ ),
    .Y(\alu/_0564_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1446_  (.A(\alu/_0560_ ),
    .B(\alu/_0564_ ),
    .Y(\alu/_0565_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1447_  (.A(\wAluA[27] ),
    .Y(\alu/_0566_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1448_  (.A(\wAluB[27] ),
    .B(\alu/_0566_ ),
    .Y(\alu/_0567_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1449_  (.A(\alu/_0567_ ),
    .Y(\alu/_0568_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1450_  (.A(\alu/_0566_ ),
    .B(\wAluB[27] ),
    .Y(\alu/_0569_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1451_  (.A(\alu/_0568_ ),
    .B(\alu/_0569_ ),
    .Y(\alu/_0570_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1452_  (.A(\wAluA[26] ),
    .Y(\alu/_0571_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1453_  (.A(\wAluB[26] ),
    .B(\alu/_0571_ ),
    .Y(\alu/_0572_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1454_  (.A(\alu/_0572_ ),
    .Y(\alu/_0573_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1455_  (.A(\alu/_0571_ ),
    .B(\wAluB[26] ),
    .Y(\alu/_0574_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1456_  (.A(\alu/_0573_ ),
    .B(\alu/_0574_ ),
    .Y(\alu/_0575_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1457_  (.A(\alu/_0570_ ),
    .B(\alu/_0575_ ),
    .Y(\alu/_0576_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1458_  (.A(\alu/_0565_ ),
    .B(\alu/_0576_ ),
    .Y(\alu/_0577_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1459_  (.A(net192),
    .Y(\alu/_0578_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1460_  (.A(\wAluB[31] ),
    .B(\alu/_0578_ ),
    .Y(\alu/_0579_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1461_  (.A(\alu/_0578_ ),
    .B(\wAluB[31] ),
    .Y(\alu/_0580_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1462_  (.A(\alu/_0580_ ),
    .Y(\alu/_0581_ ));
 sky130_fd_sc_hd__nor2_2 \alu/_1463_  (.A(\alu/_0579_ ),
    .B(\alu/_0581_ ),
    .Y(\alu/_0582_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1464_  (.A(\alu/_0582_ ),
    .Y(\alu/_0583_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1465_  (.A(\wAluA[30] ),
    .Y(\alu/_0584_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1466_  (.A(\wAluB[30] ),
    .B(\alu/_0584_ ),
    .Y(\alu/_0585_ ));
 sky130_fd_sc_hd__and2_1 \alu/_1467_  (.A(\alu/_0584_ ),
    .B(\wAluB[30] ),
    .X(\alu/_0586_ ));
 sky130_fd_sc_hd__or2_2 \alu/_1468_  (.A(\alu/_0585_ ),
    .B(\alu/_0586_ ),
    .X(\alu/_0587_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1469_  (.A(\alu/_0583_ ),
    .B(\alu/_0587_ ),
    .Y(\alu/_0588_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1470_  (.A(\wAluA[29] ),
    .Y(\alu/_0589_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1471_  (.A(\wAluB[29] ),
    .B(\alu/_0589_ ),
    .X(\alu/_0590_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1472_  (.A(\alu/_0589_ ),
    .B(\wAluB[29] ),
    .Y(\alu/_0591_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1473_  (.A(\alu/_0590_ ),
    .B(\alu/_0591_ ),
    .Y(\alu/_0592_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1474_  (.A(\wAluB[28] ),
    .Y(\alu/_0593_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1475_  (.A(net236),
    .B(\alu/_0593_ ),
    .X(\alu/_0594_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1476_  (.A(\alu/_0593_ ),
    .B(net236),
    .Y(\alu/_0595_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1477_  (.A(\alu/_0594_ ),
    .B(\alu/_0595_ ),
    .Y(\alu/_0596_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1478_  (.A(\alu/_0592_ ),
    .B(\alu/_0596_ ),
    .Y(\alu/_0597_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1479_  (.A(\alu/_0588_ ),
    .B(\alu/_0597_ ),
    .Y(\alu/_0598_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1480_  (.A(\alu/_0577_ ),
    .B(\alu/_0598_ ),
    .Y(\alu/_0599_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1481_  (.A(\wAluA[19] ),
    .Y(\alu/_0600_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1482_  (.A(\wAluB[19] ),
    .Y(\alu/_0601_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1483_  (.A(\alu/_0600_ ),
    .B(\alu/_0601_ ),
    .Y(\alu/_0602_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1484_  (.A(\wAluA[19] ),
    .B(\wAluB[19] ),
    .Y(\alu/_0603_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1485_  (.A(\alu/_0602_ ),
    .B(\alu/_0603_ ),
    .Y(\alu/_0604_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1486_  (.A(\alu/_0604_ ),
    .Y(\alu/_0605_ ));
 sky130_fd_sc_hd__inv_4 \alu/_1487_  (.A(\wAluA[18] ),
    .Y(\alu/_0606_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1488_  (.A(\wAluB[18] ),
    .B(\alu/_0606_ ),
    .X(\alu/_0607_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1489_  (.A(\alu/_0606_ ),
    .B(\wAluB[18] ),
    .Y(\alu/_0608_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1490_  (.A(\alu/_0607_ ),
    .B(\alu/_0608_ ),
    .Y(\alu/_0609_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1491_  (.A(\alu/_0605_ ),
    .B(\alu/_0609_ ),
    .Y(\alu/_0610_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1492_  (.A(\wAluA[16] ),
    .B(\wAluB[16] ),
    .Y(\alu/_0611_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1493_  (.A(\wAluA[16] ),
    .B(\wAluB[16] ),
    .Y(\alu/_0612_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1494_  (.A(\alu/_0612_ ),
    .Y(\alu/_0613_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1495_  (.A(\alu/_0611_ ),
    .B(\alu/_0613_ ),
    .Y(\alu/_0614_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1496_  (.A(\wAluA[17] ),
    .Y(\alu/_0615_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1497_  (.A(\wAluB[17] ),
    .Y(\alu/_0616_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1498_  (.A(\alu/_0615_ ),
    .B(\alu/_0616_ ),
    .Y(\alu/_0617_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1499_  (.A(\wAluA[17] ),
    .B(\wAluB[17] ),
    .Y(\alu/_0618_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1500_  (.A(\alu/_0617_ ),
    .B(\alu/_0618_ ),
    .Y(\alu/_0619_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1501_  (.A(\alu/_0619_ ),
    .Y(\alu/_0620_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1502_  (.A(\alu/_0614_ ),
    .B(\alu/_0620_ ),
    .Y(\alu/_0621_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1503_  (.A(\alu/_0610_ ),
    .B(\alu/_0621_ ),
    .Y(\alu/_0622_ ));
 sky130_fd_sc_hd__inv_4 \alu/_1504_  (.A(\wAluA[23] ),
    .Y(\alu/_0623_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1505_  (.A(\wAluB[23] ),
    .B(\alu/_0623_ ),
    .X(\alu/_0624_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1506_  (.A(\alu/_0623_ ),
    .B(\wAluB[23] ),
    .Y(\alu/_0625_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1507_  (.A(\alu/_0624_ ),
    .B(\alu/_0625_ ),
    .Y(\alu/_0626_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1508_  (.A(net193),
    .Y(\alu/_0627_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1509_  (.A(\wAluB[22] ),
    .B(\alu/_0627_ ),
    .X(\alu/_0628_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1510_  (.A(\alu/_0627_ ),
    .B(\wAluB[22] ),
    .Y(\alu/_0629_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1511_  (.A(\alu/_0628_ ),
    .B(\alu/_0629_ ),
    .Y(\alu/_0630_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1512_  (.A(\alu/_0626_ ),
    .B(\alu/_0630_ ),
    .Y(\alu/_0631_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1513_  (.A(\wAluA[21] ),
    .Y(\alu/_0632_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1514_  (.A(\wAluB[21] ),
    .Y(\alu/_0633_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1515_  (.A(\alu/_0632_ ),
    .B(\alu/_0633_ ),
    .Y(\alu/_0634_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1516_  (.A(\wAluA[21] ),
    .B(\wAluB[21] ),
    .Y(\alu/_0635_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1517_  (.A(\alu/_0634_ ),
    .B(\alu/_0635_ ),
    .Y(\alu/_0636_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1518_  (.A(\alu/_0636_ ),
    .Y(\alu/_0637_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1519_  (.A(\wAluA[20] ),
    .Y(\alu/_0638_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1520_  (.A(\wAluB[20] ),
    .Y(\alu/_0639_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1521_  (.A(\alu/_0638_ ),
    .B(\alu/_0639_ ),
    .Y(\alu/_0640_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1522_  (.A(\wAluA[20] ),
    .B(\wAluB[20] ),
    .Y(\alu/_0641_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1523_  (.A(\alu/_0640_ ),
    .B(\alu/_0641_ ),
    .Y(\alu/_0642_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1524_  (.A(\alu/_0642_ ),
    .Y(\alu/_0643_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1525_  (.A(\alu/_0637_ ),
    .B(\alu/_0643_ ),
    .Y(\alu/_0644_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1526_  (.A(\alu/_0631_ ),
    .B(\alu/_0644_ ),
    .Y(\alu/_0645_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1527_  (.A(\alu/_0622_ ),
    .B(\alu/_0645_ ),
    .Y(\alu/_0646_ ));
 sky130_fd_sc_hd__and2_1 \alu/_1528_  (.A(\alu/_0599_ ),
    .B(\alu/_0646_ ),
    .X(\alu/_0647_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1529_  (.A(\wFunct3_aluIn[1] ),
    .Y(\alu/_0648_ ));
 sky130_fd_sc_hd__o31a_2 \alu/_1530_  (.A1(op_consShf),
    .A2(r_type),
    .A3(net897),
    .B1(\wFunct7_aluIn[5] ),
    .X(\alu/_0649_ ));
 sky130_fd_sc_hd__nor2_2 \alu/_1531_  (.A(\wFunct3_aluIn[0] ),
    .B(\alu/_0649_ ),
    .Y(\alu/_0650_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1532_  (.A(\alu/_0650_ ),
    .Y(\alu/_0651_ ));
 sky130_fd_sc_hd__a2111o_1 \alu/_1533_  (.A1(\alu/_0554_ ),
    .A2(\alu/_0647_ ),
    .B1(\wFunct3_aluIn[2] ),
    .C1(\alu/_0648_ ),
    .D1(\alu/_0651_ ),
    .X(\alu/_0652_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1534_  (.A(\alu/_0652_ ),
    .Y(\alu/_0653_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1535_  (.A(\alu/_0610_ ),
    .Y(\alu/_0654_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \alu/_1536_  (.A(\alu/_0619_ ),
    .X(\alu/_0655_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1537_  (.A(\wAluA[16] ),
    .Y(\alu/_0656_ ));
 sky130_fd_sc_hd__and3_1 \alu/_1538_  (.A(\alu/_0655_ ),
    .B(\alu/_0656_ ),
    .C(\wAluB[16] ),
    .X(\alu/_0657_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_1539_  (.A1(\alu/_0615_ ),
    .A2(\wAluB[17] ),
    .B1(\alu/_0657_ ),
    .Y(\alu/_0658_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1540_  (.A(\alu/_0600_ ),
    .B(\wAluB[19] ),
    .Y(\alu/_0659_ ));
 sky130_fd_sc_hd__o221ai_1 \alu/_1541_  (.A1(\alu/_0605_ ),
    .A2(\alu/_0608_ ),
    .B1(\alu/_0654_ ),
    .B2(\alu/_0658_ ),
    .C1(\alu/_0659_ ),
    .Y(\alu/_0660_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1542_  (.A(\alu/_0645_ ),
    .Y(\alu/_0661_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1543_  (.A(\alu/_0660_ ),
    .B(\alu/_0661_ ),
    .Y(\alu/_0662_ ));
 sky130_fd_sc_hd__buf_6 \alu/_1544_  (.A(\alu/_0626_ ),
    .X(\alu/_0663_ ));
 sky130_fd_sc_hd__buf_6 \alu/_1545_  (.A(\alu/_0636_ ),
    .X(\alu/_0664_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1546_  (.A(\wAluA[21] ),
    .B(\alu/_0633_ ),
    .Y(\alu/_0665_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_1547_  (.A1(\alu/_0664_ ),
    .A2(\alu/_0638_ ),
    .A3(\wAluB[20] ),
    .B1(\alu/_0665_ ),
    .X(\alu/_0666_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1548_  (.A(\alu/_0666_ ),
    .B(\alu/_0631_ ),
    .Y(\alu/_0667_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_1549_  (.A1(\alu/_0663_ ),
    .A2(\alu/_0629_ ),
    .B1(\alu/_0625_ ),
    .C1(\alu/_0667_ ),
    .X(\alu/_0668_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1550_  (.A(\alu/_0662_ ),
    .B(\alu/_0668_ ),
    .Y(\alu/_0669_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1551_  (.A(\wAluB[25] ),
    .B(\alu/_0555_ ),
    .Y(\alu/_0670_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1552_  (.A(\alu/_0670_ ),
    .Y(\alu/_0671_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1553_  (.A1(\wAluA[25] ),
    .A2(\alu/_0556_ ),
    .B1(\alu/_0563_ ),
    .Y(\alu/_0672_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1554_  (.A(\alu/_0569_ ),
    .B(\alu/_0574_ ),
    .Y(\alu/_0673_ ));
 sky130_fd_sc_hd__a32o_1 \alu/_1555_  (.A1(\alu/_0576_ ),
    .A2(\alu/_0671_ ),
    .A3(\alu/_0672_ ),
    .B1(\alu/_0568_ ),
    .B2(\alu/_0673_ ),
    .X(\alu/_0674_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1556_  (.A1(\alu/_0582_ ),
    .A2(\alu/_0586_ ),
    .B1(\alu/_0581_ ),
    .X(\alu/_0675_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1557_  (.A(\alu/_0594_ ),
    .B(\alu/_0591_ ),
    .Y(\alu/_0676_ ));
 sky130_fd_sc_hd__and3_1 \alu/_1558_  (.A(\alu/_0588_ ),
    .B(\alu/_0590_ ),
    .C(\alu/_0676_ ),
    .X(\alu/_0677_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1559_  (.A(\alu/_0675_ ),
    .B(\alu/_0677_ ),
    .X(\alu/_0678_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_1560_  (.A1(\alu/_0674_ ),
    .A2(\alu/_0588_ ),
    .A3(\alu/_0597_ ),
    .B1(\alu/_0678_ ),
    .X(\alu/_0679_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_1561_  (.A1(\alu/_0669_ ),
    .A2(\alu/_0599_ ),
    .B1(\alu/_0679_ ),
    .Y(\alu/_0680_ ));
 sky130_fd_sc_hd__o31a_1 \alu/_1562_  (.A1(\wAluA[12] ),
    .A2(\alu/_0508_ ),
    .A3(\alu/_0506_ ),
    .B1(\alu/_0503_ ),
    .X(\alu/_0681_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_1563_  (.A1(\alu/_0521_ ),
    .A2(\alu/_0519_ ),
    .B1(\alu/_0517_ ),
    .X(\alu/_0682_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1564_  (.A1(\alu/_0323_ ),
    .A2(\alu/_0313_ ),
    .B1(\alu/_0302_ ),
    .Y(\alu/_0683_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1565_  (.A(\alu/_0683_ ),
    .B(\alu/_0482_ ),
    .Y(\alu/_0684_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1566_  (.A(\alu/_0440_ ),
    .B(\alu/_0419_ ),
    .X(\alu/_0685_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_1567_  (.A1(\alu/_0684_ ),
    .A2(\alu/_0408_ ),
    .A3(\alu/_0685_ ),
    .B1(\alu/_0526_ ),
    .X(\alu/_0686_ ));
 sky130_fd_sc_hd__o311a_1 \alu/_1568_  (.A1(\alu/_0519_ ),
    .A2(\alu/_0524_ ),
    .A3(\alu/_0681_ ),
    .B1(\alu/_0682_ ),
    .C1(\alu/_0686_ ),
    .X(\alu/_0687_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1569_  (.A1(\alu/_0547_ ),
    .A2(\alu/_0543_ ),
    .B1(\alu/_0541_ ),
    .X(\alu/_0688_ ));
 sky130_fd_sc_hd__o221a_1 \alu/_1570_  (.A1(\alu/_0529_ ),
    .A2(\alu/_0537_ ),
    .B1(\alu/_0688_ ),
    .B2(\alu/_0539_ ),
    .C1(\alu/_0534_ ),
    .X(\alu/_0689_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1571_  (.A1(\alu/_0206_ ),
    .A2(\alu/_0185_ ),
    .B1(\alu/_0153_ ),
    .Y(\alu/_0690_ ));
 sky130_fd_sc_hd__inv_4 \alu/_1572_  (.A(net234),
    .Y(\alu/_0691_ ));
 sky130_fd_sc_hd__buf_6 \alu/_1573_  (.A(\alu/_0691_ ),
    .X(\alu/_0692_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1574_  (.A(\alu/_0692_ ),
    .B(\wAluA[0] ),
    .Y(\alu/_0693_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1575_  (.A(\alu/_0693_ ),
    .B(net211),
    .Y(\alu/_0694_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1576_  (.A(\alu/_0694_ ),
    .B(\wAluA[1] ),
    .Y(\alu/_0695_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1577_  (.A(net211),
    .B(\alu/_0693_ ),
    .Y(\alu/_0696_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1578_  (.A(\alu/_0696_ ),
    .Y(\alu/_0697_ ));
 sky130_fd_sc_hd__and3_1 \alu/_1579_  (.A(\alu/_0249_ ),
    .B(\alu/_0695_ ),
    .C(\alu/_0697_ ),
    .X(\alu/_0698_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1580_  (.A1(\alu/_0690_ ),
    .A2(\alu/_0698_ ),
    .B1(\alu/_0553_ ),
    .Y(\alu/_0699_ ));
 sky130_fd_sc_hd__a21bo_1 \alu/_1581_  (.A1(\alu/_0689_ ),
    .A2(\alu/_0699_ ),
    .B1_N(\alu/_0527_ ),
    .X(\alu/_0700_ ));
 sky130_fd_sc_hd__a21bo_1 \alu/_1582_  (.A1(\alu/_0687_ ),
    .A2(\alu/_0700_ ),
    .B1_N(\alu/_0647_ ),
    .X(\alu/_0701_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_1583_  (.A(\alu/_0680_ ),
    .B(\alu/_0701_ ),
    .C(\alu/_0582_ ),
    .Y(\alu/_0702_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_1584_  (.A(\alu/_0653_ ),
    .B(\alu/_0702_ ),
    .C(\alu/_0580_ ),
    .Y(\alu/_0703_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1585_  (.A(\alu/_0217_ ),
    .X(\alu/_0704_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1586_  (.A(\alu/_0704_ ),
    .X(\alu/_0705_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1587_  (.A0(\alu/_0546_ ),
    .A1(\alu/_0540_ ),
    .S(net225),
    .X(\alu/_0706_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1588_  (.A0(\alu/_0528_ ),
    .A1(\alu/_0533_ ),
    .S(net225),
    .X(\alu/_0707_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1589_  (.A0(\alu/_0706_ ),
    .A1(\alu/_0707_ ),
    .S(net208),
    .X(\alu/_0708_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1590_  (.A(\alu/_0164_ ),
    .X(\alu/_0709_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1591_  (.A(\alu/_0709_ ),
    .X(\alu/_0710_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1592_  (.A(\alu/_0710_ ),
    .X(\alu/_0711_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1593_  (.A0(\alu/_0196_ ),
    .A1(\alu/_0143_ ),
    .S(net226),
    .X(\alu/_0712_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1594_  (.A(net226),
    .B(net191),
    .Y(\alu/_0713_ ));
 sky130_fd_sc_hd__and2_1 \alu/_1595_  (.A(\alu/_0693_ ),
    .B(\alu/_0713_ ),
    .X(\alu/_0714_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1596_  (.A(\alu/_0100_ ),
    .X(\alu/_0715_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1597_  (.A(\alu/_0715_ ),
    .X(\alu/_0716_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1598_  (.A0(\alu/_0712_ ),
    .A1(\alu/_0714_ ),
    .S(\alu/_0716_ ),
    .X(\alu/_0717_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1599_  (.A(net175),
    .B(\alu/_0717_ ),
    .X(\alu/_0718_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_1600_  (.A1(\alu/_0705_ ),
    .A2(\alu/_0708_ ),
    .B1(\alu/_0711_ ),
    .C1(\alu/_0718_ ),
    .X(\alu/_0719_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1601_  (.A(\alu/_0710_ ),
    .X(\alu/_0720_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1602_  (.A(\alu/_0720_ ),
    .X(\alu/_0721_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1603_  (.A0(net194),
    .A1(\wAluA[9] ),
    .S(net228),
    .X(\alu/_0722_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1604_  (.A0(\wAluA[10] ),
    .A1(net237),
    .S(net222),
    .X(\alu/_0723_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1605_  (.A0(\alu/_0722_ ),
    .A1(\alu/_0723_ ),
    .S(net208),
    .X(\alu/_0724_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1606_  (.A0(\wAluA[12] ),
    .A1(\wAluA[13] ),
    .S(net223),
    .X(\alu/_0725_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1607_  (.A0(\wAluA[14] ),
    .A1(\wAluA[15] ),
    .S(net223),
    .X(\alu/_0726_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1608_  (.A0(\alu/_0725_ ),
    .A1(\alu/_0726_ ),
    .S(net209),
    .X(\alu/_0727_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1609_  (.A0(\alu/_0724_ ),
    .A1(\alu/_0727_ ),
    .S(net175),
    .X(\alu/_0728_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1610_  (.A(\wFunct3_aluIn[2] ),
    .Y(\alu/_0729_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1611_  (.A(\wFunct3_aluIn[1] ),
    .B(\alu/_0729_ ),
    .Y(\alu/_0730_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1612_  (.A(\alu/_0730_ ),
    .B(\wFunct3_aluIn[0] ),
    .Y(\alu/_0731_ ));
 sky130_fd_sc_hd__nor2_2 \alu/_1613_  (.A(net169),
    .B(\alu/_0731_ ),
    .Y(\alu/_0732_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1614_  (.A(\alu/_0732_ ),
    .X(\alu/_0733_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1615_  (.A1(\alu/_0721_ ),
    .A2(\alu/_0728_ ),
    .B1(\alu/_0733_ ),
    .Y(\alu/_0734_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1616_  (.A(\wFunct3_aluIn[0] ),
    .Y(\alu/_0735_ ));
 sky130_fd_sc_hd__nor2_2 \alu/_1617_  (.A(\alu/_0735_ ),
    .B(\alu/_0649_ ),
    .Y(\alu/_0736_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1618_  (.A(\wFunct3_aluIn[2] ),
    .B(\wFunct3_aluIn[1] ),
    .Y(\alu/_0737_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1619_  (.A(\alu/_0737_ ),
    .Y(\alu/_0738_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1620_  (.A(\alu/_0736_ ),
    .B(\alu/_0738_ ),
    .Y(\alu/_0739_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1621_  (.A(\alu/_0739_ ),
    .X(\alu/_0740_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1622_  (.A(\alu/_0740_ ),
    .X(\alu/_0741_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1623_  (.A(net176),
    .B(\alu/_0697_ ),
    .Y(\alu/_0742_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1624_  (.A(\alu/_0742_ ),
    .B(\alu/_0710_ ),
    .Y(\alu/_0743_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1625_  (.A(\wFunct3_aluIn[2] ),
    .B(\wFunct3_aluIn[1] ),
    .Y(\alu/_0744_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1626_  (.A(\alu/_0736_ ),
    .B(\alu/_0744_ ),
    .Y(\alu/_0745_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1627_  (.A(net171),
    .B(\alu/_0745_ ),
    .Y(\alu/_0746_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1628_  (.A(\alu/_0746_ ),
    .Y(\alu/_0747_ ));
 sky130_fd_sc_hd__o22a_1 \alu/_1629_  (.A1(\alu/_0057_ ),
    .A2(\alu/_0741_ ),
    .B1(\alu/_0743_ ),
    .B2(\alu/_0747_ ),
    .X(\alu/_0748_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1630_  (.A1(\alu/_0719_ ),
    .A2(\alu/_0734_ ),
    .B1(\alu/_0748_ ),
    .Y(\alu/_0749_ ));
 sky130_fd_sc_hd__or3b_1 \alu/_1631_  (.A(\wFunct3_aluIn[2] ),
    .B(\alu/_0648_ ),
    .C_N(\alu/_0736_ ),
    .X(\alu/_0750_ ));
 sky130_fd_sc_hd__nand2b_1 \alu/_1632_  (.A_N(\wAluA[0] ),
    .B(net226),
    .Y(\alu/_0751_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1633_  (.A(\alu/_0132_ ),
    .B(\alu/_0751_ ),
    .Y(\alu/_0752_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1634_  (.A(\alu/_0100_ ),
    .B(net191),
    .Y(\alu/_0753_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1635_  (.A(\alu/_0752_ ),
    .B(\alu/_0753_ ),
    .Y(\alu/_0754_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1636_  (.A(\alu/_0754_ ),
    .B(\alu/_0249_ ),
    .Y(\alu/_0755_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1637_  (.A(net176),
    .B(\alu/_0196_ ),
    .Y(\alu/_0756_ ));
 sky130_fd_sc_hd__a21boi_1 \alu/_1638_  (.A1(\alu/_0756_ ),
    .A2(\alu/_0153_ ),
    .B1_N(\alu/_0174_ ),
    .Y(\alu/_0757_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1639_  (.A(\alu/_0755_ ),
    .B(\alu/_0757_ ),
    .Y(\alu/_0758_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1640_  (.A(\alu/_0758_ ),
    .B(\alu/_0553_ ),
    .Y(\alu/_0759_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1641_  (.A(net173),
    .B(\alu/_0546_ ),
    .Y(\alu/_0760_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1642_  (.A1(\alu/_0760_ ),
    .A2(\alu/_0543_ ),
    .B1(\alu/_0541_ ),
    .X(\alu/_0761_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1643_  (.A1(\alu/_0531_ ),
    .A2(\alu/_0537_ ),
    .B1(\alu/_0536_ ),
    .Y(\alu/_0762_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_1644_  (.A1(\alu/_0761_ ),
    .A2(\alu/_0538_ ),
    .B1(\alu/_0762_ ),
    .Y(\alu/_0763_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1645_  (.A(\alu/_0759_ ),
    .B(\alu/_0763_ ),
    .Y(\alu/_0764_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1646_  (.A(\alu/_0764_ ),
    .B(\alu/_0527_ ),
    .Y(\alu/_0765_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1647_  (.A1(\alu/_0344_ ),
    .A2(\alu/_0313_ ),
    .B1(\alu/_0281_ ),
    .Y(\alu/_0766_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1648_  (.A(\alu/_0766_ ),
    .B(\alu/_0482_ ),
    .Y(\alu/_0767_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_1649_  (.A1(\alu/_0461_ ),
    .A2(\alu/_0419_ ),
    .B1(\alu/_0387_ ),
    .X(\alu/_0768_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1650_  (.A(\alu/_0767_ ),
    .B(\alu/_0768_ ),
    .Y(\alu/_0769_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1651_  (.A(\alu/_0526_ ),
    .Y(\alu/_0770_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1652_  (.A(\alu/_0508_ ),
    .B(\wAluA[12] ),
    .Y(\alu/_0771_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1653_  (.A1(\alu/_0771_ ),
    .A2(\alu/_0506_ ),
    .B1(\alu/_0505_ ),
    .Y(\alu/_0772_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1654_  (.A(\alu/_0772_ ),
    .B(\alu/_0525_ ),
    .Y(\alu/_0773_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_1655_  (.A1(\alu/_0523_ ),
    .A2(\alu/_0519_ ),
    .B1(\alu/_0515_ ),
    .X(\alu/_0774_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1656_  (.A(\alu/_0773_ ),
    .B(\alu/_0774_ ),
    .Y(\alu/_0775_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_1657_  (.A1(\alu/_0769_ ),
    .A2(\alu/_0770_ ),
    .B1(\alu/_0775_ ),
    .Y(\alu/_0776_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1658_  (.A(\alu/_0765_ ),
    .B(\alu/_0776_ ),
    .Y(\alu/_0777_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1659_  (.A(\alu/_0777_ ),
    .B(\alu/_0646_ ),
    .Y(\alu/_0778_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1660_  (.A(\wAluB[16] ),
    .Y(\alu/_0779_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1661_  (.A(\alu/_0779_ ),
    .B(\wAluA[16] ),
    .Y(\alu/_0780_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1662_  (.A(\alu/_0616_ ),
    .B(\wAluA[17] ),
    .Y(\alu/_0781_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1663_  (.A1(\alu/_0780_ ),
    .A2(\alu/_0620_ ),
    .B1(\alu/_0781_ ),
    .Y(\alu/_0782_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1664_  (.A(\alu/_0782_ ),
    .Y(\alu/_0783_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1665_  (.A(\alu/_0601_ ),
    .B(\wAluA[19] ),
    .Y(\alu/_0784_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_1666_  (.A1(\alu/_0607_ ),
    .A2(\alu/_0605_ ),
    .B1(\alu/_0784_ ),
    .X(\alu/_0785_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1667_  (.A1(\alu/_0654_ ),
    .A2(\alu/_0783_ ),
    .B1(\alu/_0785_ ),
    .Y(\alu/_0786_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1668_  (.A(\wAluB[21] ),
    .B(\alu/_0632_ ),
    .Y(\alu/_0787_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_1669_  (.A1(\alu/_0664_ ),
    .A2(\wAluA[20] ),
    .A3(\alu/_0639_ ),
    .B1(\alu/_0787_ ),
    .X(\alu/_0788_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1670_  (.A(\alu/_0788_ ),
    .B(\alu/_0631_ ),
    .Y(\alu/_0789_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_1671_  (.A1(\alu/_0628_ ),
    .A2(\alu/_0663_ ),
    .B1(\alu/_0624_ ),
    .X(\alu/_0790_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1672_  (.A(\alu/_0789_ ),
    .B(\alu/_0790_ ),
    .Y(\alu/_0791_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_1673_  (.A1(\alu/_0786_ ),
    .A2(\alu/_0661_ ),
    .B1(\alu/_0791_ ),
    .Y(\alu/_0792_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1674_  (.A(\alu/_0778_ ),
    .B(\alu/_0792_ ),
    .Y(\alu/_0793_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1675_  (.A(\alu/_0570_ ),
    .Y(\alu/_0794_ ));
 sky130_fd_sc_hd__o21ai_2 \alu/_1676_  (.A1(\alu/_0562_ ),
    .A2(\alu/_0560_ ),
    .B1(\alu/_0671_ ),
    .Y(\alu/_0795_ ));
 sky130_fd_sc_hd__a221oi_4 \alu/_1677_  (.A1(\alu/_0794_ ),
    .A2(\alu/_0572_ ),
    .B1(\alu/_0795_ ),
    .B2(\alu/_0576_ ),
    .C1(\alu/_0567_ ),
    .Y(\alu/_0796_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_1678_  (.A1(\alu/_0595_ ),
    .A2(\alu/_0592_ ),
    .B1(\alu/_0590_ ),
    .X(\alu/_0797_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_1679_  (.A1(\alu/_0585_ ),
    .A2(\alu/_0580_ ),
    .B1(\alu/_0579_ ),
    .Y(\alu/_0798_ ));
 sky130_fd_sc_hd__o31a_1 \alu/_1680_  (.A1(\alu/_0583_ ),
    .A2(\alu/_0587_ ),
    .A3(\alu/_0797_ ),
    .B1(\alu/_0798_ ),
    .X(\alu/_0799_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1681_  (.A1(\alu/_0598_ ),
    .A2(\alu/_0796_ ),
    .B1(\alu/_0799_ ),
    .Y(\alu/_0800_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1682_  (.A1(\alu/_0599_ ),
    .A2(\alu/_0793_ ),
    .B1(\alu/_0800_ ),
    .X(\alu/_0801_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1683_  (.A(\alu/_0750_ ),
    .B(\alu/_0801_ ),
    .Y(\alu/_0802_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1684_  (.A(\alu/_0731_ ),
    .Y(\alu/_0803_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1685_  (.A(\alu/_0803_ ),
    .B(net170),
    .Y(\alu/_0804_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1686_  (.A(\alu/_0720_ ),
    .X(\alu/_0805_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1687_  (.A0(\wAluA[24] ),
    .A1(\wAluA[25] ),
    .S(net229),
    .X(\alu/_0806_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1688_  (.A0(\wAluA[26] ),
    .A1(\wAluA[27] ),
    .S(net230),
    .X(\alu/_0807_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1689_  (.A0(\alu/_0806_ ),
    .A1(\alu/_0807_ ),
    .S(net215),
    .X(\alu/_0808_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1690_  (.A(\alu/_0691_ ),
    .B(\wAluA[30] ),
    .Y(\alu/_0809_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1691_  (.A1(\alu/_0692_ ),
    .A2(\alu/_0578_ ),
    .B1(\alu/_0809_ ),
    .Y(\alu/_0810_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1692_  (.A(\alu/_0692_ ),
    .B(net236),
    .Y(\alu/_0811_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1693_  (.A(net231),
    .B(\wAluA[29] ),
    .Y(\alu/_0812_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1694_  (.A(\alu/_0811_ ),
    .B(\alu/_0812_ ),
    .Y(\alu/_0813_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1695_  (.A0(\alu/_0810_ ),
    .A1(\alu/_0813_ ),
    .S(\alu/_0100_ ),
    .X(\alu/_0814_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1696_  (.A0(\alu/_0808_ ),
    .A1(\alu/_0814_ ),
    .S(net185),
    .X(\alu/_0815_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1697_  (.A(\alu/_0217_ ),
    .X(\alu/_0816_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1698_  (.A(\alu/_0816_ ),
    .X(\alu/_0817_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1699_  (.A(\alu/_0817_ ),
    .X(\alu/_0818_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1700_  (.A0(\wAluA[20] ),
    .A1(\wAluA[21] ),
    .S(net229),
    .X(\alu/_0819_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1701_  (.A0(net193),
    .A1(\wAluA[23] ),
    .S(net230),
    .X(\alu/_0820_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1702_  (.A0(\alu/_0819_ ),
    .A1(\alu/_0820_ ),
    .S(net214),
    .X(\alu/_0821_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1703_  (.A(\alu/_0715_ ),
    .X(\alu/_0822_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1704_  (.A(\alu/_0822_ ),
    .X(\alu/_0823_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1705_  (.A0(\wAluA[18] ),
    .A1(\wAluA[19] ),
    .S(net229),
    .X(\alu/_0824_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1706_  (.A0(\alu/_0656_ ),
    .A1(\alu/_0615_ ),
    .S(net233),
    .X(\alu/_0825_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1707_  (.A(\alu/_0716_ ),
    .X(\alu/_0826_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1708_  (.A(\alu/_0825_ ),
    .B(\alu/_0826_ ),
    .Y(\alu/_0827_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1709_  (.A1(\alu/_0823_ ),
    .A2(\alu/_0824_ ),
    .B1(\alu/_0827_ ),
    .Y(\alu/_0828_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1710_  (.A(\alu/_0828_ ),
    .B(\alu/_0818_ ),
    .Y(\alu/_0829_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1711_  (.A1(\alu/_0818_ ),
    .A2(\alu/_0821_ ),
    .B1(\alu/_0829_ ),
    .Y(\alu/_0830_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1712_  (.A(\alu/_0710_ ),
    .X(\alu/_0831_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1713_  (.A(\alu/_0831_ ),
    .X(\alu/_0832_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1714_  (.A(\alu/_0830_ ),
    .B(\alu/_0832_ ),
    .Y(\alu/_0833_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1715_  (.A1(\alu/_0805_ ),
    .A2(\alu/_0815_ ),
    .B1(\alu/_0833_ ),
    .Y(\alu/_0834_ ));
 sky130_fd_sc_hd__buf_6 \alu/_1716_  (.A(\alu/_0649_ ),
    .X(\alu/_0835_ ));
 sky130_fd_sc_hd__a2111o_1 \alu/_1717_  (.A1(\alu/_0835_ ),
    .A2(\wFunct3_aluIn[2] ),
    .B1(\wFunct3_aluIn[0] ),
    .C1(\wFunct3_aluIn[1] ),
    .D1(\alu/_0068_ ),
    .X(\alu/_0836_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1718_  (.A(\alu/_0650_ ),
    .B(\alu/_0738_ ),
    .Y(\alu/_0837_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1719_  (.A(\alu/_0837_ ),
    .X(\alu/_0838_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1720_  (.A1(\alu/_0836_ ),
    .A2(\alu/_0838_ ),
    .B1(\alu/_0079_ ),
    .X(\alu/_0839_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1721_  (.A1(\alu/_0804_ ),
    .A2(\alu/_0834_ ),
    .B1(\alu/_0839_ ),
    .Y(\alu/_0840_ ));
 sky130_fd_sc_hd__nor3_1 \alu/_1722_  (.A(\alu/_0749_ ),
    .B(\alu/_0802_ ),
    .C(\alu/_0840_ ),
    .Y(\alu/_0841_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1723_  (.A(\alu/_0703_ ),
    .B(\alu/_0841_ ),
    .Y(\wAluOut[0] ));
 sky130_fd_sc_hd__nor2_1 \alu/_1724_  (.A(net234),
    .B(\alu/_0578_ ),
    .Y(\alu/_0842_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1725_  (.A(net234),
    .B(\wAluA[30] ),
    .Y(\alu/_0843_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1726_  (.A1(net234),
    .A2(\alu/_0589_ ),
    .B1(\alu/_0843_ ),
    .Y(\alu/_0844_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1727_  (.A(\alu/_0715_ ),
    .X(\alu/_0845_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1728_  (.A(\alu/_0844_ ),
    .B(\alu/_0845_ ),
    .Y(\alu/_0846_ ));
 sky130_fd_sc_hd__a21bo_1 \alu/_1729_  (.A1(net218),
    .A2(\alu/_0842_ ),
    .B1_N(\alu/_0846_ ),
    .X(\alu/_0847_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1730_  (.A0(\wAluA[25] ),
    .A1(\wAluA[26] ),
    .S(net232),
    .X(\alu/_0848_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1731_  (.A0(\wAluA[27] ),
    .A1(\wAluA[28] ),
    .S(net231),
    .X(\alu/_0849_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1732_  (.A0(\alu/_0848_ ),
    .A1(\alu/_0849_ ),
    .S(net216),
    .X(\alu/_0850_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1733_  (.A(\alu/_0816_ ),
    .X(\alu/_0851_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1734_  (.A(\alu/_0850_ ),
    .B(\alu/_0851_ ),
    .Y(\alu/_0852_ ));
 sky130_fd_sc_hd__a21bo_1 \alu/_1735_  (.A1(net184),
    .A2(\alu/_0847_ ),
    .B1_N(\alu/_0852_ ),
    .X(\alu/_0853_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1736_  (.A(\alu/_0853_ ),
    .B(net201),
    .Y(\alu/_0854_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1737_  (.A0(\wAluA[19] ),
    .A1(\wAluA[20] ),
    .S(net229),
    .X(\alu/_0855_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1738_  (.A0(\alu/_0615_ ),
    .A1(\alu/_0606_ ),
    .S(net233),
    .X(\alu/_0856_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1739_  (.A(\alu/_0716_ ),
    .X(\alu/_0857_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1740_  (.A(\alu/_0856_ ),
    .B(\alu/_0857_ ),
    .Y(\alu/_0858_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1741_  (.A1(\alu/_0826_ ),
    .A2(\alu/_0855_ ),
    .B1(\alu/_0858_ ),
    .Y(\alu/_0859_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1742_  (.A0(\wAluA[21] ),
    .A1(net193),
    .S(net230),
    .X(\alu/_0860_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1743_  (.A0(\wAluA[23] ),
    .A1(\wAluA[24] ),
    .S(net232),
    .X(\alu/_0861_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1744_  (.A0(\alu/_0860_ ),
    .A1(\alu/_0861_ ),
    .S(net216),
    .X(\alu/_0862_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1745_  (.A(\alu/_0862_ ),
    .B(net183),
    .Y(\alu/_0863_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1746_  (.A1(net183),
    .A2(\alu/_0859_ ),
    .B1(\alu/_0863_ ),
    .Y(\alu/_0864_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1747_  (.A(\alu/_0864_ ),
    .B(\alu/_0720_ ),
    .Y(\alu/_0865_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1748_  (.A(\alu/_0854_ ),
    .B(\alu/_0865_ ),
    .Y(\alu/_0866_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1749_  (.A(\alu/_0736_ ),
    .B(\alu/_0730_ ),
    .Y(\alu/_0867_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1750_  (.A(\alu/_0867_ ),
    .Y(\alu/_0868_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1751_  (.A(\alu/_0866_ ),
    .B(\alu/_0868_ ),
    .Y(\alu/_0869_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1752_  (.A(\alu/_0851_ ),
    .X(\alu/_0870_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1753_  (.A(net216),
    .B(net192),
    .Y(\alu/_0871_ ));
 sky130_fd_sc_hd__and2_1 \alu/_1754_  (.A(\alu/_0846_ ),
    .B(\alu/_0871_ ),
    .X(\alu/_0872_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1755_  (.A1(\alu/_0870_ ),
    .A2(\alu/_0872_ ),
    .B1(\alu/_0852_ ),
    .Y(\alu/_0873_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1756_  (.A(\alu/_0873_ ),
    .B(net201),
    .Y(\alu/_0874_ ));
 sky130_fd_sc_hd__and3_1 \alu/_1757_  (.A(\alu/_0835_ ),
    .B(\wFunct3_aluIn[0] ),
    .C(\alu/_0730_ ),
    .X(\alu/_0875_ ));
 sky130_fd_sc_hd__clkinvlp_2 \alu/_1758_  (.A(\alu/_0875_ ),
    .Y(\alu/_0876_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1759_  (.A(\alu/_0876_ ),
    .X(\alu/_0877_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1760_  (.A1(\alu/_0865_ ),
    .A2(\alu/_0874_ ),
    .B1(\alu/_0877_ ),
    .X(\alu/_0878_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1761_  (.A(\alu/_0548_ ),
    .X(\alu/_0879_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1762_  (.A(\alu/_0879_ ),
    .X(\alu/_0880_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1763_  (.A1(\alu/_0869_ ),
    .A2(\alu/_0878_ ),
    .B1(\alu/_0880_ ),
    .X(\alu/_0881_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1764_  (.A(net191),
    .B(net209),
    .Y(\alu/_0882_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1765_  (.A(\alu/_0746_ ),
    .X(\alu/_0883_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1766_  (.A(\alu/_0691_ ),
    .B(net191),
    .Y(\alu/_0884_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1767_  (.A(\alu/_0884_ ),
    .B(\alu/_0057_ ),
    .Y(\alu/_0885_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1768_  (.A(\alu/_0885_ ),
    .B(\alu/_0716_ ),
    .Y(\alu/_0886_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1769_  (.A(\alu/_0886_ ),
    .Y(\alu/_0887_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1770_  (.A(\alu/_0704_ ),
    .X(\alu/_0888_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1771_  (.A(\alu/_0887_ ),
    .B(\alu/_0888_ ),
    .Y(\alu/_0889_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1772_  (.A(net198),
    .B(\alu/_0889_ ),
    .Y(\alu/_0890_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1773_  (.A(\alu/_0883_ ),
    .B(\alu/_0890_ ),
    .Y(\alu/_0891_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1774_  (.A(\alu/_0650_ ),
    .B(\alu/_0730_ ),
    .Y(\alu/_0892_ ));
 sky130_fd_sc_hd__clkbuf_4 \alu/_1775_  (.A(\alu/_0892_ ),
    .X(\alu/_0893_ ));
 sky130_fd_sc_hd__o22a_1 \alu/_1776_  (.A1(\alu/_0121_ ),
    .A2(\alu/_0741_ ),
    .B1(\alu/_0132_ ),
    .B2(\alu/_0893_ ),
    .X(\alu/_0894_ ));
 sky130_fd_sc_hd__and3_1 \alu/_1777_  (.A(\alu/_0835_ ),
    .B(\alu/_0735_ ),
    .C(\alu/_0744_ ),
    .X(\alu/_0895_ ));
 sky130_fd_sc_hd__clkbuf_4 \alu/_1778_  (.A(\alu/_0895_ ),
    .X(\alu/_0896_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1779_  (.A(\alu/_0751_ ),
    .B(\alu/_0132_ ),
    .X(\alu/_0897_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1780_  (.A(\alu/_0650_ ),
    .B(\alu/_0744_ ),
    .Y(\alu/_0898_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1781_  (.A(\alu/_0898_ ),
    .Y(\alu/_0899_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1782_  (.A(\alu/_0132_ ),
    .B(\alu/_0057_ ),
    .Y(\alu/_0900_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1783_  (.A(\alu/_0057_ ),
    .B(\alu/_0132_ ),
    .X(\alu/_0901_ ));
 sky130_fd_sc_hd__and3_1 \alu/_1784_  (.A(\alu/_0899_ ),
    .B(\alu/_0900_ ),
    .C(\alu/_0901_ ),
    .X(\alu/_0902_ ));
 sky130_fd_sc_hd__a31oi_1 \alu/_1785_  (.A1(\alu/_0752_ ),
    .A2(\alu/_0896_ ),
    .A3(\alu/_0897_ ),
    .B1(\alu/_0902_ ),
    .Y(\alu/_0903_ ));
 sky130_fd_sc_hd__o2111a_1 \alu/_1786_  (.A1(\alu/_0882_ ),
    .A2(\alu/_0838_ ),
    .B1(\alu/_0891_ ),
    .C1(\alu/_0894_ ),
    .D1(\alu/_0903_ ),
    .X(\alu/_0904_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1787_  (.A0(\alu/_0291_ ),
    .A1(\alu/_0429_ ),
    .S(net222),
    .X(\alu/_0905_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1788_  (.A0(\alu/_0397_ ),
    .A1(\alu/_0507_ ),
    .S(net222),
    .X(\alu/_0906_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1789_  (.A0(\alu/_0905_ ),
    .A1(\alu/_0906_ ),
    .S(net208),
    .X(\alu/_0907_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1790_  (.A0(\alu/_0502_ ),
    .A1(\alu/_0520_ ),
    .S(net222),
    .X(\alu/_0908_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1791_  (.A0(\alu/_0516_ ),
    .A1(\alu/_0656_ ),
    .S(net225),
    .X(\alu/_0909_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1792_  (.A0(\alu/_0908_ ),
    .A1(\alu/_0909_ ),
    .S(net213),
    .X(\alu/_0910_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1793_  (.A0(\alu/_0907_ ),
    .A1(\alu/_0910_ ),
    .S(net178),
    .X(\alu/_0911_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1794_  (.A(\alu/_0732_ ),
    .Y(\alu/_0912_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1795_  (.A(\alu/_0912_ ),
    .X(\alu/_0913_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1796_  (.A0(\wAluA[7] ),
    .A1(\wAluA[8] ),
    .S(net227),
    .X(\alu/_0914_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1797_  (.A0(\alu/_0540_ ),
    .A1(\alu/_0528_ ),
    .S(net225),
    .X(\alu/_0915_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1798_  (.A(\alu/_0915_ ),
    .B(\alu/_0823_ ),
    .Y(\alu/_0916_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1799_  (.A1(\alu/_0823_ ),
    .A2(\alu/_0914_ ),
    .B1(\alu/_0916_ ),
    .Y(\alu/_0917_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1800_  (.A(\alu/_0692_ ),
    .B(\wAluA[3] ),
    .Y(\alu/_0918_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_1801_  (.A1(\alu/_0692_ ),
    .A2(\alu/_0546_ ),
    .B1(\alu/_0918_ ),
    .X(\alu/_0919_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1802_  (.A(net227),
    .B(\wAluA[2] ),
    .Y(\alu/_0920_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_1803_  (.A1(\alu/_0884_ ),
    .A2(\alu/_0920_ ),
    .A3(\alu/_0826_ ),
    .B1(net179),
    .X(\alu/_0921_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1804_  (.A1(net211),
    .A2(\alu/_0919_ ),
    .B1(\alu/_0921_ ),
    .X(\alu/_0922_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_1805_  (.A1(\alu/_0705_ ),
    .A2(\alu/_0917_ ),
    .B1(\alu/_0711_ ),
    .C1(\alu/_0922_ ),
    .X(\alu/_0923_ ));
 sky130_fd_sc_hd__a211o_1 \alu/_1806_  (.A1(\alu/_0911_ ),
    .A2(net196),
    .B1(\alu/_0913_ ),
    .C1(\alu/_0923_ ),
    .X(\alu/_0924_ ));
 sky130_fd_sc_hd__nand3_4 \alu/_1807_  (.A(\alu/_0881_ ),
    .B(\alu/_0904_ ),
    .C(\alu/_0924_ ),
    .Y(\wAluOut[1] ));
 sky130_fd_sc_hd__nand2_1 \alu/_1808_  (.A(\alu/_0196_ ),
    .B(\alu/_0217_ ),
    .Y(\alu/_0925_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1809_  (.A(\wAluA[2] ),
    .B(net175),
    .Y(\alu/_0926_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1810_  (.A(\alu/_0925_ ),
    .B(\alu/_0926_ ),
    .Y(\alu/_0927_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1811_  (.A(\alu/_0892_ ),
    .X(\alu/_0928_ ));
 sky130_fd_sc_hd__clkbuf_4 \alu/_1812_  (.A(\alu/_0928_ ),
    .X(\alu/_0929_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1813_  (.A(\alu/_0739_ ),
    .Y(\alu/_0930_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1814_  (.A(\alu/_0926_ ),
    .Y(\alu/_0931_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1815_  (.A(\alu/_0837_ ),
    .Y(\alu/_0932_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1816_  (.A(\alu/_0932_ ),
    .X(\alu/_0933_ ));
 sky130_fd_sc_hd__a22o_1 \alu/_1817_  (.A1(\alu/_0930_ ),
    .A2(\alu/_0931_ ),
    .B1(\alu/_0925_ ),
    .B2(\alu/_0933_ ),
    .X(\alu/_0934_ ));
 sky130_fd_sc_hd__buf_6 \alu/_1818_  (.A(\alu/_0895_ ),
    .X(\alu/_0935_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1819_  (.A(\alu/_0754_ ),
    .B(\alu/_0927_ ),
    .Y(\alu/_0936_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1820_  (.A(\alu/_0927_ ),
    .B(\alu/_0754_ ),
    .X(\alu/_0937_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1821_  (.A1(\alu/_0057_ ),
    .A2(\alu/_0882_ ),
    .B1(\alu/_0121_ ),
    .Y(\alu/_0938_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_1822_  (.A1(\alu/_0238_ ),
    .A2(\alu/_0938_ ),
    .B1(\alu/_0899_ ),
    .X(\alu/_0939_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1823_  (.A(\alu/_0938_ ),
    .B(\alu/_0238_ ),
    .Y(\alu/_0940_ ));
 sky130_fd_sc_hd__a32o_1 \alu/_1824_  (.A1(\alu/_0935_ ),
    .A2(\alu/_0936_ ),
    .A3(\alu/_0937_ ),
    .B1(\alu/_0939_ ),
    .B2(\alu/_0940_ ),
    .X(\alu/_0941_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1825_  (.A(\alu/_0934_ ),
    .B(\alu/_0941_ ),
    .Y(\alu/_0942_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1826_  (.A0(\alu/_0824_ ),
    .A1(\alu/_0819_ ),
    .S(net217),
    .X(\alu/_0943_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1827_  (.A0(\alu/_0820_ ),
    .A1(\alu/_0806_ ),
    .S(net214),
    .X(\alu/_0944_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1828_  (.A0(\alu/_0943_ ),
    .A1(\alu/_0944_ ),
    .S(net183),
    .X(\alu/_0945_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1829_  (.A(\alu/_0709_ ),
    .X(\alu/_0946_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1830_  (.A(\alu/_0946_ ),
    .X(\alu/_0947_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1831_  (.A(\alu/_0945_ ),
    .B(\alu/_0947_ ),
    .Y(\alu/_0948_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1832_  (.A(\alu/_0810_ ),
    .B(\alu/_0715_ ),
    .Y(\alu/_0949_ ));
 sky130_fd_sc_hd__and2_1 \alu/_1833_  (.A(\alu/_0949_ ),
    .B(\alu/_0871_ ),
    .X(\alu/_0950_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1834_  (.A0(\alu/_0807_ ),
    .A1(\alu/_0813_ ),
    .S(net218),
    .X(\alu/_0951_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1835_  (.A(\alu/_0951_ ),
    .B(\alu/_0870_ ),
    .Y(\alu/_0952_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1836_  (.A1(\alu/_0870_ ),
    .A2(\alu/_0950_ ),
    .B1(\alu/_0952_ ),
    .Y(\alu/_0953_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1837_  (.A(\alu/_0953_ ),
    .B(net205),
    .Y(\alu/_0954_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1838_  (.A(\alu/_0948_ ),
    .B(\alu/_0954_ ),
    .Y(\alu/_0955_ ));
 sky130_fd_sc_hd__buf_6 \alu/_1839_  (.A(\alu/_0875_ ),
    .X(\alu/_0956_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1840_  (.A(\alu/_0955_ ),
    .B(\alu/_0956_ ),
    .Y(\alu/_0957_ ));
 sky130_fd_sc_hd__o21ai_2 \alu/_1841_  (.A1(\alu/_0870_ ),
    .A2(\alu/_0949_ ),
    .B1(\alu/_0952_ ),
    .Y(\alu/_0958_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1842_  (.A(\alu/_0958_ ),
    .B(net205),
    .Y(\alu/_0959_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1843_  (.A(\alu/_0948_ ),
    .B(\alu/_0959_ ),
    .Y(\alu/_0960_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1844_  (.A(\alu/_0960_ ),
    .B(\alu/_0868_ ),
    .Y(\alu/_0961_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1845_  (.A(\alu/_0957_ ),
    .B(\alu/_0961_ ),
    .Y(\alu/_0962_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1846_  (.A(\alu/_0962_ ),
    .B(net173),
    .Y(\alu/_0963_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1847_  (.A0(\alu/_0723_ ),
    .A1(\alu/_0725_ ),
    .S(net209),
    .X(\alu/_0964_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1848_  (.A(\alu/_0726_ ),
    .B(\alu/_0857_ ),
    .Y(\alu/_0965_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1849_  (.A1(\alu/_0826_ ),
    .A2(\alu/_0825_ ),
    .B1(\alu/_0965_ ),
    .Y(\alu/_0966_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1850_  (.A0(\alu/_0964_ ),
    .A1(\alu/_0966_ ),
    .S(net177),
    .X(\alu/_0967_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_1851_  (.A(\alu/_0967_ ),
    .B(net195),
    .C(\alu/_0803_ ),
    .Y(\alu/_0968_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1852_  (.A0(\alu/_0706_ ),
    .A1(\alu/_0712_ ),
    .S(\alu/_0857_ ),
    .X(\alu/_0969_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1853_  (.A(net202),
    .B(\alu/_0731_ ),
    .Y(\alu/_0970_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1854_  (.A(\alu/_0970_ ),
    .Y(\alu/_0971_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1855_  (.A(\alu/_0707_ ),
    .B(\alu/_0857_ ),
    .Y(\alu/_0972_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1856_  (.A1(\alu/_0826_ ),
    .A2(\alu/_0722_ ),
    .B1(\alu/_0972_ ),
    .Y(\alu/_0973_ ));
 sky130_fd_sc_hd__and2_1 \alu/_1857_  (.A(\alu/_0973_ ),
    .B(net177),
    .X(\alu/_0974_ ));
 sky130_fd_sc_hd__a211o_1 \alu/_1858_  (.A1(\alu/_0969_ ),
    .A2(\alu/_0818_ ),
    .B1(\alu/_0971_ ),
    .C1(\alu/_0974_ ),
    .X(\alu/_0975_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1859_  (.A(\alu/_0745_ ),
    .X(\alu/_0976_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1860_  (.A(net196),
    .B(\alu/_0976_ ),
    .Y(\alu/_0977_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1861_  (.A1(net227),
    .A2(\alu/_0196_ ),
    .B1(\alu/_0713_ ),
    .Y(\alu/_0978_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_1862_  (.A1(net210),
    .A2(\alu/_0978_ ),
    .B1(\alu/_0694_ ),
    .X(\alu/_0979_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1863_  (.A(\alu/_0979_ ),
    .B(\alu/_0817_ ),
    .Y(\alu/_0980_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1864_  (.A(\alu/_0980_ ),
    .Y(\alu/_0981_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1865_  (.A(\alu/_0977_ ),
    .B(\alu/_0981_ ),
    .Y(\alu/_0982_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_1866_  (.A1(\alu/_0968_ ),
    .A2(\alu/_0975_ ),
    .A3(\alu/_0982_ ),
    .B1(net173),
    .X(\alu/_0983_ ));
 sky130_fd_sc_hd__o2111ai_4 \alu/_1867_  (.A1(\alu/_0927_ ),
    .A2(\alu/_0929_ ),
    .B1(\alu/_0942_ ),
    .C1(\alu/_0963_ ),
    .D1(\alu/_0983_ ),
    .Y(\wAluOut[2] ));
 sky130_fd_sc_hd__nand2_1 \alu/_1868_  (.A(\alu/_0905_ ),
    .B(net208),
    .Y(\alu/_0984_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1869_  (.A1(net208),
    .A2(\alu/_0914_ ),
    .B1(\alu/_0984_ ),
    .Y(\alu/_0985_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1870_  (.A(\alu/_0831_ ),
    .X(\alu/_0986_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1871_  (.A1(\alu/_0915_ ),
    .A2(net208),
    .B1(net175),
    .X(\alu/_0987_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1872_  (.A1(\alu/_0823_ ),
    .A2(\alu/_0919_ ),
    .B1(\alu/_0987_ ),
    .X(\alu/_0988_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_1873_  (.A1(\alu/_0705_ ),
    .A2(\alu/_0985_ ),
    .B1(\alu/_0986_ ),
    .C1(\alu/_0988_ ),
    .X(\alu/_0989_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1874_  (.A0(\alu/_0906_ ),
    .A1(\alu/_0908_ ),
    .S(net209),
    .X(\alu/_0990_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1875_  (.A0(\alu/_0909_ ),
    .A1(\alu/_0856_ ),
    .S(net209),
    .X(\alu/_0991_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1876_  (.A0(\alu/_0990_ ),
    .A1(\alu/_0991_ ),
    .S(net177),
    .X(\alu/_0992_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1877_  (.A1(\alu/_0992_ ),
    .A2(net196),
    .B1(\alu/_0913_ ),
    .X(\alu/_0993_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1878_  (.A(\alu/_0143_ ),
    .B(\alu/_0164_ ),
    .Y(\alu/_0994_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1879_  (.A(\wAluA[3] ),
    .B(net197),
    .Y(\alu/_0995_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1880_  (.A(\alu/_0994_ ),
    .B(\alu/_0995_ ),
    .Y(\alu/_0996_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_1881_  (.A1(\alu/_0940_ ),
    .A2(\alu/_0926_ ),
    .B1(\alu/_0996_ ),
    .Y(\alu/_0997_ ));
 sky130_fd_sc_hd__or3b_1 \alu/_1882_  (.A(\alu/_0185_ ),
    .B(\alu/_0931_ ),
    .C_N(\alu/_0940_ ),
    .X(\alu/_0998_ ));
 sky130_fd_sc_hd__or3b_2 \alu/_1883_  (.A(\alu/_0898_ ),
    .B(\alu/_0997_ ),
    .C_N(\alu/_0998_ ),
    .X(\alu/_0999_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1884_  (.A(net217),
    .B(\alu/_0855_ ),
    .X(\alu/_1000_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1885_  (.A1(\alu/_0822_ ),
    .A2(\alu/_0860_ ),
    .B1(\alu/_1000_ ),
    .Y(\alu/_1001_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1886_  (.A0(\alu/_0848_ ),
    .A1(\alu/_0861_ ),
    .S(\alu/_0715_ ),
    .X(\alu/_1002_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1887_  (.A(\alu/_1002_ ),
    .B(net184),
    .Y(\alu/_1003_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1888_  (.A1(net184),
    .A2(\alu/_1001_ ),
    .B1(\alu/_1003_ ),
    .Y(\alu/_1004_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1889_  (.A(\alu/_1004_ ),
    .B(\alu/_0710_ ),
    .Y(\alu/_1005_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1890_  (.A(\alu/_0842_ ),
    .B(\alu/_0845_ ),
    .Y(\alu/_1006_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1891_  (.A0(\alu/_0849_ ),
    .A1(\alu/_0844_ ),
    .S(net216),
    .X(\alu/_1007_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1892_  (.A(\alu/_1007_ ),
    .B(\alu/_0704_ ),
    .Y(\alu/_1008_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1893_  (.A1(\alu/_0851_ ),
    .A2(\alu/_1006_ ),
    .B1(\alu/_1008_ ),
    .Y(\alu/_1009_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1894_  (.A(\alu/_1009_ ),
    .B(net202),
    .Y(\alu/_1010_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1895_  (.A1(\alu/_1005_ ),
    .A2(\alu/_1010_ ),
    .B1(\alu/_0867_ ),
    .X(\alu/_1011_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1896_  (.A(net185),
    .B(\wAluA[31] ),
    .Y(\alu/_1012_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1897_  (.A(\alu/_1008_ ),
    .B(\alu/_1012_ ),
    .Y(\alu/_1013_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1898_  (.A(\alu/_1013_ ),
    .B(net201),
    .Y(\alu/_1014_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1899_  (.A1(\alu/_1005_ ),
    .A2(\alu/_1014_ ),
    .B1(\alu/_0876_ ),
    .X(\alu/_1015_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1900_  (.A(\alu/_1011_ ),
    .B(\alu/_1015_ ),
    .Y(\alu/_1016_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1901_  (.A(\alu/_1016_ ),
    .B(net173),
    .Y(\alu/_1017_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1902_  (.A(\alu/_0746_ ),
    .X(\alu/_1018_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1903_  (.A(\alu/_0918_ ),
    .B(\alu/_0920_ ),
    .Y(\alu/_1019_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1904_  (.A0(\alu/_1019_ ),
    .A1(\alu/_0885_ ),
    .S(net210),
    .X(\alu/_1020_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1905_  (.A(\alu/_1020_ ),
    .B(\alu/_0888_ ),
    .Y(\alu/_1021_ ));
 sky130_fd_sc_hd__nor2_2 \alu/_1906_  (.A(net204),
    .B(\alu/_1021_ ),
    .Y(\alu/_1022_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1907_  (.A(\alu/_0996_ ),
    .B(\alu/_0929_ ),
    .Y(\alu/_1023_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1908_  (.A(\alu/_0936_ ),
    .B(\alu/_0227_ ),
    .Y(\alu/_1024_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1909_  (.A(\alu/_0996_ ),
    .B(\alu/_1024_ ),
    .X(\alu/_1025_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1910_  (.A(\alu/_1024_ ),
    .B(\alu/_0996_ ),
    .Y(\alu/_1026_ ));
 sky130_fd_sc_hd__and3_1 \alu/_1911_  (.A(\alu/_1025_ ),
    .B(\alu/_0935_ ),
    .C(\alu/_1026_ ),
    .X(\alu/_1027_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1912_  (.A(\alu/_0995_ ),
    .Y(\alu/_1028_ ));
 sky130_fd_sc_hd__a22o_1 \alu/_1913_  (.A1(\alu/_0930_ ),
    .A2(\alu/_1028_ ),
    .B1(\alu/_0994_ ),
    .B2(\alu/_0933_ ),
    .X(\alu/_1029_ ));
 sky130_fd_sc_hd__a2111oi_2 \alu/_1914_  (.A1(\alu/_1018_ ),
    .A2(\alu/_1022_ ),
    .B1(\alu/_1023_ ),
    .C1(\alu/_1027_ ),
    .D1(\alu/_1029_ ),
    .Y(\alu/_1030_ ));
 sky130_fd_sc_hd__o2111ai_4 \alu/_1915_  (.A1(\alu/_0989_ ),
    .A2(\alu/_0993_ ),
    .B1(\alu/_0999_ ),
    .C1(\alu/_1017_ ),
    .D1(\alu/_1030_ ),
    .Y(\wAluOut[3] ));
 sky130_fd_sc_hd__mux2_1 \alu/_1916_  (.A0(\wAluA[4] ),
    .A1(\wAluA[3] ),
    .S(net226),
    .X(\alu/_1031_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1917_  (.A0(\alu/_1031_ ),
    .A1(\alu/_0978_ ),
    .S(net210),
    .X(\alu/_1032_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1918_  (.A0(\alu/_1032_ ),
    .A1(\alu/_0696_ ),
    .S(net179),
    .X(\alu/_1033_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1919_  (.A(\alu/_1033_ ),
    .B(\alu/_0986_ ),
    .Y(\alu/_1034_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1920_  (.A1(net173),
    .A2(\wAluA[4] ),
    .B1(\alu/_0933_ ),
    .Y(\alu/_1035_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1921_  (.A(net170),
    .B(\wAluA[4] ),
    .Y(\alu/_1036_ ));
 sky130_fd_sc_hd__o22a_1 \alu/_1922_  (.A1(\alu/_1036_ ),
    .A2(\alu/_0741_ ),
    .B1(\alu/_0551_ ),
    .B2(\alu/_0929_ ),
    .X(\alu/_1037_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1923_  (.A(\alu/_0727_ ),
    .B(\alu/_0888_ ),
    .Y(\alu/_1038_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1924_  (.A1(\alu/_0888_ ),
    .A2(\alu/_0828_ ),
    .B1(\alu/_1038_ ),
    .Y(\alu/_1039_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1925_  (.A(\alu/_0724_ ),
    .B(net175),
    .Y(\alu/_1040_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1926_  (.A1(net175),
    .A2(\alu/_0708_ ),
    .B1(\alu/_1040_ ),
    .Y(\alu/_1041_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1927_  (.A0(\alu/_1039_ ),
    .A1(\alu/_1041_ ),
    .S(\alu/_0946_ ),
    .X(\alu/_1042_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1928_  (.A(\alu/_1042_ ),
    .B(\alu/_0733_ ),
    .Y(\alu/_1043_ ));
 sky130_fd_sc_hd__o2111a_1 \alu/_1929_  (.A1(\alu/_0747_ ),
    .A2(\alu/_1034_ ),
    .B1(\alu/_1035_ ),
    .C1(\alu/_1037_ ),
    .D1(\alu/_1043_ ),
    .X(\alu/_1044_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1930_  (.A(\alu/_0814_ ),
    .B(\alu/_0816_ ),
    .Y(\alu/_1045_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1931_  (.A0(\alu/_0821_ ),
    .A1(\alu/_0808_ ),
    .S(net183),
    .X(\alu/_1046_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_1932_  (.A(\alu/_0710_ ),
    .X(\alu/_1047_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1933_  (.A(\alu/_1046_ ),
    .B(\alu/_1047_ ),
    .Y(\alu/_1048_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_1934_  (.A1(\alu/_0947_ ),
    .A2(\alu/_1045_ ),
    .B1(\alu/_1048_ ),
    .X(\alu/_1049_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1935_  (.A(\alu/_1045_ ),
    .B(\alu/_1012_ ),
    .Y(\alu/_1050_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1936_  (.A(\alu/_1050_ ),
    .B(net202),
    .Y(\alu/_1051_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1937_  (.A1(\alu/_1048_ ),
    .A2(\alu/_1051_ ),
    .B1(\alu/_0877_ ),
    .X(\alu/_1052_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1938_  (.A1(\alu/_0867_ ),
    .A2(\alu/_1049_ ),
    .B1(\alu/_1052_ ),
    .Y(\alu/_1053_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1939_  (.A(\alu/_1053_ ),
    .B(net170),
    .Y(\alu/_1054_ ));
 sky130_fd_sc_hd__clkbuf_4 \alu/_1940_  (.A(\alu/_0896_ ),
    .X(\alu/_1055_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1941_  (.A(\alu/_0758_ ),
    .Y(\alu/_1056_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1942_  (.A(\alu/_0550_ ),
    .B(\alu/_1056_ ),
    .Y(\alu/_1057_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1943_  (.A(\alu/_1057_ ),
    .Y(\alu/_1058_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1944_  (.A(\alu/_1056_ ),
    .B(\alu/_0550_ ),
    .Y(\alu/_1059_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1945_  (.A(\alu/_0899_ ),
    .X(\alu/_1060_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1946_  (.A(\alu/_0996_ ),
    .B(\alu/_0927_ ),
    .Y(\alu/_1061_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1947_  (.A(\alu/_1061_ ),
    .B(\alu/_0938_ ),
    .Y(\alu/_1062_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_1948_  (.A1(\alu/_0994_ ),
    .A2(\alu/_0931_ ),
    .B1(\alu/_1028_ ),
    .Y(\alu/_1063_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1949_  (.A(\alu/_1062_ ),
    .B(\alu/_1063_ ),
    .Y(\alu/_1064_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1950_  (.A(\alu/_0550_ ),
    .B(\alu/_1064_ ),
    .X(\alu/_1065_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1951_  (.A(\alu/_1064_ ),
    .B(\alu/_0550_ ),
    .Y(\alu/_1066_ ));
 sky130_fd_sc_hd__and3_1 \alu/_1952_  (.A(\alu/_1060_ ),
    .B(\alu/_1065_ ),
    .C(\alu/_1066_ ),
    .X(\alu/_1067_ ));
 sky130_fd_sc_hd__a31oi_2 \alu/_1953_  (.A1(\alu/_1055_ ),
    .A2(\alu/_1058_ ),
    .A3(\alu/_1059_ ),
    .B1(\alu/_1067_ ),
    .Y(\alu/_1068_ ));
 sky130_fd_sc_hd__nand3_4 \alu/_1954_  (.A(\alu/_1044_ ),
    .B(\alu/_1054_ ),
    .C(\alu/_1068_ ),
    .Y(\wAluOut[4] ));
 sky130_fd_sc_hd__nand2_1 \alu/_1955_  (.A(\alu/_1058_ ),
    .B(\alu/_0549_ ),
    .Y(\alu/_1069_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1956_  (.A(\alu/_0545_ ),
    .B(\alu/_1069_ ),
    .X(\alu/_1070_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1957_  (.A(\alu/_1069_ ),
    .B(\alu/_0545_ ),
    .Y(\alu/_1071_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1958_  (.A(\alu/_1066_ ),
    .B(\alu/_1036_ ),
    .Y(\alu/_1072_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1959_  (.A(\alu/_0544_ ),
    .B(\alu/_1072_ ),
    .X(\alu/_1073_ ));
 sky130_fd_sc_hd__clkbuf_4 \alu/_1960_  (.A(\alu/_0898_ ),
    .X(\alu/_1074_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_1961_  (.A1(\alu/_1072_ ),
    .A2(\alu/_0544_ ),
    .B1(\alu/_1074_ ),
    .Y(\alu/_1075_ ));
 sky130_fd_sc_hd__a32o_1 \alu/_1962_  (.A1(\alu/_1070_ ),
    .A2(\alu/_0896_ ),
    .A3(\alu/_1071_ ),
    .B1(\alu/_1073_ ),
    .B2(\alu/_1075_ ),
    .X(\alu/_1076_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1963_  (.A0(\alu/_0907_ ),
    .A1(\alu/_0917_ ),
    .S(\alu/_0888_ ),
    .X(\alu/_1077_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1964_  (.A(\alu/_1077_ ),
    .B(\alu/_0721_ ),
    .Y(\alu/_1078_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1965_  (.A0(\alu/_0910_ ),
    .A1(\alu/_0859_ ),
    .S(net177),
    .X(\alu/_1079_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1966_  (.A(\alu/_1079_ ),
    .B(net195),
    .Y(\alu/_1080_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1967_  (.A(\wAluA[5] ),
    .B(\wAluB[5] ),
    .Y(\alu/_1081_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1968_  (.A(\wAluA[5] ),
    .B(\wAluB[5] ),
    .Y(\alu/_1082_ ));
 sky130_fd_sc_hd__buf_2 \alu/_1969_  (.A(\alu/_0739_ ),
    .X(\alu/_1083_ ));
 sky130_fd_sc_hd__o22a_1 \alu/_1970_  (.A1(\alu/_1082_ ),
    .A2(\alu/_1083_ ),
    .B1(\alu/_0545_ ),
    .B2(\alu/_0928_ ),
    .X(\alu/_1084_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1971_  (.A0(\wAluA[5] ),
    .A1(\wAluA[4] ),
    .S(net227),
    .X(\alu/_1085_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1972_  (.A(\alu/_0845_ ),
    .B(\alu/_1019_ ),
    .X(\alu/_1086_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1973_  (.A1(net211),
    .A2(\alu/_1085_ ),
    .B1(\alu/_1086_ ),
    .Y(\alu/_1087_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1974_  (.A(\alu/_0887_ ),
    .B(net180),
    .Y(\alu/_1088_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1975_  (.A1(net179),
    .A2(\alu/_1087_ ),
    .B1(\alu/_1088_ ),
    .Y(\alu/_1089_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1976_  (.A(\alu/_1089_ ),
    .B(\alu/_0946_ ),
    .Y(\alu/_1090_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1977_  (.A(\alu/_0747_ ),
    .B(\alu/_1090_ ),
    .X(\alu/_1091_ ));
 sky130_fd_sc_hd__o211ai_1 \alu/_1978_  (.A1(\alu/_1081_ ),
    .A2(\alu/_0838_ ),
    .B1(\alu/_1084_ ),
    .C1(\alu/_1091_ ),
    .Y(\alu/_1092_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_1979_  (.A1(\alu/_0733_ ),
    .A2(\alu/_1078_ ),
    .A3(\alu/_1080_ ),
    .B1(\alu/_1092_ ),
    .X(\alu/_1093_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_1980_  (.A(\alu/_1076_ ),
    .B(\alu/_1093_ ),
    .Y(\alu/_1094_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_1981_  (.A0(\alu/_0850_ ),
    .A1(\alu/_0862_ ),
    .S(\alu/_0704_ ),
    .X(\alu/_1095_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1982_  (.A(\alu/_1095_ ),
    .B(\alu/_1047_ ),
    .Y(\alu/_1096_ ));
 sky130_fd_sc_hd__and2_1 \alu/_1983_  (.A(\alu/_0871_ ),
    .B(\alu/_1012_ ),
    .X(\alu/_1097_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1984_  (.A1(net184),
    .A2(\alu/_0846_ ),
    .B1(\alu/_1097_ ),
    .Y(\alu/_1098_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1985_  (.A(\alu/_1098_ ),
    .B(net201),
    .Y(\alu/_1099_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_1986_  (.A1(\alu/_1096_ ),
    .A2(\alu/_1099_ ),
    .B1(\alu/_0877_ ),
    .X(\alu/_1100_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1987_  (.A(\alu/_0847_ ),
    .B(\alu/_0851_ ),
    .Y(\alu/_1101_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1988_  (.A1(\alu/_0832_ ),
    .A2(\alu/_1101_ ),
    .B1(\alu/_1096_ ),
    .Y(\alu/_1102_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1989_  (.A(\alu/_1102_ ),
    .B(\alu/_0868_ ),
    .Y(\alu/_1103_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1990_  (.A(\alu/_1100_ ),
    .B(\alu/_1103_ ),
    .Y(\alu/_1104_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1991_  (.A(\alu/_1104_ ),
    .B(net170),
    .Y(\alu/_1105_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_1992_  (.A(\alu/_1094_ ),
    .B(\alu/_1105_ ),
    .Y(\wAluOut[5] ));
 sky130_fd_sc_hd__a21o_1 \alu/_1993_  (.A1(\alu/_1036_ ),
    .A2(\alu/_1082_ ),
    .B1(\alu/_1081_ ),
    .X(\alu/_1106_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_1994_  (.A1(\alu/_0545_ ),
    .A2(\alu/_1066_ ),
    .B1(\alu/_1106_ ),
    .Y(\alu/_1107_ ));
 sky130_fd_sc_hd__or2_1 \alu/_1995_  (.A(\alu/_0532_ ),
    .B(\alu/_1107_ ),
    .X(\alu/_1108_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1996_  (.A(\alu/_1107_ ),
    .B(\alu/_0532_ ),
    .Y(\alu/_1109_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1997_  (.A(\alu/_1108_ ),
    .B(\alu/_1109_ ),
    .Y(\alu/_1110_ ));
 sky130_fd_sc_hd__inv_2 \alu/_1998_  (.A(\alu/_0532_ ),
    .Y(\alu/_1111_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_1999_  (.A(\alu/_1071_ ),
    .B(\alu/_0542_ ),
    .Y(\alu/_1112_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2000_  (.A(\alu/_1111_ ),
    .B(\alu/_1112_ ),
    .X(\alu/_1113_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_2001_  (.A(\alu/_0935_ ),
    .X(\alu/_1114_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2002_  (.A(\alu/_1112_ ),
    .B(\alu/_1111_ ),
    .Y(\alu/_1115_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2003_  (.A(\alu/_1113_ ),
    .B(\alu/_1114_ ),
    .C(\alu/_1115_ ),
    .Y(\alu/_1116_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2004_  (.A0(\alu/_0944_ ),
    .A1(\alu/_0951_ ),
    .S(net186),
    .X(\alu/_1117_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2005_  (.A(\alu/_1117_ ),
    .B(\alu/_0720_ ),
    .Y(\alu/_1118_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2006_  (.A(net188),
    .B(\alu/_0949_ ),
    .X(\alu/_1119_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2007_  (.A(\alu/_1119_ ),
    .B(\alu/_1097_ ),
    .Y(\alu/_1120_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2008_  (.A(\alu/_1120_ ),
    .B(net205),
    .Y(\alu/_1121_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2009_  (.A1(\alu/_1118_ ),
    .A2(\alu/_1121_ ),
    .B1(\alu/_0877_ ),
    .X(\alu/_1122_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2010_  (.A1(\alu/_0986_ ),
    .A2(\alu/_1119_ ),
    .B1(\alu/_1118_ ),
    .Y(\alu/_1123_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2011_  (.A(\alu/_1123_ ),
    .B(\alu/_0868_ ),
    .Y(\alu/_1124_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_2012_  (.A(\alu/_1122_ ),
    .B(\alu/_1124_ ),
    .Y(\alu/_1125_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2013_  (.A(\alu/_1125_ ),
    .B(net169),
    .Y(\alu/_1126_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2014_  (.A0(\wAluA[6] ),
    .A1(\wAluA[5] ),
    .S(net226),
    .X(\alu/_1127_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2015_  (.A(net210),
    .B(\alu/_1127_ ),
    .X(\alu/_1128_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2016_  (.A1(\alu/_0857_ ),
    .A2(\alu/_1031_ ),
    .B1(\alu/_1128_ ),
    .Y(\alu/_1129_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2017_  (.A(\alu/_0979_ ),
    .B(net180),
    .Y(\alu/_1130_ ));
 sky130_fd_sc_hd__o21ai_2 \alu/_2018_  (.A1(net179),
    .A2(\alu/_1129_ ),
    .B1(\alu/_1130_ ),
    .Y(\alu/_1131_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2019_  (.A(\alu/_1131_ ),
    .B(\alu/_0720_ ),
    .Y(\alu/_1132_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2020_  (.A(\wAluA[6] ),
    .B(\wAluB[6] ),
    .Y(\alu/_1133_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_2021_  (.A(\alu/_0740_ ),
    .X(\alu/_1134_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_2022_  (.A(\alu/_0892_ ),
    .X(\alu/_1135_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_2023_  (.A(\alu/_0932_ ),
    .X(\alu/_1136_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2024_  (.A1(\wAluA[6] ),
    .A2(\wAluB[6] ),
    .B1(\alu/_1136_ ),
    .Y(\alu/_1137_ ));
 sky130_fd_sc_hd__o221a_1 \alu/_2025_  (.A1(\alu/_1133_ ),
    .A2(\alu/_1134_ ),
    .B1(\alu/_1111_ ),
    .B2(\alu/_1135_ ),
    .C1(\alu/_1137_ ),
    .X(\alu/_1138_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2026_  (.A(net177),
    .B(\alu/_0973_ ),
    .Y(\alu/_1139_ ));
 sky130_fd_sc_hd__a211o_1 \alu/_2027_  (.A1(\alu/_0964_ ),
    .A2(net177),
    .B1(net195),
    .C1(\alu/_1139_ ),
    .X(\alu/_1140_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2028_  (.A(net183),
    .B(\alu/_0966_ ),
    .X(\alu/_1141_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2029_  (.A1(\alu/_0818_ ),
    .A2(\alu/_0943_ ),
    .B1(\alu/_1141_ ),
    .Y(\alu/_1142_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2030_  (.A(\alu/_1142_ ),
    .B(net195),
    .Y(\alu/_1143_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2031_  (.A(\alu/_1140_ ),
    .B(\alu/_0733_ ),
    .C(\alu/_1143_ ),
    .Y(\alu/_1144_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2032_  (.A1(\alu/_0747_ ),
    .A2(\alu/_1132_ ),
    .B1(\alu/_1138_ ),
    .C1(\alu/_1144_ ),
    .X(\alu/_1145_ ));
 sky130_fd_sc_hd__o2111ai_4 \alu/_2033_  (.A1(\alu/_1074_ ),
    .A2(\alu/_1110_ ),
    .B1(\alu/_1116_ ),
    .C1(\alu/_1126_ ),
    .D1(\alu/_1145_ ),
    .Y(\wAluOut[6] ));
 sky130_fd_sc_hd__mux2_1 \alu/_2034_  (.A0(\alu/_0990_ ),
    .A1(\alu/_0985_ ),
    .S(\alu/_0817_ ),
    .X(\alu/_1146_ ));
 sky130_fd_sc_hd__and2_1 \alu/_2035_  (.A(\alu/_1146_ ),
    .B(\alu/_0711_ ),
    .X(\alu/_1147_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2036_  (.A0(\alu/_0991_ ),
    .A1(\alu/_1001_ ),
    .S(net178),
    .X(\alu/_1148_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2037_  (.A1(\alu/_1148_ ),
    .A2(net196),
    .B1(\alu/_0913_ ),
    .X(\alu/_1149_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2038_  (.A0(net190),
    .A1(\wAluA[6] ),
    .S(net227),
    .X(\alu/_1150_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2039_  (.A0(\alu/_1150_ ),
    .A1(\alu/_1085_ ),
    .S(net212),
    .X(\alu/_1151_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2040_  (.A0(\alu/_1151_ ),
    .A1(\alu/_1020_ ),
    .S(net181),
    .X(\alu/_1152_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2041_  (.A(\alu/_1152_ ),
    .B(\alu/_1047_ ),
    .Y(\alu/_1153_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2042_  (.A(net190),
    .B(\wAluB[7] ),
    .Y(\alu/_1154_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_2043_  (.A(\alu/_0739_ ),
    .X(\alu/_1155_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2044_  (.A(\alu/_0537_ ),
    .Y(\alu/_1156_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2045_  (.A1(net190),
    .A2(\wAluB[7] ),
    .B1(\alu/_1136_ ),
    .Y(\alu/_1157_ ));
 sky130_fd_sc_hd__o221a_1 \alu/_2046_  (.A1(\alu/_1154_ ),
    .A2(\alu/_1155_ ),
    .B1(\alu/_1156_ ),
    .B2(\alu/_0928_ ),
    .C1(\alu/_1157_ ),
    .X(\alu/_1158_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_2047_  (.A1(\alu/_0747_ ),
    .A2(\alu/_1153_ ),
    .B1(\alu/_1158_ ),
    .X(\alu/_1159_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2048_  (.A1(\alu/_1147_ ),
    .A2(\alu/_1149_ ),
    .B1(\alu/_1159_ ),
    .Y(\alu/_1160_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2049_  (.A(\alu/_1002_ ),
    .B(\alu/_0817_ ),
    .Y(\alu/_1161_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2050_  (.A(\alu/_1007_ ),
    .B(net184),
    .Y(\alu/_1162_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2051_  (.A(\alu/_1161_ ),
    .B(\alu/_1162_ ),
    .Y(\alu/_1163_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2052_  (.A(net201),
    .B(net192),
    .Y(\alu/_1164_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2053_  (.A(\alu/_1164_ ),
    .Y(\alu/_1165_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_2054_  (.A(\alu/_1165_ ),
    .X(\alu/_1166_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2055_  (.A1(\alu/_1163_ ),
    .A2(\alu/_0831_ ),
    .B1(\alu/_1166_ ),
    .X(\alu/_1167_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2056_  (.A(net183),
    .B(\alu/_1006_ ),
    .Y(\alu/_1168_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2057_  (.A0(\alu/_1163_ ),
    .A1(\alu/_1168_ ),
    .S(net202),
    .X(\alu/_1169_ ));
 sky130_fd_sc_hd__a22oi_1 \alu/_2058_  (.A1(\alu/_1167_ ),
    .A2(\alu/_0956_ ),
    .B1(\alu/_1169_ ),
    .B2(\alu/_0868_ ),
    .Y(\alu/_1170_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2059_  (.A(\alu/_0880_ ),
    .B(\alu/_1170_ ),
    .Y(\alu/_1171_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2060_  (.A(\alu/_1160_ ),
    .B(\alu/_1171_ ),
    .Y(\alu/_1172_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2061_  (.A(\alu/_1115_ ),
    .B(\alu/_0531_ ),
    .Y(\alu/_1173_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2062_  (.A1(\alu/_1156_ ),
    .A2(\alu/_1173_ ),
    .B1(\alu/_1114_ ),
    .Y(\alu/_1174_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2063_  (.A1(\alu/_1156_ ),
    .A2(\alu/_1173_ ),
    .B1(\alu/_1174_ ),
    .X(\alu/_1175_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2064_  (.A1(\alu/_1109_ ),
    .A2(\alu/_1133_ ),
    .B1(\alu/_1156_ ),
    .X(\alu/_1176_ ));
 sky130_fd_sc_hd__buf_2 \alu/_2065_  (.A(\alu/_0899_ ),
    .X(\alu/_1177_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2066_  (.A(\alu/_1176_ ),
    .B(\alu/_1177_ ),
    .Y(\alu/_1178_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2067_  (.A1(\alu/_1133_ ),
    .A2(\alu/_1156_ ),
    .A3(\alu/_1109_ ),
    .B1(\alu/_1178_ ),
    .X(\alu/_1179_ ));
 sky130_fd_sc_hd__nand3_4 \alu/_2068_  (.A(\alu/_1172_ ),
    .B(\alu/_1175_ ),
    .C(\alu/_1179_ ),
    .Y(\wAluOut[7] ));
 sky130_fd_sc_hd__mux2_1 \alu/_2069_  (.A0(net194),
    .A1(net190),
    .S(net228),
    .X(\alu/_1180_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2070_  (.A0(\alu/_1180_ ),
    .A1(\alu/_1127_ ),
    .S(net210),
    .X(\alu/_1181_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2071_  (.A0(\alu/_1181_ ),
    .A1(\alu/_1032_ ),
    .S(net179),
    .X(\alu/_1182_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2072_  (.A0(\alu/_1182_ ),
    .A1(\alu/_0742_ ),
    .S(net197),
    .X(\alu/_1183_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2073_  (.A(\alu/_1183_ ),
    .B(\alu/_1018_ ),
    .Y(\alu/_1184_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2074_  (.A(net194),
    .B(\wAluB[8] ),
    .Y(\alu/_1185_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2075_  (.A(\alu/_0355_ ),
    .Y(\alu/_1186_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2076_  (.A1(net194),
    .A2(\wAluB[8] ),
    .B1(\alu/_1136_ ),
    .Y(\alu/_1187_ ));
 sky130_fd_sc_hd__o221a_1 \alu/_2077_  (.A1(\alu/_1185_ ),
    .A2(\alu/_1134_ ),
    .B1(\alu/_1186_ ),
    .B2(\alu/_1135_ ),
    .C1(\alu/_1187_ ),
    .X(\alu/_1188_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2078_  (.A(\alu/_0830_ ),
    .B(net197),
    .Y(\alu/_1189_ ));
 sky130_fd_sc_hd__o211ai_1 \alu/_2079_  (.A1(net197),
    .A2(\alu/_0728_ ),
    .B1(\alu/_0732_ ),
    .C1(\alu/_1189_ ),
    .Y(\alu/_1190_ ));
 sky130_fd_sc_hd__and3_1 \alu/_2080_  (.A(\alu/_1184_ ),
    .B(\alu/_1188_ ),
    .C(\alu/_1190_ ),
    .X(\alu/_1191_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2081_  (.A(\alu/_0764_ ),
    .B(\alu/_1186_ ),
    .Y(\alu/_1192_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_2082_  (.A(\alu/_0935_ ),
    .X(\alu/_1193_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2083_  (.A(\alu/_1192_ ),
    .B(\alu/_1193_ ),
    .Y(\alu/_1194_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2084_  (.A1(\alu/_0355_ ),
    .A2(\alu/_0759_ ),
    .A3(\alu/_0763_ ),
    .B1(\alu/_1194_ ),
    .X(\alu/_1195_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2085_  (.A(\alu/_0875_ ),
    .B(net192),
    .Y(\alu/_1196_ ));
 sky130_fd_sc_hd__a2bb2o_1 \alu/_2086_  (.A1_N(\alu/_0947_ ),
    .A2_N(\alu/_1196_ ),
    .B1(\alu/_0970_ ),
    .B2(\alu/_0815_ ),
    .X(\alu/_1197_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2087_  (.A(\alu/_0532_ ),
    .B(\alu/_0537_ ),
    .Y(\alu/_1198_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2088_  (.A(\alu/_0544_ ),
    .B(\alu/_0550_ ),
    .Y(\alu/_1199_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2089_  (.A(\alu/_1198_ ),
    .B(\alu/_1199_ ),
    .Y(\alu/_1200_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2090_  (.A(\alu/_1064_ ),
    .B(\alu/_1200_ ),
    .Y(\alu/_1201_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2091_  (.A(\alu/_1198_ ),
    .B(\alu/_1106_ ),
    .Y(\alu/_1202_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2092_  (.A1(\alu/_1133_ ),
    .A2(\alu/_1156_ ),
    .B1(\alu/_1154_ ),
    .Y(\alu/_1203_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2093_  (.A(\alu/_1202_ ),
    .B(\alu/_1203_ ),
    .Y(\alu/_1204_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2094_  (.A(\alu/_1201_ ),
    .B(\alu/_1204_ ),
    .Y(\alu/_1205_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2095_  (.A(\alu/_1205_ ),
    .B(\alu/_0355_ ),
    .Y(\alu/_1206_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2096_  (.A(\alu/_1206_ ),
    .B(\alu/_1060_ ),
    .Y(\alu/_1207_ ));
 sky130_fd_sc_hd__o21ba_1 \alu/_2097_  (.A1(\alu/_0355_ ),
    .A2(\alu/_1205_ ),
    .B1_N(\alu/_1207_ ),
    .X(\alu/_1208_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2098_  (.A1(\alu/_1197_ ),
    .A2(net169),
    .B1(\alu/_1208_ ),
    .Y(\alu/_1209_ ));
 sky130_fd_sc_hd__nand3_4 \alu/_2099_  (.A(\alu/_1191_ ),
    .B(\alu/_1195_ ),
    .C(\alu/_1209_ ),
    .Y(\wAluOut[8] ));
 sky130_fd_sc_hd__nor2_1 \alu/_2100_  (.A(\alu/_0720_ ),
    .B(\alu/_0864_ ),
    .Y(\alu/_1210_ ));
 sky130_fd_sc_hd__a211o_1 \alu/_2101_  (.A1(\alu/_0911_ ),
    .A2(\alu/_1047_ ),
    .B1(\alu/_0913_ ),
    .C1(\alu/_1210_ ),
    .X(\alu/_1211_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2102_  (.A(\alu/_0889_ ),
    .Y(\alu/_1212_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2103_  (.A0(\wAluA[9] ),
    .A1(\wAluA[8] ),
    .S(net228),
    .X(\alu/_1213_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2104_  (.A(net213),
    .B(\alu/_1213_ ),
    .X(\alu/_1214_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2105_  (.A1(\alu/_0857_ ),
    .A2(\alu/_1150_ ),
    .B1(\alu/_1214_ ),
    .Y(\alu/_1215_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2106_  (.A0(\alu/_1215_ ),
    .A1(\alu/_1087_ ),
    .S(net180),
    .X(\alu/_1216_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2107_  (.A(\alu/_1216_ ),
    .B(\alu/_0832_ ),
    .Y(\alu/_1217_ ));
 sky130_fd_sc_hd__o211ai_1 \alu/_2108_  (.A1(\alu/_0805_ ),
    .A2(\alu/_1212_ ),
    .B1(\alu/_0883_ ),
    .C1(\alu/_1217_ ),
    .Y(\alu/_1218_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2109_  (.A(\wAluA[9] ),
    .B(\wAluB[9] ),
    .Y(\alu/_1219_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2110_  (.A(\alu/_0313_ ),
    .Y(\alu/_1220_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2111_  (.A(\wAluA[9] ),
    .B(\wAluB[9] ),
    .Y(\alu/_1221_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2112_  (.A(\alu/_1221_ ),
    .B(\alu/_0740_ ),
    .X(\alu/_1222_ ));
 sky130_fd_sc_hd__o221a_1 \alu/_2113_  (.A1(\alu/_1219_ ),
    .A2(\alu/_0838_ ),
    .B1(\alu/_1220_ ),
    .B2(\alu/_1135_ ),
    .C1(\alu/_1222_ ),
    .X(\alu/_1223_ ));
 sky130_fd_sc_hd__and3_1 \alu/_2114_  (.A(\alu/_1211_ ),
    .B(\alu/_1218_ ),
    .C(\alu/_1223_ ),
    .X(\alu/_1224_ ));
 sky130_fd_sc_hd__nor2_2 \alu/_2115_  (.A(\alu/_0971_ ),
    .B(\alu/_0835_ ),
    .Y(\alu/_1225_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_2116_  (.A(\alu/_0831_ ),
    .X(\alu/_1226_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2117_  (.A1(\alu/_0873_ ),
    .A2(\alu/_1226_ ),
    .B1(\alu/_1166_ ),
    .Y(\alu/_1227_ ));
 sky130_fd_sc_hd__o2bb2ai_2 \alu/_2118_  (.A1_N(\alu/_0853_ ),
    .A2_N(\alu/_1225_ ),
    .B1(\alu/_0877_ ),
    .B2(\alu/_1227_ ),
    .Y(\alu/_1228_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2119_  (.A(\alu/_1228_ ),
    .B(net170),
    .Y(\alu/_1229_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2120_  (.A1(\alu/_1206_ ),
    .A2(\alu/_1185_ ),
    .B1(\alu/_1220_ ),
    .Y(\alu/_1230_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2121_  (.A1(\alu/_1206_ ),
    .A2(\alu/_1185_ ),
    .A3(\alu/_1220_ ),
    .B1(\alu/_1074_ ),
    .X(\alu/_1231_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2122_  (.A(\alu/_1192_ ),
    .B(\alu/_0344_ ),
    .Y(\alu/_1232_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2123_  (.A1(\alu/_1220_ ),
    .A2(\alu/_1232_ ),
    .B1(\alu/_0935_ ),
    .Y(\alu/_1233_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2124_  (.A1(\alu/_1220_ ),
    .A2(\alu/_1232_ ),
    .B1(\alu/_1233_ ),
    .X(\alu/_1234_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_2125_  (.A1(\alu/_1230_ ),
    .A2(\alu/_1231_ ),
    .B1(\alu/_1234_ ),
    .X(\alu/_1235_ ));
 sky130_fd_sc_hd__nand3_4 \alu/_2126_  (.A(\alu/_1224_ ),
    .B(\alu/_1229_ ),
    .C(\alu/_1235_ ),
    .Y(\wAluOut[9] ));
 sky130_fd_sc_hd__nor2_1 \alu/_2127_  (.A(net195),
    .B(\alu/_0967_ ),
    .Y(\alu/_1236_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2128_  (.A1(\alu/_0805_ ),
    .A2(\alu/_0945_ ),
    .B1(\alu/_0733_ ),
    .Y(\alu/_1237_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2129_  (.A0(\alu/_0429_ ),
    .A1(\alu/_0291_ ),
    .S(net222),
    .X(\alu/_1238_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2130_  (.A(\alu/_1238_ ),
    .B(\alu/_0716_ ),
    .Y(\alu/_1239_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2131_  (.A1(\alu/_0822_ ),
    .A2(\alu/_1180_ ),
    .B1(\alu/_1239_ ),
    .Y(\alu/_1240_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2132_  (.A0(\alu/_1129_ ),
    .A1(\alu/_1240_ ),
    .S(\alu/_0817_ ),
    .X(\alu/_1241_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2133_  (.A(\alu/_1241_ ),
    .B(\alu/_0805_ ),
    .Y(\alu/_1242_ ));
 sky130_fd_sc_hd__o211ai_2 \alu/_2134_  (.A1(\alu/_0721_ ),
    .A2(\alu/_0981_ ),
    .B1(\alu/_1018_ ),
    .C1(\alu/_1242_ ),
    .Y(\alu/_1243_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2135_  (.A(\wAluA[10] ),
    .B(\wAluB[10] ),
    .Y(\alu/_1244_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2136_  (.A(\alu/_0472_ ),
    .Y(\alu/_1245_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2137_  (.A1(\wAluA[10] ),
    .A2(\wAluB[10] ),
    .B1(\alu/_0933_ ),
    .Y(\alu/_1246_ ));
 sky130_fd_sc_hd__o221a_1 \alu/_2138_  (.A1(\alu/_1244_ ),
    .A2(\alu/_1134_ ),
    .B1(\alu/_1245_ ),
    .B2(\alu/_0893_ ),
    .C1(\alu/_1246_ ),
    .X(\alu/_1247_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2139_  (.A1(\alu/_1236_ ),
    .A2(\alu/_1237_ ),
    .B1(\alu/_1243_ ),
    .C1(\alu/_1247_ ),
    .X(\alu/_1248_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2140_  (.A1(\alu/_0953_ ),
    .A2(\alu/_1226_ ),
    .B1(\alu/_1166_ ),
    .Y(\alu/_1249_ ));
 sky130_fd_sc_hd__o2bb2ai_4 \alu/_2141_  (.A1_N(\alu/_0958_ ),
    .A2_N(\alu/_1225_ ),
    .B1(\alu/_0877_ ),
    .B2(\alu/_1249_ ),
    .Y(\alu/_1250_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2142_  (.A(\alu/_1250_ ),
    .B(net169),
    .Y(\alu/_1251_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2143_  (.A1(\alu/_0764_ ),
    .A2(\alu/_0366_ ),
    .B1(\alu/_0766_ ),
    .X(\alu/_1252_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2144_  (.A(\alu/_1252_ ),
    .B(\alu/_1245_ ),
    .Y(\alu/_1253_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2145_  (.A(\alu/_1245_ ),
    .B(\alu/_1252_ ),
    .X(\alu/_1254_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2146_  (.A1(\alu/_1185_ ),
    .A2(\alu/_1221_ ),
    .B1(\alu/_1219_ ),
    .Y(\alu/_1255_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2147_  (.A(\alu/_1255_ ),
    .Y(\alu/_1256_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2148_  (.A(\alu/_1220_ ),
    .B(\alu/_1186_ ),
    .Y(\alu/_1257_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2149_  (.A(\alu/_1205_ ),
    .B(\alu/_1257_ ),
    .Y(\alu/_1258_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2150_  (.A1(\alu/_1258_ ),
    .A2(\alu/_1256_ ),
    .B1(\alu/_1245_ ),
    .X(\alu/_1259_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2151_  (.A(\alu/_1259_ ),
    .B(\alu/_1060_ ),
    .Y(\alu/_1260_ ));
 sky130_fd_sc_hd__a31oi_1 \alu/_2152_  (.A1(\alu/_1245_ ),
    .A2(\alu/_1256_ ),
    .A3(\alu/_1258_ ),
    .B1(\alu/_1260_ ),
    .Y(\alu/_1261_ ));
 sky130_fd_sc_hd__a31oi_2 \alu/_2153_  (.A1(\alu/_1055_ ),
    .A2(\alu/_1253_ ),
    .A3(\alu/_1254_ ),
    .B1(\alu/_1261_ ),
    .Y(\alu/_1262_ ));
 sky130_fd_sc_hd__nand3_4 \alu/_2154_  (.A(\alu/_1248_ ),
    .B(\alu/_1251_ ),
    .C(\alu/_1262_ ),
    .Y(\wAluOut[10] ));
 sky130_fd_sc_hd__nand2_1 \alu/_2155_  (.A(\alu/_0397_ ),
    .B(\alu/_0376_ ),
    .Y(\alu/_1263_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2156_  (.A(net237),
    .B(\wAluB[11] ),
    .Y(\alu/_1264_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_2157_  (.A(\alu/_1263_ ),
    .B(\alu/_1264_ ),
    .Y(\alu/_1265_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2158_  (.A1(\alu/_1259_ ),
    .A2(\alu/_1244_ ),
    .B1(\alu/_1265_ ),
    .Y(\alu/_1266_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2159_  (.A1(\alu/_1259_ ),
    .A2(\alu/_1265_ ),
    .A3(\alu/_1244_ ),
    .B1(\alu/_1074_ ),
    .X(\alu/_1267_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2160_  (.A(\alu/_1253_ ),
    .B(\alu/_0461_ ),
    .Y(\alu/_1268_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2161_  (.A1(\alu/_1265_ ),
    .A2(\alu/_1268_ ),
    .B1(\alu/_1193_ ),
    .Y(\alu/_1269_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2162_  (.A1(\alu/_1265_ ),
    .A2(\alu/_1268_ ),
    .B1(\alu/_1269_ ),
    .X(\alu/_1270_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2163_  (.A1(\alu/_1013_ ),
    .A2(\alu/_0831_ ),
    .B1(\alu/_1166_ ),
    .X(\alu/_1271_ ));
 sky130_fd_sc_hd__a22o_1 \alu/_2164_  (.A1(\alu/_1009_ ),
    .A2(\alu/_1225_ ),
    .B1(\alu/_1271_ ),
    .B2(\alu/_0956_ ),
    .X(\alu/_1272_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2165_  (.A1(\alu/_0947_ ),
    .A2(\alu/_1004_ ),
    .B1(\alu/_0732_ ),
    .Y(\alu/_1273_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2166_  (.A1(\alu/_1226_ ),
    .A2(\alu/_0992_ ),
    .B1(\alu/_1273_ ),
    .X(\alu/_1274_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2167_  (.A0(\wAluA[11] ),
    .A1(\wAluA[10] ),
    .S(net223),
    .X(\alu/_1275_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2168_  (.A0(\alu/_1275_ ),
    .A1(\alu/_1213_ ),
    .S(net212),
    .X(\alu/_1276_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2169_  (.A0(\alu/_1276_ ),
    .A1(\alu/_1151_ ),
    .S(net181),
    .X(\alu/_1277_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2170_  (.A(\alu/_1277_ ),
    .B(\alu/_0986_ ),
    .Y(\alu/_1278_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2171_  (.A1(\alu/_0986_ ),
    .A2(\alu/_1021_ ),
    .B1(\alu/_1278_ ),
    .Y(\alu/_1279_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2172_  (.A(\alu/_1279_ ),
    .B(\alu/_1018_ ),
    .Y(\alu/_1280_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_2173_  (.A(\alu/_0892_ ),
    .X(\alu/_1281_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2174_  (.A(\alu/_0933_ ),
    .B(\alu/_1263_ ),
    .Y(\alu/_1282_ ));
 sky130_fd_sc_hd__o221a_1 \alu/_2175_  (.A1(\alu/_1264_ ),
    .A2(\alu/_1134_ ),
    .B1(\alu/_1265_ ),
    .B2(\alu/_1281_ ),
    .C1(\alu/_1282_ ),
    .X(\alu/_1283_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2176_  (.A(\alu/_1274_ ),
    .B(\alu/_1280_ ),
    .C(\alu/_1283_ ),
    .Y(\alu/_1284_ ));
 sky130_fd_sc_hd__a21oi_2 \alu/_2177_  (.A1(\alu/_1272_ ),
    .A2(net172),
    .B1(\alu/_1284_ ),
    .Y(\alu/_1285_ ));
 sky130_fd_sc_hd__o211ai_4 \alu/_2178_  (.A1(\alu/_1266_ ),
    .A2(\alu/_1267_ ),
    .B1(\alu/_1270_ ),
    .C1(\alu/_1285_ ),
    .Y(\wAluOut[11] ));
 sky130_fd_sc_hd__a31o_1 \alu/_2179_  (.A1(\alu/_0764_ ),
    .A2(\alu/_0366_ ),
    .A3(\alu/_0482_ ),
    .B1(\alu/_0769_ ),
    .X(\alu/_1286_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2180_  (.A(\alu/_1286_ ),
    .B(\alu/_0511_ ),
    .Y(\alu/_1287_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2181_  (.A(\alu/_0511_ ),
    .B(\alu/_1286_ ),
    .X(\alu/_1288_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2182_  (.A(\alu/_1265_ ),
    .B(\alu/_1245_ ),
    .Y(\alu/_1289_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2183_  (.A(\alu/_1289_ ),
    .B(\alu/_1255_ ),
    .Y(\alu/_1290_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2184_  (.A(net237),
    .B(\wAluB[11] ),
    .Y(\alu/_1291_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_2185_  (.A1(\alu/_1244_ ),
    .A2(\alu/_1291_ ),
    .B1(\alu/_1264_ ),
    .X(\alu/_1292_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2186_  (.A(\alu/_1290_ ),
    .B(\alu/_1292_ ),
    .Y(\alu/_1293_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2187_  (.A1(\alu/_1205_ ),
    .A2(\alu/_1257_ ),
    .A3(\alu/_1289_ ),
    .B1(\alu/_1293_ ),
    .X(\alu/_1294_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2188_  (.A(\alu/_0512_ ),
    .B(\alu/_1294_ ),
    .X(\alu/_1295_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2189_  (.A(\alu/_1294_ ),
    .B(\alu/_0512_ ),
    .Y(\alu/_1296_ ));
 sky130_fd_sc_hd__and3_1 \alu/_2190_  (.A(\alu/_1295_ ),
    .B(\alu/_1060_ ),
    .C(\alu/_1296_ ),
    .X(\alu/_1297_ ));
 sky130_fd_sc_hd__a31oi_1 \alu/_2191_  (.A1(\alu/_1055_ ),
    .A2(\alu/_1287_ ),
    .A3(\alu/_1288_ ),
    .B1(\alu/_1297_ ),
    .Y(\alu/_1298_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2192_  (.A0(\wAluA[12] ),
    .A1(net237),
    .S(net223),
    .X(\alu/_1299_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2193_  (.A(\alu/_1299_ ),
    .B(\alu/_0822_ ),
    .Y(\alu/_1300_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2194_  (.A1(\alu/_0822_ ),
    .A2(\alu/_1238_ ),
    .B1(\alu/_1300_ ),
    .Y(\alu/_1301_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2195_  (.A0(\alu/_1181_ ),
    .A1(\alu/_1301_ ),
    .S(\alu/_0816_ ),
    .X(\alu/_1302_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2196_  (.A0(\alu/_1302_ ),
    .A1(\alu/_1033_ ),
    .S(net198),
    .X(\alu/_1303_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2197_  (.A(\alu/_1303_ ),
    .B(\alu/_1018_ ),
    .Y(\alu/_1304_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2198_  (.A(net195),
    .B(\alu/_1039_ ),
    .X(\alu/_1305_ ));
 sky130_fd_sc_hd__o211ai_1 \alu/_2199_  (.A1(\alu/_0832_ ),
    .A2(\alu/_1046_ ),
    .B1(\alu/_0732_ ),
    .C1(\alu/_1305_ ),
    .Y(\alu/_1306_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2200_  (.A(\alu/_1225_ ),
    .Y(\alu/_1307_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2201_  (.A1(\alu/_1050_ ),
    .A2(\alu/_0709_ ),
    .B1(\alu/_1166_ ),
    .X(\alu/_1308_ ));
 sky130_fd_sc_hd__a2bb2o_1 \alu/_2202_  (.A1_N(\alu/_1045_ ),
    .A2_N(\alu/_1307_ ),
    .B1(\alu/_0956_ ),
    .B2(\alu/_1308_ ),
    .X(\alu/_1309_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2203_  (.A(\alu/_1309_ ),
    .B(net172),
    .Y(\alu/_1310_ ));
 sky130_fd_sc_hd__and3_1 \alu/_2204_  (.A(\alu/_1304_ ),
    .B(\alu/_1306_ ),
    .C(\alu/_1310_ ),
    .X(\alu/_1311_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2205_  (.A(\alu/_0933_ ),
    .B(\alu/_0509_ ),
    .Y(\alu/_1312_ ));
 sky130_fd_sc_hd__o221a_1 \alu/_2206_  (.A1(\alu/_0510_ ),
    .A2(\alu/_0741_ ),
    .B1(\alu/_0511_ ),
    .B2(\alu/_0929_ ),
    .C1(\alu/_1312_ ),
    .X(\alu/_1313_ ));
 sky130_fd_sc_hd__nand3_2 \alu/_2207_  (.A(\alu/_1298_ ),
    .B(\alu/_1311_ ),
    .C(\alu/_1313_ ),
    .Y(\wAluOut[12] ));
 sky130_fd_sc_hd__a21o_1 \alu/_2208_  (.A1(\alu/_1098_ ),
    .A2(\alu/_0709_ ),
    .B1(\alu/_1165_ ),
    .X(\alu/_1314_ ));
 sky130_fd_sc_hd__a2bb2o_2 \alu/_2209_  (.A1_N(\alu/_1307_ ),
    .A2_N(\alu/_1101_ ),
    .B1(\alu/_0956_ ),
    .B2(\alu/_1314_ ),
    .X(\alu/_1315_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2210_  (.A(\wAluA[13] ),
    .B(\wAluB[13] ),
    .Y(\alu/_1316_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2211_  (.A(\alu/_1316_ ),
    .Y(\alu/_1317_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2212_  (.A(\alu/_0502_ ),
    .B(\alu/_0504_ ),
    .Y(\alu/_1318_ ));
 sky130_fd_sc_hd__a22o_1 \alu/_2213_  (.A1(\alu/_0930_ ),
    .A2(\alu/_1317_ ),
    .B1(\alu/_1318_ ),
    .B2(\alu/_1136_ ),
    .X(\alu/_1319_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2214_  (.A(\alu/_1318_ ),
    .B(\alu/_1316_ ),
    .Y(\alu/_1320_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2215_  (.A(\alu/_1320_ ),
    .B(\alu/_0929_ ),
    .Y(\alu/_1321_ ));
 sky130_fd_sc_hd__a211o_1 \alu/_2216_  (.A1(\alu/_1315_ ),
    .A2(net169),
    .B1(\alu/_1319_ ),
    .C1(\alu/_1321_ ),
    .X(\alu/_1322_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2217_  (.A(\alu/_0947_ ),
    .B(\alu/_1095_ ),
    .Y(\alu/_1323_ ));
 sky130_fd_sc_hd__a211o_1 \alu/_2218_  (.A1(\alu/_0832_ ),
    .A2(\alu/_1079_ ),
    .B1(\alu/_0913_ ),
    .C1(\alu/_1323_ ),
    .X(\alu/_1324_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2219_  (.A0(\alu/_0502_ ),
    .A1(\alu/_0507_ ),
    .S(net222),
    .X(\alu/_1325_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2220_  (.A(\alu/_1325_ ),
    .B(\alu/_0845_ ),
    .Y(\alu/_1326_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2221_  (.A1(\alu/_0845_ ),
    .A2(\alu/_1275_ ),
    .B1(\alu/_1326_ ),
    .Y(\alu/_1327_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2222_  (.A(net180),
    .B(\alu/_1327_ ),
    .X(\alu/_1328_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_2223_  (.A1(\alu/_0888_ ),
    .A2(\alu/_1215_ ),
    .B1(\alu/_1328_ ),
    .X(\alu/_1329_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2224_  (.A(\alu/_1089_ ),
    .B(net199),
    .Y(\alu/_1330_ ));
 sky130_fd_sc_hd__o21ai_2 \alu/_2225_  (.A1(net199),
    .A2(\alu/_1329_ ),
    .B1(\alu/_1330_ ),
    .Y(\alu/_1331_ ));
 sky130_fd_sc_hd__buf_2 \alu/_2226_  (.A(\alu/_0746_ ),
    .X(\alu/_1332_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2227_  (.A(\alu/_1331_ ),
    .B(\alu/_1332_ ),
    .Y(\alu/_1333_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2228_  (.A(\alu/_1324_ ),
    .B(\alu/_1333_ ),
    .Y(\alu/_1334_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2229_  (.A(\alu/_1322_ ),
    .B(\alu/_1334_ ),
    .Y(\alu/_1335_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2230_  (.A(\alu/_1287_ ),
    .B(\alu/_0771_ ),
    .Y(\alu/_1336_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2231_  (.A1(\alu/_1320_ ),
    .A2(\alu/_1336_ ),
    .B1(\alu/_1114_ ),
    .Y(\alu/_1337_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2232_  (.A1(\alu/_1320_ ),
    .A2(\alu/_1336_ ),
    .B1(\alu/_1337_ ),
    .X(\alu/_1338_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2233_  (.A(\alu/_1296_ ),
    .B(\alu/_0510_ ),
    .Y(\alu/_1339_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2234_  (.A1(\alu/_0506_ ),
    .A2(\alu/_1339_ ),
    .B1(\alu/_1177_ ),
    .Y(\alu/_1340_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2235_  (.A1(\alu/_0506_ ),
    .A2(\alu/_1339_ ),
    .B1(\alu/_1340_ ),
    .X(\alu/_0000_ ));
 sky130_fd_sc_hd__nand3_2 \alu/_2236_  (.A(\alu/_1335_ ),
    .B(\alu/_1338_ ),
    .C(\alu/_0000_ ),
    .Y(\wAluOut[13] ));
 sky130_fd_sc_hd__nand2_1 \alu/_2237_  (.A(\alu/_1142_ ),
    .B(\alu/_1226_ ),
    .Y(\alu/_0001_ ));
 sky130_fd_sc_hd__o211ai_1 \alu/_2238_  (.A1(\alu/_1226_ ),
    .A2(\alu/_1117_ ),
    .B1(\alu/_0732_ ),
    .C1(\alu/_0001_ ),
    .Y(\alu/_0002_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2239_  (.A(\alu/_1299_ ),
    .B(net212),
    .Y(\alu/_0003_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2240_  (.A0(\wAluA[14] ),
    .A1(\wAluA[13] ),
    .S(net223),
    .X(\alu/_0004_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2241_  (.A(\alu/_0004_ ),
    .B(\alu/_0716_ ),
    .Y(\alu/_0005_ ));
 sky130_fd_sc_hd__and2_1 \alu/_2242_  (.A(\alu/_0003_ ),
    .B(\alu/_0005_ ),
    .X(\alu/_0006_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2243_  (.A(\alu/_0704_ ),
    .B(\alu/_1240_ ),
    .X(\alu/_0007_ ));
 sky130_fd_sc_hd__o21ai_2 \alu/_2244_  (.A1(net180),
    .A2(\alu/_0006_ ),
    .B1(\alu/_0007_ ),
    .Y(\alu/_0008_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2245_  (.A(\alu/_0946_ ),
    .B(\alu/_1131_ ),
    .X(\alu/_0009_ ));
 sky130_fd_sc_hd__o211ai_1 \alu/_2246_  (.A1(net203),
    .A2(\alu/_0008_ ),
    .B1(\alu/_0883_ ),
    .C1(\alu/_0009_ ),
    .Y(\alu/_0010_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2247_  (.A1(\alu/_1120_ ),
    .A2(\alu/_0709_ ),
    .B1(\alu/_1166_ ),
    .X(\alu/_0011_ ));
 sky130_fd_sc_hd__a2bb2o_1 \alu/_2248_  (.A1_N(\alu/_1119_ ),
    .A2_N(\alu/_1307_ ),
    .B1(\alu/_0956_ ),
    .B2(\alu/_0011_ ),
    .X(\alu/_0012_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2249_  (.A(\alu/_0012_ ),
    .B(net171),
    .Y(\alu/_0013_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2250_  (.A(\wAluA[14] ),
    .B(\wAluB[14] ),
    .Y(\alu/_0014_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2251_  (.A(\alu/_0524_ ),
    .Y(\alu/_0015_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2252_  (.A1(\wAluA[14] ),
    .A2(\wAluB[14] ),
    .B1(\alu/_1136_ ),
    .Y(\alu/_0016_ ));
 sky130_fd_sc_hd__o221a_1 \alu/_2253_  (.A1(\alu/_0014_ ),
    .A2(\alu/_1083_ ),
    .B1(\alu/_0015_ ),
    .B2(\alu/_0928_ ),
    .C1(\alu/_0016_ ),
    .X(\alu/_0017_ ));
 sky130_fd_sc_hd__and4_2 \alu/_2254_  (.A(\alu/_0002_ ),
    .B(\alu/_0010_ ),
    .C(\alu/_0013_ ),
    .D(\alu/_0017_ ),
    .X(\alu/_0018_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2255_  (.A1(\alu/_1286_ ),
    .A2(\alu/_0513_ ),
    .B1(\alu/_0772_ ),
    .X(\alu/_0019_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2256_  (.A(\alu/_0015_ ),
    .B(\alu/_0019_ ),
    .X(\alu/_0020_ ));
 sky130_fd_sc_hd__buf_2 \alu/_2257_  (.A(\alu/_1193_ ),
    .X(\alu/_0021_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2258_  (.A(\alu/_0019_ ),
    .B(\alu/_0015_ ),
    .Y(\alu/_0022_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2259_  (.A(\alu/_0020_ ),
    .B(\alu/_0021_ ),
    .C(\alu/_0022_ ),
    .Y(\alu/_0023_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2260_  (.A(\alu/_1320_ ),
    .B(\alu/_0511_ ),
    .Y(\alu/_0024_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2261_  (.A1(\alu/_0510_ ),
    .A2(\alu/_1320_ ),
    .B1(\alu/_1316_ ),
    .Y(\alu/_0025_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2262_  (.A1(\alu/_1294_ ),
    .A2(\alu/_0024_ ),
    .B1(\alu/_0025_ ),
    .X(\alu/_0026_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2263_  (.A(\alu/_0524_ ),
    .B(\alu/_0026_ ),
    .X(\alu/_0027_ ));
 sky130_fd_sc_hd__buf_2 \alu/_2264_  (.A(\alu/_1177_ ),
    .X(\alu/_0028_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2265_  (.A(\alu/_0026_ ),
    .B(\alu/_0524_ ),
    .Y(\alu/_0029_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2266_  (.A(\alu/_0027_ ),
    .B(\alu/_0028_ ),
    .C(\alu/_0029_ ),
    .Y(\alu/_0030_ ));
 sky130_fd_sc_hd__nand3_2 \alu/_2267_  (.A(\alu/_0018_ ),
    .B(\alu/_0023_ ),
    .C(\alu/_0030_ ),
    .Y(\wAluOut[14] ));
 sky130_fd_sc_hd__inv_2 \alu/_2268_  (.A(\alu/_0519_ ),
    .Y(\alu/_0031_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2269_  (.A1(\alu/_0029_ ),
    .A2(\alu/_0014_ ),
    .B1(\alu/_0031_ ),
    .X(\alu/_0032_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2270_  (.A(\alu/_0029_ ),
    .B(\alu/_0031_ ),
    .C(\alu/_0014_ ),
    .Y(\alu/_0033_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2271_  (.A(\alu/_0032_ ),
    .B(\alu/_0028_ ),
    .C(\alu/_0033_ ),
    .Y(\alu/_0034_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2272_  (.A(\alu/_0022_ ),
    .B(\alu/_0523_ ),
    .Y(\alu/_0035_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2273_  (.A(\alu/_0035_ ),
    .B(\alu/_0031_ ),
    .Y(\alu/_0036_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2274_  (.A(\alu/_0022_ ),
    .B(\alu/_0519_ ),
    .C(\alu/_0523_ ),
    .Y(\alu/_0037_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2275_  (.A(\alu/_0036_ ),
    .B(\alu/_0021_ ),
    .C(\alu/_0037_ ),
    .Y(\alu/_0038_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2276_  (.A0(\alu/_0516_ ),
    .A1(\alu/_0520_ ),
    .S(net225),
    .X(\alu/_0039_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2277_  (.A(\alu/_0039_ ),
    .B(\alu/_0715_ ),
    .Y(\alu/_0040_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2278_  (.A(\alu/_1325_ ),
    .B(net212),
    .Y(\alu/_0041_ ));
 sky130_fd_sc_hd__and2_1 \alu/_2279_  (.A(\alu/_0040_ ),
    .B(\alu/_0041_ ),
    .X(\alu/_0042_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2280_  (.A0(\alu/_1276_ ),
    .A1(\alu/_0042_ ),
    .S(\alu/_0217_ ),
    .X(\alu/_0043_ ));
 sky130_fd_sc_hd__mux2_2 \alu/_2281_  (.A0(\alu/_0043_ ),
    .A1(\alu/_1152_ ),
    .S(net198),
    .X(\alu/_0044_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2282_  (.A(\wAluA[15] ),
    .B(\wAluB[15] ),
    .Y(\alu/_0045_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2283_  (.A(\alu/_1168_ ),
    .B(\alu/_0709_ ),
    .Y(\alu/_0046_ ));
 sky130_fd_sc_hd__or3_1 \alu/_2284_  (.A(\alu/_0804_ ),
    .B(\alu/_0046_ ),
    .C(\alu/_0835_ ),
    .X(\alu/_0047_ ));
 sky130_fd_sc_hd__or2_2 \alu/_2285_  (.A(\alu/_0548_ ),
    .B(\alu/_1196_ ),
    .X(\alu/_0048_ ));
 sky130_fd_sc_hd__buf_6 \alu/_2286_  (.A(\alu/_0048_ ),
    .X(\alu/_0049_ ));
 sky130_fd_sc_hd__o211ai_1 \alu/_2287_  (.A1(\alu/_0045_ ),
    .A2(\alu/_0741_ ),
    .B1(\alu/_0047_ ),
    .C1(\alu/_0049_ ),
    .Y(\alu/_0050_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2288_  (.A(\alu/_1148_ ),
    .B(\alu/_0805_ ),
    .Y(\alu/_0051_ ));
 sky130_fd_sc_hd__o211ai_2 \alu/_2289_  (.A1(\alu/_0805_ ),
    .A2(\alu/_1163_ ),
    .B1(\alu/_0733_ ),
    .C1(\alu/_0051_ ),
    .Y(\alu/_0052_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2290_  (.A(\wAluA[15] ),
    .B(\wAluB[15] ),
    .Y(\alu/_0053_ ));
 sky130_fd_sc_hd__o22a_1 \alu/_2291_  (.A1(\alu/_0053_ ),
    .A2(\alu/_0838_ ),
    .B1(\alu/_0031_ ),
    .B2(\alu/_0929_ ),
    .X(\alu/_0054_ ));
 sky130_fd_sc_hd__nand3b_1 \alu/_2292_  (.A_N(\alu/_0050_ ),
    .B(\alu/_0052_ ),
    .C(\alu/_0054_ ),
    .Y(\alu/_0055_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2293_  (.A1(\alu/_1332_ ),
    .A2(\alu/_0044_ ),
    .B1(\alu/_0055_ ),
    .Y(\alu/_0056_ ));
 sky130_fd_sc_hd__nand3_2 \alu/_2294_  (.A(\alu/_0034_ ),
    .B(\alu/_0038_ ),
    .C(\alu/_0056_ ),
    .Y(\wAluOut[15] ));
 sky130_fd_sc_hd__mux2_2 \alu/_2295_  (.A0(\wAluA[16] ),
    .A1(\wAluA[15] ),
    .S(net224),
    .X(\alu/_0058_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2296_  (.A0(\alu/_0058_ ),
    .A1(\alu/_0004_ ),
    .S(net212),
    .X(\alu/_0059_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2297_  (.A0(\alu/_0059_ ),
    .A1(\alu/_1301_ ),
    .S(net181),
    .X(\alu/_0060_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2298_  (.A(\alu/_0711_ ),
    .B(\alu/_1182_ ),
    .X(\alu/_0061_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2299_  (.A1(net198),
    .A2(\alu/_0060_ ),
    .B1(\alu/_1332_ ),
    .C1(\alu/_0061_ ),
    .X(\alu/_0062_ ));
 sky130_fd_sc_hd__a2111o_1 \alu/_2300_  (.A1(\alu/_0648_ ),
    .A2(\alu/_0613_ ),
    .B1(\alu/_0729_ ),
    .C1(\alu/_0611_ ),
    .D1(\alu/_0651_ ),
    .X(\alu/_0063_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_2301_  (.A(\alu/_0048_ ),
    .X(\alu/_0064_ ));
 sky130_fd_sc_hd__or3_1 \alu/_2302_  (.A(\alu/_0548_ ),
    .B(\alu/_0743_ ),
    .C(\alu/_0745_ ),
    .X(\alu/_0065_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2303_  (.A1(\alu/_0612_ ),
    .A2(\alu/_0741_ ),
    .B1(\alu/_0064_ ),
    .C1(\alu/_0065_ ),
    .X(\alu/_0066_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2304_  (.A1(\alu/_0913_ ),
    .A2(\alu/_0834_ ),
    .B1(\alu/_0063_ ),
    .C1(\alu/_0066_ ),
    .X(\alu/_0067_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2305_  (.A(\alu/_0614_ ),
    .Y(\alu/_0069_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2306_  (.A(\alu/_0069_ ),
    .B(\alu/_0777_ ),
    .X(\alu/_0070_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2307_  (.A(\alu/_0777_ ),
    .B(\alu/_0069_ ),
    .Y(\alu/_0071_ ));
 sky130_fd_sc_hd__and3_1 \alu/_2308_  (.A(\alu/_0070_ ),
    .B(\alu/_0935_ ),
    .C(\alu/_0071_ ),
    .X(\alu/_0072_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2309_  (.A(\alu/_1257_ ),
    .B(\alu/_1289_ ),
    .Y(\alu/_0073_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2310_  (.A(\alu/_0518_ ),
    .B(\alu/_0524_ ),
    .Y(\alu/_0074_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2311_  (.A(\alu/_0074_ ),
    .Y(\alu/_0075_ ));
 sky130_fd_sc_hd__and2_1 \alu/_2312_  (.A(\alu/_0075_ ),
    .B(\alu/_0024_ ),
    .X(\alu/_0076_ ));
 sky130_fd_sc_hd__nor2b_1 \alu/_2313_  (.A(\alu/_0073_ ),
    .B_N(\alu/_0076_ ),
    .Y(\alu/_0077_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2314_  (.A(\alu/_1205_ ),
    .B(\alu/_0077_ ),
    .Y(\alu/_0078_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2315_  (.A(\alu/_0025_ ),
    .B(\alu/_0075_ ),
    .Y(\alu/_0080_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_2316_  (.A1(\alu/_0014_ ),
    .A2(\alu/_0053_ ),
    .B1(\alu/_0045_ ),
    .X(\alu/_0081_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2317_  (.A(\alu/_0080_ ),
    .B(\alu/_0081_ ),
    .Y(\alu/_0082_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2318_  (.A1(\alu/_1293_ ),
    .A2(\alu/_0076_ ),
    .B1(\alu/_0082_ ),
    .Y(\alu/_0083_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_2319_  (.A(\alu/_0078_ ),
    .B(\alu/_0083_ ),
    .Y(\alu/_0084_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2320_  (.A(\alu/_0614_ ),
    .B(\alu/_0084_ ),
    .X(\alu/_0085_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2321_  (.A(\alu/_0084_ ),
    .B(\alu/_0614_ ),
    .Y(\alu/_0086_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2322_  (.A(\alu/_0085_ ),
    .B(\alu/_1177_ ),
    .C(\alu/_0086_ ),
    .Y(\alu/_0087_ ));
 sky130_fd_sc_hd__and2b_1 \alu/_2323_  (.A_N(\alu/_0072_ ),
    .B(\alu/_0087_ ),
    .X(\alu/_0088_ ));
 sky130_fd_sc_hd__nand3b_4 \alu/_2324_  (.A_N(\alu/_0062_ ),
    .B(\alu/_0067_ ),
    .C(\alu/_0088_ ),
    .Y(\wAluOut[16] ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2325_  (.A1(\alu/_0869_ ),
    .A2(\alu/_0878_ ),
    .B1(net172),
    .Y(\alu/_0090_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2326_  (.A(\alu/_1216_ ),
    .B(net198),
    .Y(\alu/_0091_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2327_  (.A0(\alu/_0615_ ),
    .A1(\alu/_0656_ ),
    .S(net233),
    .X(\alu/_0092_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2328_  (.A0(\alu/_0092_ ),
    .A1(\alu/_0039_ ),
    .S(net220),
    .X(\alu/_0093_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2329_  (.A(\alu/_0816_ ),
    .B(\alu/_1327_ ),
    .X(\alu/_0094_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2330_  (.A1(net187),
    .A2(\alu/_0093_ ),
    .B1(\alu/_0094_ ),
    .Y(\alu/_0095_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2331_  (.A(net198),
    .B(\alu/_0095_ ),
    .X(\alu/_0096_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2332_  (.A(\alu/_0091_ ),
    .B(\alu/_0096_ ),
    .C(\alu/_0879_ ),
    .Y(\alu/_0097_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2333_  (.A(\alu/_0890_ ),
    .B(net171),
    .Y(\alu/_0098_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2334_  (.A1(\alu/_0097_ ),
    .A2(\alu/_0098_ ),
    .B1(\alu/_0976_ ),
    .X(\alu/_0099_ ));
 sky130_fd_sc_hd__o2bb2a_1 \alu/_2335_  (.A1_N(\alu/_0617_ ),
    .A2_N(\alu/_1136_ ),
    .B1(\alu/_0618_ ),
    .B2(\alu/_1083_ ),
    .X(\alu/_0101_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2336_  (.A1(\alu/_0655_ ),
    .A2(\alu/_0893_ ),
    .B1(\alu/_0064_ ),
    .C1(\alu/_0101_ ),
    .X(\alu/_0102_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2337_  (.A(\alu/_0099_ ),
    .B(\alu/_0102_ ),
    .Y(\alu/_0103_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2338_  (.A(\alu/_0090_ ),
    .B(\alu/_0103_ ),
    .Y(\alu/_0104_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2339_  (.A(\alu/_0071_ ),
    .B(\alu/_0780_ ),
    .Y(\alu/_0105_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2340_  (.A1(\alu/_0655_ ),
    .A2(\alu/_0105_ ),
    .B1(\alu/_1193_ ),
    .Y(\alu/_0106_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2341_  (.A1(\alu/_0655_ ),
    .A2(\alu/_0105_ ),
    .B1(\alu/_0106_ ),
    .X(\alu/_0107_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2342_  (.A1(\alu/_0086_ ),
    .A2(\alu/_0612_ ),
    .B1(\alu/_0655_ ),
    .X(\alu/_0108_ ));
 sky130_fd_sc_hd__buf_2 \alu/_2343_  (.A(\alu/_0899_ ),
    .X(\alu/_0109_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2344_  (.A(\alu/_0108_ ),
    .B(\alu/_0109_ ),
    .Y(\alu/_0110_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2345_  (.A1(\alu/_0612_ ),
    .A2(\alu/_0655_ ),
    .A3(\alu/_0086_ ),
    .B1(\alu/_0110_ ),
    .X(\alu/_0112_ ));
 sky130_fd_sc_hd__nand3_2 \alu/_2346_  (.A(\alu/_0104_ ),
    .B(\alu/_0107_ ),
    .C(\alu/_0112_ ),
    .Y(\wAluOut[17] ));
 sky130_fd_sc_hd__nor2_1 \alu/_2347_  (.A(\alu/_0619_ ),
    .B(\alu/_0069_ ),
    .Y(\alu/_0113_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2348_  (.A(\alu/_0084_ ),
    .B(\alu/_0113_ ),
    .Y(\alu/_0114_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_2349_  (.A1(\alu/_0612_ ),
    .A2(\alu/_0619_ ),
    .B1(\alu/_0618_ ),
    .X(\alu/_0115_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2350_  (.A(\alu/_0114_ ),
    .B(\alu/_0115_ ),
    .Y(\alu/_0116_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2351_  (.A(\alu/_0609_ ),
    .B(\alu/_0116_ ),
    .X(\alu/_0117_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2352_  (.A(\alu/_0116_ ),
    .B(\alu/_0609_ ),
    .Y(\alu/_0118_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2353_  (.A(\alu/_0117_ ),
    .B(\alu/_0118_ ),
    .Y(\alu/_0119_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2354_  (.A(\wAluA[18] ),
    .B(\wAluB[18] ),
    .Y(\alu/_0120_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2355_  (.A(\alu/_0120_ ),
    .B(\alu/_1083_ ),
    .X(\alu/_0122_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2356_  (.A(\wAluA[18] ),
    .B(\wAluB[18] ),
    .Y(\alu/_0123_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2357_  (.A(\alu/_0609_ ),
    .Y(\alu/_0124_ ));
 sky130_fd_sc_hd__o22a_1 \alu/_2358_  (.A1(\alu/_0123_ ),
    .A2(\alu/_0838_ ),
    .B1(\alu/_0124_ ),
    .B2(\alu/_1135_ ),
    .X(\alu/_0125_ ));
 sky130_fd_sc_hd__o2111a_1 \alu/_2359_  (.A1(\alu/_0879_ ),
    .A2(\alu/_0982_ ),
    .B1(\alu/_0122_ ),
    .C1(\alu/_0064_ ),
    .D1(\alu/_0125_ ),
    .X(\alu/_0126_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2360_  (.A(\alu/_0777_ ),
    .B(\alu/_0621_ ),
    .Y(\alu/_0127_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2361_  (.A(\alu/_0127_ ),
    .B(\alu/_0783_ ),
    .Y(\alu/_0128_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2362_  (.A(\alu/_0128_ ),
    .B(\alu/_0124_ ),
    .Y(\alu/_0129_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2363_  (.A(\alu/_0129_ ),
    .B(\alu/_0896_ ),
    .Y(\alu/_0130_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2364_  (.A1(\alu/_0609_ ),
    .A2(\alu/_0783_ ),
    .A3(\alu/_0127_ ),
    .B1(\alu/_0130_ ),
    .X(\alu/_0131_ ));
 sky130_fd_sc_hd__mux2_2 \alu/_2365_  (.A0(\wAluA[18] ),
    .A1(\wAluA[17] ),
    .S(net224),
    .X(\alu/_0133_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2366_  (.A(\alu/_0133_ ),
    .Y(\alu/_0134_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2367_  (.A(\alu/_0134_ ),
    .B(\alu/_0823_ ),
    .Y(\alu/_0135_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2368_  (.A1(\alu/_0823_ ),
    .A2(\alu/_0058_ ),
    .B1(\alu/_0135_ ),
    .Y(\alu/_0136_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2369_  (.A(\alu/_0851_ ),
    .B(\alu/_0006_ ),
    .X(\alu/_0137_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2370_  (.A1(net188),
    .A2(\alu/_0136_ ),
    .B1(\alu/_0137_ ),
    .Y(\alu/_0138_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2371_  (.A(\alu/_0745_ ),
    .Y(\alu/_0139_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2372_  (.A(\alu/_1241_ ),
    .B(net205),
    .Y(\alu/_0140_ ));
 sky130_fd_sc_hd__o211ai_1 \alu/_2373_  (.A1(net205),
    .A2(\alu/_0138_ ),
    .B1(\alu/_0139_ ),
    .C1(\alu/_0140_ ),
    .Y(\alu/_0141_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2374_  (.A(\alu/_0141_ ),
    .B(\alu/_0957_ ),
    .C(\alu/_0961_ ),
    .Y(\alu/_0142_ ));
 sky130_fd_sc_hd__buf_2 \alu/_2375_  (.A(\alu/_0880_ ),
    .X(\alu/_0144_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_2376_  (.A(\alu/_0142_ ),
    .B(\alu/_0144_ ),
    .Y(\alu/_0145_ ));
 sky130_fd_sc_hd__o2111ai_4 \alu/_2377_  (.A1(\alu/_1074_ ),
    .A2(\alu/_0119_ ),
    .B1(\alu/_0126_ ),
    .C1(\alu/_0131_ ),
    .D1(\alu/_0145_ ),
    .Y(\wAluOut[18] ));
 sky130_fd_sc_hd__mux2_1 \alu/_2378_  (.A0(\alu/_0600_ ),
    .A1(\alu/_0606_ ),
    .S(net229),
    .X(\alu/_0146_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2379_  (.A(\alu/_0845_ ),
    .B(\alu/_0092_ ),
    .X(\alu/_0147_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2380_  (.A1(net220),
    .A2(\alu/_0146_ ),
    .B1(\alu/_0147_ ),
    .Y(\alu/_0148_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2381_  (.A(\alu/_0851_ ),
    .B(\alu/_0042_ ),
    .X(\alu/_0149_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2382_  (.A1(net188),
    .A2(\alu/_0148_ ),
    .B1(\alu/_0149_ ),
    .Y(\alu/_0150_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2383_  (.A(\alu/_1277_ ),
    .B(net204),
    .Y(\alu/_0151_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2384_  (.A1(net204),
    .A2(\alu/_0150_ ),
    .B1(\alu/_0151_ ),
    .Y(\alu/_0152_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_2385_  (.A1(\alu/_0879_ ),
    .A2(\alu/_1022_ ),
    .B1(\alu/_0139_ ),
    .X(\alu/_0154_ ));
 sky130_fd_sc_hd__o21ai_2 \alu/_2386_  (.A1(net171),
    .A2(\alu/_0152_ ),
    .B1(\alu/_0154_ ),
    .Y(\alu/_0155_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_2387_  (.A(\alu/_0548_ ),
    .X(\alu/_0156_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2388_  (.A(\alu/_1016_ ),
    .B(\alu/_0156_ ),
    .Y(\alu/_0157_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_2389_  (.A(\alu/_0604_ ),
    .X(\alu/_0158_ ));
 sky130_fd_sc_hd__o2bb2a_1 \alu/_2390_  (.A1_N(\alu/_0602_ ),
    .A2_N(\alu/_0932_ ),
    .B1(\alu/_0603_ ),
    .B2(\alu/_0740_ ),
    .X(\alu/_0159_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2391_  (.A1(\alu/_0158_ ),
    .A2(\alu/_1135_ ),
    .B1(\alu/_0048_ ),
    .C1(\alu/_0159_ ),
    .X(\alu/_0160_ ));
 sky130_fd_sc_hd__and3_1 \alu/_2392_  (.A(\alu/_0155_ ),
    .B(\alu/_0157_ ),
    .C(\alu/_0160_ ),
    .X(\alu/_0161_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2393_  (.A1(\alu/_0118_ ),
    .A2(\alu/_0120_ ),
    .B1(\alu/_0158_ ),
    .X(\alu/_0162_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2394_  (.A(\alu/_0162_ ),
    .B(\alu/_0109_ ),
    .Y(\alu/_0163_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2395_  (.A1(\alu/_0158_ ),
    .A2(\alu/_0120_ ),
    .A3(\alu/_0118_ ),
    .B1(\alu/_0163_ ),
    .X(\alu/_0165_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2396_  (.A(\alu/_0129_ ),
    .B(\alu/_0607_ ),
    .Y(\alu/_0166_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2397_  (.A1(\alu/_0158_ ),
    .A2(\alu/_0166_ ),
    .B1(\alu/_1114_ ),
    .Y(\alu/_0167_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2398_  (.A1(\alu/_0158_ ),
    .A2(\alu/_0166_ ),
    .B1(\alu/_0167_ ),
    .X(\alu/_0168_ ));
 sky130_fd_sc_hd__nand3_4 \alu/_2399_  (.A(\alu/_0161_ ),
    .B(\alu/_0165_ ),
    .C(\alu/_0168_ ),
    .Y(\wAluOut[19] ));
 sky130_fd_sc_hd__nor2_1 \alu/_2400_  (.A(\alu/_0711_ ),
    .B(\alu/_1302_ ),
    .Y(\alu/_0169_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2401_  (.A0(\wAluA[20] ),
    .A1(\wAluA[19] ),
    .S(net229),
    .X(\alu/_0170_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2402_  (.A0(\alu/_0170_ ),
    .A1(\alu/_0133_ ),
    .S(net220),
    .X(\alu/_0171_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2403_  (.A0(\alu/_0171_ ),
    .A1(\alu/_0059_ ),
    .S(net187),
    .X(\alu/_0172_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2404_  (.A(net203),
    .B(\alu/_0172_ ),
    .Y(\alu/_0173_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2405_  (.A1(\alu/_0169_ ),
    .A2(\alu/_0173_ ),
    .B1(\alu/_0880_ ),
    .Y(\alu/_0175_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2406_  (.A1(\alu/_1034_ ),
    .A2(net171),
    .B1(\alu/_0976_ ),
    .Y(\alu/_0176_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2407_  (.A(\alu/_0175_ ),
    .B(\alu/_0176_ ),
    .Y(\alu/_0177_ ));
 sky130_fd_sc_hd__o2bb2a_1 \alu/_2408_  (.A1_N(\alu/_0640_ ),
    .A2_N(\alu/_0932_ ),
    .B1(\alu/_0641_ ),
    .B2(\alu/_1155_ ),
    .X(\alu/_0178_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2409_  (.A1(\alu/_0642_ ),
    .A2(\alu/_0893_ ),
    .B1(\alu/_0064_ ),
    .C1(\alu/_0178_ ),
    .X(\alu/_0179_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2410_  (.A(\alu/_0177_ ),
    .B(\alu/_0179_ ),
    .Y(\alu/_0180_ ));
 sky130_fd_sc_hd__a21oi_2 \alu/_2411_  (.A1(\alu/_1053_ ),
    .A2(\alu/_0144_ ),
    .B1(\alu/_0180_ ),
    .Y(\alu/_0181_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2412_  (.A(\alu/_0609_ ),
    .B(\alu/_0605_ ),
    .Y(\alu/_0182_ ));
 sky130_fd_sc_hd__nand2b_1 \alu/_2413_  (.A_N(\alu/_0182_ ),
    .B(\alu/_0113_ ),
    .Y(\alu/_0183_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2414_  (.A(\alu/_0183_ ),
    .Y(\alu/_0184_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2415_  (.A(\alu/_0084_ ),
    .B(\alu/_0184_ ),
    .Y(\alu/_0186_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_2416_  (.A1(\alu/_0120_ ),
    .A2(\alu/_0158_ ),
    .B1(\alu/_0603_ ),
    .X(\alu/_0187_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2417_  (.A1(\alu/_0182_ ),
    .A2(\alu/_0115_ ),
    .B1(\alu/_0187_ ),
    .Y(\alu/_0188_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2418_  (.A(\alu/_0188_ ),
    .Y(\alu/_0189_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2419_  (.A(\alu/_0186_ ),
    .B(\alu/_0189_ ),
    .Y(\alu/_0190_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2420_  (.A(\alu/_0190_ ),
    .Y(\alu/_0191_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2421_  (.A(\alu/_0642_ ),
    .B(\alu/_0191_ ),
    .Y(\alu/_0192_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2422_  (.A1(\alu/_0643_ ),
    .A2(\alu/_0190_ ),
    .B1(\alu/_1060_ ),
    .Y(\alu/_0193_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2423_  (.A(\alu/_0192_ ),
    .B(\alu/_0193_ ),
    .X(\alu/_0194_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2424_  (.A(\alu/_0786_ ),
    .Y(\alu/_0195_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2425_  (.A(\alu/_0622_ ),
    .Y(\alu/_0197_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2426_  (.A(\alu/_0777_ ),
    .B(\alu/_0197_ ),
    .Y(\alu/_0198_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2427_  (.A(\alu/_0198_ ),
    .B(\alu/_0195_ ),
    .Y(\alu/_0199_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2428_  (.A(\alu/_0199_ ),
    .B(\alu/_0642_ ),
    .Y(\alu/_0200_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2429_  (.A(\alu/_0200_ ),
    .B(\alu/_1193_ ),
    .Y(\alu/_0201_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2430_  (.A1(\alu/_0643_ ),
    .A2(\alu/_0195_ ),
    .A3(\alu/_0198_ ),
    .B1(\alu/_0201_ ),
    .X(\alu/_0202_ ));
 sky130_fd_sc_hd__nand3_2 \alu/_2431_  (.A(\alu/_0181_ ),
    .B(\alu/_0194_ ),
    .C(\alu/_0202_ ),
    .Y(\wAluOut[20] ));
 sky130_fd_sc_hd__mux2_2 \alu/_2432_  (.A0(\alu/_0632_ ),
    .A1(\alu/_0638_ ),
    .S(net224),
    .X(\alu/_0203_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2433_  (.A0(\alu/_0203_ ),
    .A1(\alu/_0146_ ),
    .S(net219),
    .X(\alu/_0204_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2434_  (.A0(\alu/_0204_ ),
    .A1(\alu/_0093_ ),
    .S(net189),
    .X(\alu/_0205_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2435_  (.A(\alu/_0205_ ),
    .B(\alu/_0711_ ),
    .Y(\alu/_0207_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2436_  (.A(\alu/_1329_ ),
    .B(net199),
    .Y(\alu/_0208_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2437_  (.A(\alu/_0207_ ),
    .B(\alu/_0208_ ),
    .C(\alu/_0879_ ),
    .Y(\alu/_0209_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2438_  (.A1(\alu/_0156_ ),
    .A2(\alu/_1090_ ),
    .B1(\alu/_0209_ ),
    .Y(\alu/_0210_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2439_  (.A(\alu/_0210_ ),
    .B(\alu/_0139_ ),
    .Y(\alu/_0211_ ));
 sky130_fd_sc_hd__o2bb2a_1 \alu/_2440_  (.A1_N(\alu/_0634_ ),
    .A2_N(\alu/_0932_ ),
    .B1(\alu/_0635_ ),
    .B2(\alu/_1155_ ),
    .X(\alu/_0212_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2441_  (.A1(\alu/_0664_ ),
    .A2(\alu/_0893_ ),
    .B1(\alu/_0064_ ),
    .C1(\alu/_0212_ ),
    .X(\alu/_0213_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2442_  (.A(\alu/_0211_ ),
    .B(\alu/_0213_ ),
    .Y(\alu/_0214_ ));
 sky130_fd_sc_hd__a21oi_2 \alu/_2443_  (.A1(\alu/_0144_ ),
    .A2(\alu/_1104_ ),
    .B1(\alu/_0214_ ),
    .Y(\alu/_0215_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2444_  (.A1(\alu/_0642_ ),
    .A2(\alu/_0191_ ),
    .B1(\alu/_0641_ ),
    .Y(\alu/_0216_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2445_  (.A(\alu/_0637_ ),
    .B(\alu/_0216_ ),
    .X(\alu/_0218_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2446_  (.A(\alu/_0216_ ),
    .B(\alu/_0637_ ),
    .Y(\alu/_0219_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2447_  (.A(\alu/_0218_ ),
    .B(\alu/_1177_ ),
    .C(\alu/_0219_ ),
    .Y(\alu/_0220_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2448_  (.A1(\alu/_0638_ ),
    .A2(\wAluB[20] ),
    .B1(\alu/_0200_ ),
    .Y(\alu/_0221_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2449_  (.A(\alu/_0664_ ),
    .B(\alu/_0221_ ),
    .X(\alu/_0222_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2450_  (.A(\alu/_0221_ ),
    .B(\alu/_0664_ ),
    .Y(\alu/_0223_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2451_  (.A(\alu/_0222_ ),
    .B(\alu/_0021_ ),
    .C(\alu/_0223_ ),
    .Y(\alu/_0224_ ));
 sky130_fd_sc_hd__nand3_2 \alu/_2452_  (.A(\alu/_0215_ ),
    .B(\alu/_0220_ ),
    .C(\alu/_0224_ ),
    .Y(\wAluOut[21] ));
 sky130_fd_sc_hd__inv_2 \alu/_2453_  (.A(\alu/_0788_ ),
    .Y(\alu/_0225_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2454_  (.A(\alu/_0199_ ),
    .B(\alu/_0644_ ),
    .Y(\alu/_0226_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2455_  (.A(\alu/_0226_ ),
    .B(\alu/_0225_ ),
    .Y(\alu/_0228_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2456_  (.A(\alu/_0630_ ),
    .Y(\alu/_0229_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2457_  (.A(\alu/_0228_ ),
    .B(\alu/_0229_ ),
    .Y(\alu/_0230_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2458_  (.A(\alu/_0230_ ),
    .B(\alu/_1193_ ),
    .Y(\alu/_0231_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2459_  (.A1(\alu/_0630_ ),
    .A2(\alu/_0225_ ),
    .A3(\alu/_0226_ ),
    .B1(\alu/_0231_ ),
    .X(\alu/_0232_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2460_  (.A1(\alu/_1132_ ),
    .A2(net172),
    .B1(\alu/_0976_ ),
    .X(\alu/_0233_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2461_  (.A0(net193),
    .A1(\wAluA[21] ),
    .S(net230),
    .X(\alu/_0234_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2462_  (.A0(\alu/_0234_ ),
    .A1(\alu/_0170_ ),
    .S(net219),
    .X(\alu/_0235_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2463_  (.A(\alu/_0235_ ),
    .B(\alu/_0870_ ),
    .Y(\alu/_0236_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2464_  (.A1(\alu/_0870_ ),
    .A2(\alu/_0136_ ),
    .B1(\alu/_0236_ ),
    .Y(\alu/_0237_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2465_  (.A(\alu/_0237_ ),
    .B(\alu/_1047_ ),
    .Y(\alu/_0239_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2466_  (.A(\alu/_0008_ ),
    .B(net203),
    .Y(\alu/_0240_ ));
 sky130_fd_sc_hd__and3_1 \alu/_2467_  (.A(\alu/_0239_ ),
    .B(\alu/_0240_ ),
    .C(\alu/_0879_ ),
    .X(\alu/_0241_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2468_  (.A(net193),
    .B(\wAluB[22] ),
    .Y(\alu/_0242_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2469_  (.A(net193),
    .B(\wAluB[22] ),
    .Y(\alu/_0243_ ));
 sky130_fd_sc_hd__clkbuf_2 \alu/_2470_  (.A(\alu/_0837_ ),
    .X(\alu/_0244_ ));
 sky130_fd_sc_hd__o22a_1 \alu/_2471_  (.A1(\alu/_0242_ ),
    .A2(\alu/_1083_ ),
    .B1(\alu/_0243_ ),
    .B2(\alu/_0244_ ),
    .X(\alu/_0245_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2472_  (.A1(\alu/_0229_ ),
    .A2(\alu/_1281_ ),
    .B1(\alu/_0049_ ),
    .C1(\alu/_0245_ ),
    .X(\alu/_0246_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2473_  (.A1(\alu/_0233_ ),
    .A2(\alu/_0241_ ),
    .B1(\alu/_0246_ ),
    .Y(\alu/_0247_ ));
 sky130_fd_sc_hd__a21oi_2 \alu/_2474_  (.A1(\alu/_1125_ ),
    .A2(\alu/_0880_ ),
    .B1(\alu/_0247_ ),
    .Y(\alu/_0248_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2475_  (.A(\alu/_0636_ ),
    .B(\alu/_0642_ ),
    .Y(\alu/_0250_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2476_  (.A(\alu/_0190_ ),
    .B(\alu/_0250_ ),
    .Y(\alu/_0251_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_2477_  (.A1(\alu/_0641_ ),
    .A2(\alu/_0664_ ),
    .B1(\alu/_0635_ ),
    .X(\alu/_0252_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2478_  (.A(\alu/_0251_ ),
    .B(\alu/_0252_ ),
    .Y(\alu/_0253_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2479_  (.A(\alu/_0253_ ),
    .B(\alu/_0630_ ),
    .Y(\alu/_0254_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2480_  (.A(\alu/_0254_ ),
    .B(\alu/_0109_ ),
    .Y(\alu/_0255_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2481_  (.A1(\alu/_0229_ ),
    .A2(\alu/_0251_ ),
    .A3(\alu/_0252_ ),
    .B1(\alu/_0255_ ),
    .X(\alu/_0256_ ));
 sky130_fd_sc_hd__nand3_2 \alu/_2482_  (.A(\alu/_0232_ ),
    .B(\alu/_0248_ ),
    .C(\alu/_0256_ ),
    .Y(\wAluOut[22] ));
 sky130_fd_sc_hd__nor2_1 \alu/_2483_  (.A(net171),
    .B(\alu/_1170_ ),
    .Y(\alu/_0257_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2484_  (.A1(\alu/_1153_ ),
    .A2(net172),
    .B1(\alu/_0976_ ),
    .X(\alu/_0258_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2485_  (.A0(\wAluA[23] ),
    .A1(\wAluA[22] ),
    .S(net231),
    .X(\alu/_0260_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2486_  (.A(\alu/_0203_ ),
    .B(net214),
    .Y(\alu/_0261_ ));
 sky130_fd_sc_hd__o21ai_2 \alu/_2487_  (.A1(net214),
    .A2(\alu/_0260_ ),
    .B1(\alu/_0261_ ),
    .Y(\alu/_0262_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2488_  (.A(\alu/_0148_ ),
    .B(net187),
    .Y(\alu/_0263_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2489_  (.A1(net187),
    .A2(\alu/_0262_ ),
    .B1(\alu/_0263_ ),
    .Y(\alu/_0264_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2490_  (.A(net203),
    .B(\alu/_0264_ ),
    .Y(\alu/_0265_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2491_  (.A(\alu/_0947_ ),
    .B(\alu/_0043_ ),
    .Y(\alu/_0266_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_2492_  (.A1(\alu/_0265_ ),
    .A2(\alu/_0266_ ),
    .B1(\alu/_0156_ ),
    .X(\alu/_0267_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2493_  (.A(\alu/_0663_ ),
    .Y(\alu/_0268_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2494_  (.A(\wAluA[23] ),
    .B(\wAluB[23] ),
    .Y(\alu/_0269_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2495_  (.A(\wAluA[23] ),
    .B(\wAluB[23] ),
    .Y(\alu/_0271_ ));
 sky130_fd_sc_hd__o22a_1 \alu/_2496_  (.A1(\alu/_0269_ ),
    .A2(\alu/_0244_ ),
    .B1(\alu/_0271_ ),
    .B2(\alu/_1134_ ),
    .X(\alu/_0272_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2497_  (.A1(\alu/_0268_ ),
    .A2(\alu/_0893_ ),
    .B1(\alu/_0064_ ),
    .C1(\alu/_0272_ ),
    .X(\alu/_0273_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2498_  (.A1(\alu/_0258_ ),
    .A2(\alu/_0267_ ),
    .B1(\alu/_0273_ ),
    .Y(\alu/_0274_ ));
 sky130_fd_sc_hd__nor2_2 \alu/_2499_  (.A(\alu/_0257_ ),
    .B(\alu/_0274_ ),
    .Y(\alu/_0275_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2500_  (.A(\alu/_0230_ ),
    .B(\alu/_0628_ ),
    .Y(\alu/_0276_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2501_  (.A(\alu/_0268_ ),
    .B(\alu/_0276_ ),
    .X(\alu/_0277_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2502_  (.A(\alu/_0276_ ),
    .B(\alu/_0268_ ),
    .Y(\alu/_0278_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2503_  (.A(\alu/_0277_ ),
    .B(\alu/_0021_ ),
    .C(\alu/_0278_ ),
    .Y(\alu/_0279_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2504_  (.A(\alu/_0254_ ),
    .B(\alu/_0242_ ),
    .Y(\alu/_0280_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2505_  (.A(\alu/_0663_ ),
    .B(\alu/_0280_ ),
    .X(\alu/_0282_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2506_  (.A(\alu/_0280_ ),
    .B(\alu/_0663_ ),
    .Y(\alu/_0283_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2507_  (.A(\alu/_0282_ ),
    .B(\alu/_0028_ ),
    .C(\alu/_0283_ ),
    .Y(\alu/_0284_ ));
 sky130_fd_sc_hd__nand3_4 \alu/_2508_  (.A(\alu/_0275_ ),
    .B(\alu/_0279_ ),
    .C(\alu/_0284_ ),
    .Y(\wAluOut[23] ));
 sky130_fd_sc_hd__mux2_2 \alu/_2509_  (.A0(\alu/_0561_ ),
    .A1(\alu/_0623_ ),
    .S(net235),
    .X(\alu/_0285_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2510_  (.A(\alu/_0234_ ),
    .B(net219),
    .Y(\alu/_0286_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2511_  (.A1(net218),
    .A2(\alu/_0285_ ),
    .B1(\alu/_0286_ ),
    .Y(\alu/_0287_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2512_  (.A0(\alu/_0171_ ),
    .A1(\alu/_0287_ ),
    .S(\alu/_0704_ ),
    .X(\alu/_0288_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2513_  (.A0(\alu/_0060_ ),
    .A1(\alu/_0288_ ),
    .S(\alu/_0946_ ),
    .X(\alu/_0289_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2514_  (.A(\alu/_0289_ ),
    .B(\alu/_1018_ ),
    .Y(\alu/_0290_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2515_  (.A(\alu/_0548_ ),
    .B(\alu/_0976_ ),
    .Y(\alu/_0292_ ));
 sky130_fd_sc_hd__buf_4 \alu/_2516_  (.A(\alu/_0292_ ),
    .X(\alu/_0293_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2517_  (.A(\alu/_1183_ ),
    .B(\alu/_0293_ ),
    .Y(\alu/_0294_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2518_  (.A(\wAluA[24] ),
    .B(\wAluB[24] ),
    .Y(\alu/_0295_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2519_  (.A(\wAluA[24] ),
    .B(\wAluB[24] ),
    .Y(\alu/_0296_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2520_  (.A(\alu/_0564_ ),
    .Y(\alu/_0297_ ));
 sky130_fd_sc_hd__o22a_1 \alu/_2521_  (.A1(\alu/_0296_ ),
    .A2(\alu/_0837_ ),
    .B1(\alu/_0297_ ),
    .B2(\alu/_0928_ ),
    .X(\alu/_0298_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2522_  (.A1(\alu/_0295_ ),
    .A2(\alu/_1134_ ),
    .B1(\alu/_0048_ ),
    .C1(\alu/_0298_ ),
    .X(\alu/_0299_ ));
 sky130_fd_sc_hd__and3_1 \alu/_2523_  (.A(\alu/_0290_ ),
    .B(\alu/_0294_ ),
    .C(\alu/_0299_ ),
    .X(\alu/_0300_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2524_  (.A(\alu/_1197_ ),
    .B(\alu/_0144_ ),
    .Y(\alu/_0301_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2525_  (.A(\alu/_0793_ ),
    .B(\alu/_0297_ ),
    .Y(\alu/_0303_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2526_  (.A(\alu/_0297_ ),
    .B(\alu/_0793_ ),
    .X(\alu/_0304_ ));
 sky130_fd_sc_hd__and3_1 \alu/_2527_  (.A(\alu/_0250_ ),
    .B(\alu/_0626_ ),
    .C(\alu/_0630_ ),
    .X(\alu/_0305_ ));
 sky130_fd_sc_hd__and2_1 \alu/_2528_  (.A(\alu/_0184_ ),
    .B(\alu/_0305_ ),
    .X(\alu/_0306_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2529_  (.A(\alu/_0084_ ),
    .B(\alu/_0306_ ),
    .Y(\alu/_0307_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2530_  (.A(\alu/_0663_ ),
    .B(\alu/_0630_ ),
    .Y(\alu/_0308_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2531_  (.A1(\alu/_0271_ ),
    .A2(\alu/_0242_ ),
    .B1(\alu/_0269_ ),
    .X(\alu/_0309_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2532_  (.A1(\alu/_0308_ ),
    .A2(\alu/_0252_ ),
    .B1(\alu/_0309_ ),
    .Y(\alu/_0310_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2533_  (.A1(\alu/_0188_ ),
    .A2(\alu/_0305_ ),
    .B1(\alu/_0310_ ),
    .Y(\alu/_0311_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_2534_  (.A(\alu/_0307_ ),
    .B(\alu/_0311_ ),
    .Y(\alu/_0312_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2535_  (.A(\alu/_0564_ ),
    .B(\alu/_0312_ ),
    .X(\alu/_0314_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2536_  (.A(\alu/_0312_ ),
    .B(\alu/_0564_ ),
    .Y(\alu/_0315_ ));
 sky130_fd_sc_hd__and3_1 \alu/_2537_  (.A(\alu/_0314_ ),
    .B(\alu/_1060_ ),
    .C(\alu/_0315_ ),
    .X(\alu/_0316_ ));
 sky130_fd_sc_hd__a31oi_2 \alu/_2538_  (.A1(\alu/_1055_ ),
    .A2(\alu/_0303_ ),
    .A3(\alu/_0304_ ),
    .B1(\alu/_0316_ ),
    .Y(\alu/_0317_ ));
 sky130_fd_sc_hd__nand3_4 \alu/_2539_  (.A(\alu/_0300_ ),
    .B(\alu/_0301_ ),
    .C(\alu/_0317_ ),
    .Y(\wAluOut[24] ));
 sky130_fd_sc_hd__mux2_1 \alu/_2540_  (.A0(\alu/_0555_ ),
    .A1(\alu/_0561_ ),
    .S(net224),
    .X(\alu/_0318_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2541_  (.A(\alu/_0260_ ),
    .B(net214),
    .Y(\alu/_0319_ ));
 sky130_fd_sc_hd__o21ai_2 \alu/_2542_  (.A1(net214),
    .A2(\alu/_0318_ ),
    .B1(\alu/_0319_ ),
    .Y(\alu/_0320_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2543_  (.A(\alu/_0818_ ),
    .B(\alu/_0204_ ),
    .Y(\alu/_0321_ ));
 sky130_fd_sc_hd__a211o_1 \alu/_2544_  (.A1(\alu/_0705_ ),
    .A2(\alu/_0320_ ),
    .B1(net204),
    .C1(\alu/_0321_ ),
    .X(\alu/_0322_ ));
 sky130_fd_sc_hd__o211ai_2 \alu/_2545_  (.A1(\alu/_0721_ ),
    .A2(\alu/_0095_ ),
    .B1(\alu/_1332_ ),
    .C1(\alu/_0322_ ),
    .Y(\alu/_0324_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \alu/_2546_  (.A(\alu/_0559_ ),
    .X(\alu/_0325_ ));
 sky130_fd_sc_hd__o2bb2a_1 \alu/_2547_  (.A1_N(\alu/_0557_ ),
    .A2_N(\alu/_0932_ ),
    .B1(\alu/_0558_ ),
    .B2(\alu/_1155_ ),
    .X(\alu/_0326_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2548_  (.A1(\alu/_0325_ ),
    .A2(\alu/_1281_ ),
    .B1(\alu/_0049_ ),
    .C1(\alu/_0326_ ),
    .X(\alu/_0327_ ));
 sky130_fd_sc_hd__o211ai_2 \alu/_2549_  (.A1(\alu/_0721_ ),
    .A2(\alu/_1212_ ),
    .B1(\alu/_0293_ ),
    .C1(\alu/_1217_ ),
    .Y(\alu/_0328_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2550_  (.A(\alu/_0324_ ),
    .B(\alu/_0327_ ),
    .C(\alu/_0328_ ),
    .Y(\alu/_0329_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2551_  (.A1(\alu/_0144_ ),
    .A2(\alu/_1228_ ),
    .B1(\alu/_0329_ ),
    .Y(\alu/_0330_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2552_  (.A1(\alu/_0315_ ),
    .A2(\alu/_0295_ ),
    .B1(\alu/_0325_ ),
    .X(\alu/_0331_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2553_  (.A(\alu/_0331_ ),
    .B(\alu/_0109_ ),
    .Y(\alu/_0332_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2554_  (.A1(\alu/_0325_ ),
    .A2(\alu/_0295_ ),
    .A3(\alu/_0315_ ),
    .B1(\alu/_0332_ ),
    .X(\alu/_0333_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2555_  (.A(\alu/_0303_ ),
    .B(\alu/_0562_ ),
    .Y(\alu/_0335_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2556_  (.A1(\alu/_0325_ ),
    .A2(\alu/_0335_ ),
    .B1(\alu/_1114_ ),
    .Y(\alu/_0336_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2557_  (.A1(\alu/_0325_ ),
    .A2(\alu/_0335_ ),
    .B1(\alu/_0336_ ),
    .X(\alu/_0337_ ));
 sky130_fd_sc_hd__nand3_2 \alu/_2558_  (.A(\alu/_0330_ ),
    .B(\alu/_0333_ ),
    .C(\alu/_0337_ ),
    .Y(\wAluOut[25] ));
 sky130_fd_sc_hd__mux2_2 \alu/_2559_  (.A0(\alu/_0571_ ),
    .A1(\alu/_0555_ ),
    .S(net224),
    .X(\alu/_0338_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2560_  (.A0(\alu/_0338_ ),
    .A1(\alu/_0285_ ),
    .S(net218),
    .X(\alu/_0339_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2561_  (.A1(\alu/_0339_ ),
    .A2(\alu/_0818_ ),
    .B1(net205),
    .Y(\alu/_0340_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2562_  (.A(\alu/_0817_ ),
    .B(\alu/_0235_ ),
    .X(\alu/_0341_ ));
 sky130_fd_sc_hd__a22o_1 \alu/_2563_  (.A1(\alu/_0340_ ),
    .A2(\alu/_0341_ ),
    .B1(\alu/_0138_ ),
    .B2(net206),
    .X(\alu/_0342_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2564_  (.A(\alu/_0342_ ),
    .B(\alu/_1332_ ),
    .Y(\alu/_0343_ ));
 sky130_fd_sc_hd__o211ai_2 \alu/_2565_  (.A1(\alu/_0721_ ),
    .A2(\alu/_0981_ ),
    .B1(\alu/_0293_ ),
    .C1(\alu/_1242_ ),
    .Y(\alu/_0345_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2566_  (.A(\alu/_0575_ ),
    .Y(\alu/_0346_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2567_  (.A(\wAluA[26] ),
    .B(\wAluB[26] ),
    .Y(\alu/_0347_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2568_  (.A(\wAluA[26] ),
    .B(\wAluB[26] ),
    .Y(\alu/_0348_ ));
 sky130_fd_sc_hd__o22a_1 \alu/_2569_  (.A1(\alu/_0347_ ),
    .A2(\alu/_1155_ ),
    .B1(\alu/_0348_ ),
    .B2(\alu/_0244_ ),
    .X(\alu/_0349_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2570_  (.A1(\alu/_0346_ ),
    .A2(\alu/_1281_ ),
    .B1(\alu/_0049_ ),
    .C1(\alu/_0349_ ),
    .X(\alu/_0350_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2571_  (.A(\alu/_0343_ ),
    .B(\alu/_0345_ ),
    .C(\alu/_0350_ ),
    .Y(\alu/_0351_ ));
 sky130_fd_sc_hd__a21oi_2 \alu/_2572_  (.A1(\alu/_0144_ ),
    .A2(\alu/_1250_ ),
    .B1(\alu/_0351_ ),
    .Y(\alu/_0352_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2573_  (.A(\alu/_0795_ ),
    .Y(\alu/_0353_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2574_  (.A(\alu/_0793_ ),
    .B(\alu/_0565_ ),
    .Y(\alu/_0354_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2575_  (.A(\alu/_0354_ ),
    .B(\alu/_0353_ ),
    .Y(\alu/_0356_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2576_  (.A(\alu/_0356_ ),
    .B(\alu/_0346_ ),
    .Y(\alu/_0357_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2577_  (.A(\alu/_0357_ ),
    .B(\alu/_0896_ ),
    .Y(\alu/_0358_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2578_  (.A1(\alu/_0575_ ),
    .A2(\alu/_0353_ ),
    .A3(\alu/_0354_ ),
    .B1(\alu/_0358_ ),
    .X(\alu/_0359_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_2579_  (.A1(\alu/_0295_ ),
    .A2(\alu/_0559_ ),
    .B1(\alu/_0558_ ),
    .X(\alu/_0360_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2580_  (.A(\alu/_0325_ ),
    .B(\alu/_0297_ ),
    .Y(\alu/_0361_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2581_  (.A(\alu/_0312_ ),
    .B(\alu/_0361_ ),
    .Y(\alu/_0362_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2582_  (.A(\alu/_0362_ ),
    .B(\alu/_0360_ ),
    .Y(\alu/_0363_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2583_  (.A(\alu/_0363_ ),
    .B(\alu/_0575_ ),
    .Y(\alu/_0364_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2584_  (.A(\alu/_0364_ ),
    .B(\alu/_0109_ ),
    .Y(\alu/_0365_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2585_  (.A1(\alu/_0346_ ),
    .A2(\alu/_0360_ ),
    .A3(\alu/_0362_ ),
    .B1(\alu/_0365_ ),
    .X(\alu/_0367_ ));
 sky130_fd_sc_hd__nand3_4 \alu/_2586_  (.A(\alu/_0352_ ),
    .B(\alu/_0359_ ),
    .C(\alu/_0367_ ),
    .Y(\wAluOut[26] ));
 sky130_fd_sc_hd__nand2_1 \alu/_2587_  (.A(\alu/_0357_ ),
    .B(\alu/_0573_ ),
    .Y(\alu/_0368_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2588_  (.A(\alu/_0794_ ),
    .B(\alu/_0368_ ),
    .X(\alu/_0369_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2589_  (.A(\alu/_0368_ ),
    .B(\alu/_0794_ ),
    .Y(\alu/_0370_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2590_  (.A(\alu/_0369_ ),
    .B(\alu/_0021_ ),
    .C(\alu/_0370_ ),
    .Y(\alu/_0371_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2591_  (.A(\alu/_1279_ ),
    .B(\alu/_0293_ ),
    .Y(\alu/_0372_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2592_  (.A0(\wAluA[27] ),
    .A1(\wAluA[26] ),
    .S(net230),
    .X(\alu/_0373_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2593_  (.A(\alu/_0318_ ),
    .B(net215),
    .Y(\alu/_0374_ ));
 sky130_fd_sc_hd__o21ai_2 \alu/_2594_  (.A1(net215),
    .A2(\alu/_0373_ ),
    .B1(\alu/_0374_ ),
    .Y(\alu/_0375_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2595_  (.A1(\alu/_0262_ ),
    .A2(net188),
    .B1(net206),
    .X(\alu/_0377_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2596_  (.A1(\alu/_0705_ ),
    .A2(\alu/_0375_ ),
    .B1(\alu/_0377_ ),
    .Y(\alu/_0378_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2597_  (.A(\alu/_0832_ ),
    .B(\alu/_0150_ ),
    .Y(\alu/_0379_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2598_  (.A1(\alu/_0378_ ),
    .A2(\alu/_0379_ ),
    .B1(\alu/_1332_ ),
    .Y(\alu/_0380_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2599_  (.A(\wAluA[27] ),
    .B(\wAluB[27] ),
    .Y(\alu/_0381_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2600_  (.A(\wAluA[27] ),
    .B(\wAluB[27] ),
    .Y(\alu/_0382_ ));
 sky130_fd_sc_hd__o22a_1 \alu/_2601_  (.A1(\alu/_0381_ ),
    .A2(\alu/_1155_ ),
    .B1(\alu/_0382_ ),
    .B2(\alu/_0244_ ),
    .X(\alu/_0383_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2602_  (.A1(\alu/_0794_ ),
    .A2(\alu/_1281_ ),
    .B1(\alu/_0049_ ),
    .C1(\alu/_0383_ ),
    .X(\alu/_0384_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2603_  (.A(\alu/_0372_ ),
    .B(\alu/_0380_ ),
    .C(\alu/_0384_ ),
    .Y(\alu/_0385_ ));
 sky130_fd_sc_hd__a21oi_2 \alu/_2604_  (.A1(\alu/_1272_ ),
    .A2(\alu/_0880_ ),
    .B1(\alu/_0385_ ),
    .Y(\alu/_0386_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2605_  (.A(\alu/_0364_ ),
    .B(\alu/_0347_ ),
    .Y(\alu/_0388_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2606_  (.A(\alu/_0570_ ),
    .B(\alu/_0388_ ),
    .X(\alu/_0389_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2607_  (.A(\alu/_0388_ ),
    .B(\alu/_0570_ ),
    .Y(\alu/_0390_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2608_  (.A(\alu/_0389_ ),
    .B(\alu/_0028_ ),
    .C(\alu/_0390_ ),
    .Y(\alu/_0391_ ));
 sky130_fd_sc_hd__nand3_2 \alu/_2609_  (.A(\alu/_0371_ ),
    .B(\alu/_0386_ ),
    .C(\alu/_0391_ ),
    .Y(\wAluOut[27] ));
 sky130_fd_sc_hd__o21a_1 \alu/_2610_  (.A1(\alu/_0692_ ),
    .A2(\alu/_0566_ ),
    .B1(\alu/_0811_ ),
    .X(\alu/_0392_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2611_  (.A1(\alu/_0392_ ),
    .A2(\alu/_0826_ ),
    .B1(net187),
    .X(\alu/_0393_ ));
 sky130_fd_sc_hd__a21oi_1 \alu/_2612_  (.A1(\alu/_0338_ ),
    .A2(net218),
    .B1(\alu/_0393_ ),
    .Y(\alu/_0394_ ));
 sky130_fd_sc_hd__a211o_1 \alu/_2613_  (.A1(\alu/_0287_ ),
    .A2(net187),
    .B1(net203),
    .C1(\alu/_0394_ ),
    .X(\alu/_0395_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2614_  (.A1(\alu/_0986_ ),
    .A2(\alu/_0172_ ),
    .B1(\alu/_0883_ ),
    .C1(\alu/_0395_ ),
    .X(\alu/_0396_ ));
 sky130_fd_sc_hd__and2_1 \alu/_2615_  (.A(\alu/_1309_ ),
    .B(\alu/_0156_ ),
    .X(\alu/_0398_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2616_  (.A(\alu/_1303_ ),
    .B(\alu/_0293_ ),
    .Y(\alu/_0399_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2617_  (.A(\alu/_0596_ ),
    .Y(\alu/_0400_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2618_  (.A(net236),
    .B(\wAluB[28] ),
    .Y(\alu/_0401_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2619_  (.A(net236),
    .B(\wAluB[28] ),
    .Y(\alu/_0402_ ));
 sky130_fd_sc_hd__o22a_1 \alu/_2620_  (.A1(\alu/_0401_ ),
    .A2(\alu/_1083_ ),
    .B1(\alu/_0402_ ),
    .B2(\alu/_0244_ ),
    .X(\alu/_0403_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2621_  (.A1(\alu/_0400_ ),
    .A2(\alu/_1281_ ),
    .B1(\alu/_0049_ ),
    .C1(\alu/_0403_ ),
    .X(\alu/_0404_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2622_  (.A(\alu/_0399_ ),
    .B(\alu/_0404_ ),
    .Y(\alu/_0405_ ));
 sky130_fd_sc_hd__nor3_2 \alu/_2623_  (.A(\alu/_0396_ ),
    .B(\alu/_0398_ ),
    .C(\alu/_0405_ ),
    .Y(\alu/_0406_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2624_  (.A(\alu/_0577_ ),
    .Y(\alu/_0407_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2625_  (.A(\alu/_0793_ ),
    .B(\alu/_0407_ ),
    .Y(\alu/_0409_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2626_  (.A(\alu/_0409_ ),
    .B(\alu/_0796_ ),
    .Y(\alu/_0410_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2627_  (.A(\alu/_0410_ ),
    .B(\alu/_0400_ ),
    .Y(\alu/_0411_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2628_  (.A(\alu/_0411_ ),
    .B(\alu/_0896_ ),
    .Y(\alu/_0412_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2629_  (.A1(\alu/_0596_ ),
    .A2(\alu/_0796_ ),
    .A3(\alu/_0409_ ),
    .B1(\alu/_0412_ ),
    .X(\alu/_0413_ ));
 sky130_fd_sc_hd__and3_1 \alu/_2630_  (.A(\alu/_0361_ ),
    .B(\alu/_0570_ ),
    .C(\alu/_0575_ ),
    .X(\alu/_0414_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2631_  (.A(\alu/_0312_ ),
    .B(\alu/_0414_ ),
    .Y(\alu/_0415_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2632_  (.A(\alu/_0570_ ),
    .B(\alu/_0575_ ),
    .Y(\alu/_0416_ ));
 sky130_fd_sc_hd__o221a_1 \alu/_2633_  (.A1(\alu/_0794_ ),
    .A2(\alu/_0347_ ),
    .B1(\alu/_0416_ ),
    .B2(\alu/_0360_ ),
    .C1(\alu/_0381_ ),
    .X(\alu/_0417_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2634_  (.A(\alu/_0415_ ),
    .B(\alu/_0417_ ),
    .Y(\alu/_0418_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2635_  (.A(\alu/_0418_ ),
    .B(\alu/_0596_ ),
    .Y(\alu/_0420_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2636_  (.A(\alu/_0420_ ),
    .B(\alu/_0109_ ),
    .Y(\alu/_0421_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2637_  (.A1(\alu/_0400_ ),
    .A2(\alu/_0415_ ),
    .A3(\alu/_0417_ ),
    .B1(\alu/_0421_ ),
    .X(\alu/_0422_ ));
 sky130_fd_sc_hd__nand3_4 \alu/_2638_  (.A(\alu/_0406_ ),
    .B(\alu/_0413_ ),
    .C(\alu/_0422_ ),
    .Y(\wAluOut[28] ));
 sky130_fd_sc_hd__a22oi_1 \alu/_2639_  (.A1(\alu/_1315_ ),
    .A2(\alu/_0156_ ),
    .B1(\alu/_1331_ ),
    .B2(\alu/_0293_ ),
    .Y(\alu/_0423_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2640_  (.A0(\wAluA[29] ),
    .A1(net236),
    .S(net230),
    .X(\alu/_0424_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2641_  (.A0(\alu/_0424_ ),
    .A1(\alu/_0373_ ),
    .S(net215),
    .X(\alu/_0425_ ));
 sky130_fd_sc_hd__mux2_1 \alu/_2642_  (.A0(\alu/_0425_ ),
    .A1(\alu/_0320_ ),
    .S(net185),
    .X(\alu/_0426_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2643_  (.A(\alu/_0205_ ),
    .B(net202),
    .Y(\alu/_0427_ ));
 sky130_fd_sc_hd__o211ai_1 \alu/_2644_  (.A1(net201),
    .A2(\alu/_0426_ ),
    .B1(\alu/_0883_ ),
    .C1(\alu/_0427_ ),
    .Y(\alu/_0428_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2645_  (.A(\alu/_0592_ ),
    .Y(\alu/_0430_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2646_  (.A(\wAluA[29] ),
    .B(\wAluB[29] ),
    .Y(\alu/_0431_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2647_  (.A(\wAluA[29] ),
    .B(\wAluB[29] ),
    .Y(\alu/_0432_ ));
 sky130_fd_sc_hd__o22a_1 \alu/_2648_  (.A1(\alu/_0431_ ),
    .A2(\alu/_0740_ ),
    .B1(\alu/_0432_ ),
    .B2(\alu/_0837_ ),
    .X(\alu/_0433_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2649_  (.A1(\alu/_0430_ ),
    .A2(\alu/_1135_ ),
    .B1(\alu/_0048_ ),
    .C1(\alu/_0433_ ),
    .X(\alu/_0434_ ));
 sky130_fd_sc_hd__and3_1 \alu/_2650_  (.A(\alu/_0423_ ),
    .B(\alu/_0428_ ),
    .C(\alu/_0434_ ),
    .X(\alu/_0435_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2651_  (.A(\alu/_0411_ ),
    .B(\alu/_0595_ ),
    .Y(\alu/_0436_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2652_  (.A(\alu/_0430_ ),
    .B(\alu/_0436_ ),
    .X(\alu/_0437_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2653_  (.A(\alu/_0436_ ),
    .B(\alu/_0430_ ),
    .Y(\alu/_0438_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2654_  (.A(\alu/_0437_ ),
    .B(\alu/_1055_ ),
    .C(\alu/_0438_ ),
    .Y(\alu/_0439_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2655_  (.A(\alu/_0420_ ),
    .B(\alu/_0401_ ),
    .Y(\alu/_0441_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2656_  (.A(\alu/_0592_ ),
    .B(\alu/_0441_ ),
    .X(\alu/_0442_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2657_  (.A(\alu/_0441_ ),
    .B(\alu/_0592_ ),
    .Y(\alu/_0443_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2658_  (.A(\alu/_0442_ ),
    .B(\alu/_0028_ ),
    .C(\alu/_0443_ ),
    .Y(\alu/_0444_ ));
 sky130_fd_sc_hd__nand3_4 \alu/_2659_  (.A(\alu/_0435_ ),
    .B(\alu/_0439_ ),
    .C(\alu/_0444_ ),
    .Y(\wAluOut[29] ));
 sky130_fd_sc_hd__a31o_1 \alu/_2660_  (.A1(\alu/_0809_ ),
    .A2(\alu/_0812_ ),
    .A3(\alu/_0822_ ),
    .B1(net188),
    .X(\alu/_0445_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2661_  (.A1(net218),
    .A2(\alu/_0392_ ),
    .B1(\alu/_0445_ ),
    .X(\alu/_0446_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2662_  (.A(\alu/_0446_ ),
    .B(\alu/_1047_ ),
    .Y(\alu/_0447_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2663_  (.A(\alu/_0705_ ),
    .B(\alu/_0339_ ),
    .Y(\alu/_0448_ ));
 sky130_fd_sc_hd__o221ai_1 \alu/_2664_  (.A1(\alu/_0447_ ),
    .A2(\alu/_0448_ ),
    .B1(\alu/_1226_ ),
    .B2(\alu/_0237_ ),
    .C1(\alu/_0883_ ),
    .Y(\alu/_0449_ ));
 sky130_fd_sc_hd__o211ai_1 \alu/_2665_  (.A1(net203),
    .A2(\alu/_0008_ ),
    .B1(\alu/_0292_ ),
    .C1(\alu/_0009_ ),
    .Y(\alu/_0451_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2666_  (.A(\alu/_0587_ ),
    .Y(\alu/_0452_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2667_  (.A(\wAluA[30] ),
    .B(\wAluB[30] ),
    .Y(\alu/_0453_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2668_  (.A(\wAluA[30] ),
    .B(\wAluB[30] ),
    .Y(\alu/_0454_ ));
 sky130_fd_sc_hd__o22a_1 \alu/_2669_  (.A1(\alu/_0453_ ),
    .A2(\alu/_0740_ ),
    .B1(\alu/_0454_ ),
    .B2(\alu/_0837_ ),
    .X(\alu/_0455_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2670_  (.A1(\alu/_0452_ ),
    .A2(\alu/_0928_ ),
    .B1(\alu/_0048_ ),
    .C1(\alu/_0455_ ),
    .X(\alu/_0456_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2671_  (.A(\alu/_0012_ ),
    .B(\alu/_0156_ ),
    .Y(\alu/_0457_ ));
 sky130_fd_sc_hd__and4_1 \alu/_2672_  (.A(\alu/_0449_ ),
    .B(\alu/_0451_ ),
    .C(\alu/_0456_ ),
    .D(\alu/_0457_ ),
    .X(\alu/_0458_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2673_  (.A(\alu/_0410_ ),
    .B(\alu/_0597_ ),
    .Y(\alu/_0459_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2674_  (.A(\alu/_0459_ ),
    .B(\alu/_0797_ ),
    .Y(\alu/_0460_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2675_  (.A(\alu/_0452_ ),
    .B(\alu/_0460_ ),
    .X(\alu/_0462_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2676_  (.A(\alu/_0460_ ),
    .B(\alu/_0452_ ),
    .Y(\alu/_0463_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2677_  (.A(\alu/_0462_ ),
    .B(\alu/_1055_ ),
    .C(\alu/_0463_ ),
    .Y(\alu/_0464_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2678_  (.A(\alu/_0430_ ),
    .B(\alu/_0400_ ),
    .Y(\alu/_0465_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2679_  (.A(\alu/_0418_ ),
    .B(\alu/_0465_ ),
    .Y(\alu/_0466_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2680_  (.A1(\alu/_0431_ ),
    .A2(\alu/_0401_ ),
    .B1(\alu/_0432_ ),
    .X(\alu/_0467_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2681_  (.A(\alu/_0466_ ),
    .B(\alu/_0467_ ),
    .Y(\alu/_0468_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2682_  (.A(\alu/_0587_ ),
    .B(\alu/_0468_ ),
    .X(\alu/_0469_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2683_  (.A(\alu/_0468_ ),
    .B(\alu/_0587_ ),
    .Y(\alu/_0470_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2684_  (.A(\alu/_0469_ ),
    .B(\alu/_0028_ ),
    .C(\alu/_0470_ ),
    .Y(\alu/_0471_ ));
 sky130_fd_sc_hd__nand3_4 \alu/_2685_  (.A(\alu/_0458_ ),
    .B(\alu/_0464_ ),
    .C(\alu/_0471_ ),
    .Y(\wAluOut[30] ));
 sky130_fd_sc_hd__inv_2 \alu/_2686_  (.A(\alu/_0585_ ),
    .Y(\alu/_0473_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2687_  (.A(\alu/_0463_ ),
    .B(\alu/_0473_ ),
    .Y(\alu/_0474_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2688_  (.A(\alu/_0474_ ),
    .B(\alu/_0582_ ),
    .Y(\alu/_0475_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2689_  (.A(\alu/_0463_ ),
    .B(\alu/_0583_ ),
    .C(\alu/_0473_ ),
    .Y(\alu/_0476_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2690_  (.A(\alu/_0475_ ),
    .B(\alu/_0021_ ),
    .C(\alu/_0476_ ),
    .Y(\alu/_0477_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2691_  (.A(\alu/_0424_ ),
    .B(net215),
    .Y(\alu/_0478_ ));
 sky130_fd_sc_hd__o21a_1 \alu/_2692_  (.A1(net219),
    .A2(\alu/_0843_ ),
    .B1(\alu/_0816_ ),
    .X(\alu/_0479_ ));
 sky130_fd_sc_hd__a32o_1 \alu/_2693_  (.A1(\alu/_0478_ ),
    .A2(\alu/_1006_ ),
    .A3(\alu/_0479_ ),
    .B1(\alu/_0375_ ),
    .B2(net184),
    .X(\alu/_0480_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2694_  (.A(\alu/_0946_ ),
    .B(\alu/_0264_ ),
    .Y(\alu/_0481_ ));
 sky130_fd_sc_hd__a211o_1 \alu/_2695_  (.A1(\alu/_0480_ ),
    .A2(\alu/_0831_ ),
    .B1(\alu/_0747_ ),
    .C1(\alu/_0481_ ),
    .X(\alu/_0483_ ));
 sky130_fd_sc_hd__nor2_1 \alu/_2696_  (.A(net192),
    .B(\wAluB[31] ),
    .Y(\alu/_0484_ ));
 sky130_fd_sc_hd__or3_1 \alu/_2697_  (.A(\alu/_0912_ ),
    .B(\alu/_0046_ ),
    .C(\alu/_0835_ ),
    .X(\alu/_0485_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2698_  (.A(net192),
    .B(\wAluB[31] ),
    .Y(\alu/_0486_ ));
 sky130_fd_sc_hd__o221a_1 \alu/_2699_  (.A1(\alu/_0486_ ),
    .A2(\alu/_0739_ ),
    .B1(\alu/_0582_ ),
    .B2(\alu/_0892_ ),
    .C1(\alu/_1196_ ),
    .X(\alu/_0487_ ));
 sky130_fd_sc_hd__o211a_1 \alu/_2700_  (.A1(\alu/_0484_ ),
    .A2(\alu/_0244_ ),
    .B1(\alu/_0485_ ),
    .C1(\alu/_0487_ ),
    .X(\alu/_0488_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2701_  (.A(\alu/_0044_ ),
    .B(\alu/_0292_ ),
    .Y(\alu/_0489_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2702_  (.A(\alu/_0483_ ),
    .B(\alu/_0488_ ),
    .C(\alu/_0489_ ),
    .Y(\alu/_0490_ ));
 sky130_fd_sc_hd__inv_2 \alu/_2703_  (.A(\alu/_0490_ ),
    .Y(\alu/_0491_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2704_  (.A(\alu/_0470_ ),
    .B(\alu/_0453_ ),
    .Y(\alu/_0492_ ));
 sky130_fd_sc_hd__nand2_1 \alu/_2705_  (.A(\alu/_0492_ ),
    .B(\alu/_0583_ ),
    .Y(\alu/_0494_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2706_  (.A(\alu/_0470_ ),
    .B(\alu/_0582_ ),
    .C(\alu/_0453_ ),
    .Y(\alu/_0495_ ));
 sky130_fd_sc_hd__nand3_1 \alu/_2707_  (.A(\alu/_0494_ ),
    .B(\alu/_1177_ ),
    .C(\alu/_0495_ ),
    .Y(\alu/_0496_ ));
 sky130_fd_sc_hd__nand3_4 \alu/_2708_  (.A(\alu/_0477_ ),
    .B(\alu/_0491_ ),
    .C(\alu/_0496_ ),
    .Y(\wAluOut[31] ));
 sky130_fd_sc_hd__nand2_1 \alu/_2709_  (.A(\alu/_0583_ ),
    .B(wAluSextEn),
    .Y(\alu/_0497_ ));
 sky130_fd_sc_hd__o21ai_1 \alu/_2710_  (.A1(\alu/_0497_ ),
    .A2(\alu/_0801_ ),
    .B1(\alu/_1114_ ),
    .Y(\alu/_0498_ ));
 sky130_fd_sc_hd__a21o_1 \alu/_2711_  (.A1(\alu/_0801_ ),
    .A2(\alu/_0497_ ),
    .B1(\alu/_0498_ ),
    .X(\alu/_0499_ ));
 sky130_fd_sc_hd__or2_1 \alu/_2712_  (.A(\alu/_0484_ ),
    .B(\alu/_1074_ ),
    .X(\alu/_0500_ ));
 sky130_fd_sc_hd__a31o_1 \alu/_2713_  (.A1(\alu/_0470_ ),
    .A2(\alu/_0486_ ),
    .A3(\alu/_0453_ ),
    .B1(\alu/_0500_ ),
    .X(\alu/_0501_ ));
 sky130_fd_sc_hd__nand2_2 \alu/_2714_  (.A(\alu/_0499_ ),
    .B(\alu/_0501_ ),
    .Y(wAluFlag));
 sky130_fd_sc_hd__o21a_1 \brancher/_1010_  (.A1(net902),
    .A2(net323),
    .B1(\brancher/rPc_current_reg1[0] ),
    .X(\wPcReturn[0] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1011_  (.A1(net902),
    .A2(net323),
    .B1(\brancher/rPc_current_reg1[1] ),
    .X(\wPcReturn[1] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1012_  (.A1(net900),
    .A2(net321),
    .B1(\brancher/rPc_current_reg1[2] ),
    .X(\wPcReturn[2] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1013_  (.A1(net904),
    .A2(net326),
    .B1(\brancher/rPc_current_reg1[3] ),
    .X(\wPcReturn[3] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1014_  (.A1(net906),
    .A2(net321),
    .B1(\brancher/rPc_current_reg1[4] ),
    .X(\wPcReturn[4] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1015_  (.A1(net900),
    .A2(net322),
    .B1(\brancher/rPc_current_reg1[5] ),
    .X(\wPcReturn[5] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1016_  (.A1(net901),
    .A2(net321),
    .B1(\brancher/rPc_current_reg1[6] ),
    .X(\wPcReturn[6] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1017_  (.A1(net904),
    .A2(net326),
    .B1(\brancher/rPc_current_reg1[7] ),
    .X(\wPcReturn[7] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1018_  (.A1(net900),
    .A2(net322),
    .B1(\brancher/rPc_current_reg1[8] ),
    .X(\wPcReturn[8] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1019_  (.A1(net900),
    .A2(net322),
    .B1(\brancher/rPc_current_reg1[9] ),
    .X(\wPcReturn[9] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1020_  (.A1(net901),
    .A2(net321),
    .B1(\brancher/rPc_current_reg1[10] ),
    .X(\wPcReturn[10] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1021_  (.A1(net901),
    .A2(net321),
    .B1(\brancher/rPc_current_reg1[11] ),
    .X(\wPcReturn[11] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1022_  (.A1(net898),
    .A2(net320),
    .B1(\brancher/rPc_current_reg1[12] ),
    .X(\wPcReturn[12] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1023_  (.A1(net900),
    .A2(net322),
    .B1(\brancher/rPc_current_reg1[13] ),
    .X(\wPcReturn[13] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1024_  (.A1(net900),
    .A2(net322),
    .B1(\brancher/rPc_current_reg1[14] ),
    .X(\wPcReturn[14] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1025_  (.A1(net898),
    .A2(net320),
    .B1(\brancher/rPc_current_reg1[15] ),
    .X(\wPcReturn[15] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1026_  (.A1(net898),
    .A2(net320),
    .B1(\brancher/rPc_current_reg1[16] ),
    .X(\wPcReturn[16] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1027_  (.A1(net898),
    .A2(net320),
    .B1(\brancher/rPc_current_reg1[17] ),
    .X(\wPcReturn[17] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1028_  (.A1(net898),
    .A2(net320),
    .B1(\brancher/rPc_current_reg1[18] ),
    .X(\wPcReturn[18] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1029_  (.A1(net899),
    .A2(net328),
    .B1(\brancher/rPc_current_reg1[19] ),
    .X(\wPcReturn[19] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1030_  (.A1(net899),
    .A2(net328),
    .B1(\brancher/rPc_current_reg1[20] ),
    .X(\wPcReturn[20] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1031_  (.A1(net905),
    .A2(net326),
    .B1(\brancher/rPc_current_reg1[21] ),
    .X(\wPcReturn[21] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1032_  (.A1(net904),
    .A2(net326),
    .B1(\brancher/rPc_current_reg1[22] ),
    .X(\wPcReturn[22] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1033_  (.A1(net903),
    .A2(net325),
    .B1(\brancher/rPc_current_reg1[23] ),
    .X(\wPcReturn[23] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1034_  (.A1(net903),
    .A2(net325),
    .B1(\brancher/rPc_current_reg1[24] ),
    .X(\wPcReturn[24] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1035_  (.A1(net903),
    .A2(net323),
    .B1(\brancher/rPc_current_reg1[25] ),
    .X(\wPcReturn[25] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1036_  (.A1(net903),
    .A2(net324),
    .B1(\brancher/rPc_current_reg1[26] ),
    .X(\wPcReturn[26] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1037_  (.A1(net902),
    .A2(net323),
    .B1(\brancher/rPc_current_reg1[27] ),
    .X(\wPcReturn[27] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1038_  (.A1(net905),
    .A2(net327),
    .B1(\brancher/rPc_current_reg1[28] ),
    .X(\wPcReturn[28] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1039_  (.A1(net902),
    .A2(net323),
    .B1(\brancher/rPc_current_reg1[29] ),
    .X(\wPcReturn[29] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1040_  (.A1(net902),
    .A2(net323),
    .B1(\brancher/rPc_current_reg1[30] ),
    .X(\wPcReturn[30] ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1041_  (.A1(net902),
    .A2(net324),
    .B1(\brancher/rPc_current_reg1[31] ),
    .X(\wPcReturn[31] ));
 sky130_fd_sc_hd__nand2_2 \brancher/_1042_  (.A(rCond),
    .B(\brancher/rOp_b_type ),
    .Y(\brancher/_0426_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1043_  (.A(\brancher/_0426_ ),
    .Y(\brancher/_0427_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1044_  (.A(\brancher/_0427_ ),
    .X(\brancher/_0428_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1045_  (.A(\brancher/_0428_ ),
    .X(\brancher/_0429_ ));
 sky130_fd_sc_hd__buf_2 \brancher/_1046_  (.A(\brancher/_0429_ ),
    .X(\brancher/_0430_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1047_  (.A(\brancher/_0426_ ),
    .X(\brancher/_0431_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1048_  (.A(\brancher/_0431_ ),
    .X(\brancher/_0432_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1049_  (.A(net943),
    .Y(\brancher/_0433_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1050_  (.A(\brancher/_0433_ ),
    .X(\brancher/_0434_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1051_  (.A1(\brancher/_0432_ ),
    .A2(\brancher/_0434_ ),
    .B1(\brancher/rPc_current_reg3[0] ),
    .X(\brancher/_0435_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1052_  (.A(net947),
    .Y(\brancher/_0436_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1053_  (.A(net944),
    .B(\brancher/_0436_ ),
    .Y(\brancher/_0437_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1054_  (.A(\brancher/_0437_ ),
    .Y(\brancher/_0438_ ));
 sky130_fd_sc_hd__o311ai_2 \brancher/_1055_  (.A1(net135),
    .A2(net944),
    .A3(\brancher/_0430_ ),
    .B1(\brancher/_0435_ ),
    .C1(\brancher/_0438_ ),
    .Y(\brancher/_0439_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1056_  (.A(\brancher/_0439_ ),
    .Y(\wPcNextCond[0] ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \brancher/_1057_  (.A(\brancher/_0436_ ),
    .X(\brancher/_0440_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1058_  (.A(\brancher/rAdder_b[1] ),
    .B(\brancher/rPc_current_reg3[1] ),
    .X(\brancher/_0441_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1059_  (.A(\brancher/rAdder_b[1] ),
    .B(\brancher/rPc_current_reg3[1] ),
    .Y(\brancher/_0442_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1060_  (.A1(\brancher/_0441_ ),
    .A2(\brancher/_0442_ ),
    .B1(\brancher/_0431_ ),
    .X(\brancher/_0443_ ));
 sky130_fd_sc_hd__o211a_1 \brancher/_1061_  (.A1(net146),
    .A2(\brancher/_0428_ ),
    .B1(\brancher/_0440_ ),
    .C1(\brancher/_0443_ ),
    .X(\brancher/_0444_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \brancher/_1062_  (.A(\brancher/_0433_ ),
    .X(\brancher/_0445_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1063_  (.A(\brancher/rPc_current_reg3[1] ),
    .B(\brancher/rAdder_jal[1] ),
    .X(\brancher/_0446_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1064_  (.A(\brancher/rPc_current_reg3[1] ),
    .B(\brancher/rAdder_jal[1] ),
    .Y(\brancher/_0447_ ));
 sky130_fd_sc_hd__and3_1 \brancher/_1065_  (.A(\brancher/_0446_ ),
    .B(net944),
    .C(\brancher/_0447_ ),
    .X(\brancher/_0448_ ));
 sky130_fd_sc_hd__a221o_1 \brancher/_1066_  (.A1(\brancher/rAlu_result[1] ),
    .A2(\brancher/_0437_ ),
    .B1(\brancher/_0444_ ),
    .B2(\brancher/_0445_ ),
    .C1(\brancher/_0448_ ),
    .X(\wPcNextCond[1] ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1067_  (.A(\brancher/rAdder_b[2] ),
    .B(\brancher/rPc_current_reg3[2] ),
    .Y(\brancher/_0449_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1068_  (.A(\brancher/rAdder_b[2] ),
    .B(\brancher/rPc_current_reg3[2] ),
    .Y(\brancher/_0450_ ));
 sky130_fd_sc_hd__or2b_1 \brancher/_1069_  (.A(\brancher/_0449_ ),
    .B_N(\brancher/_0450_ ),
    .X(\brancher/_0451_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1070_  (.A(\brancher/_0442_ ),
    .B(\brancher/_0451_ ),
    .X(\brancher/_0452_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1071_  (.A(\brancher/_0451_ ),
    .B(\brancher/_0442_ ),
    .Y(\brancher/_0453_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1072_  (.A(net378),
    .B(\brancher/_0429_ ),
    .Y(\brancher/_0454_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1073_  (.A1(\brancher/_0452_ ),
    .A2(\brancher/_0429_ ),
    .A3(\brancher/_0453_ ),
    .B1(\brancher/_0454_ ),
    .X(\brancher/_0455_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1074_  (.A(\brancher/_0440_ ),
    .X(\brancher/_0456_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1075_  (.A(\brancher/_0456_ ),
    .X(\brancher/_0457_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1076_  (.A(\brancher/_0433_ ),
    .X(\brancher/_0458_ ));
 sky130_fd_sc_hd__buf_2 \brancher/_1077_  (.A(\brancher/_0458_ ),
    .X(\brancher/_0459_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1078_  (.A(\brancher/_0447_ ),
    .Y(\brancher/_0460_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1079_  (.A(\brancher/rPc_current_reg3[2] ),
    .B(\brancher/rAdder_jal[2] ),
    .Y(\brancher/_0461_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1080_  (.A(\brancher/rPc_current_reg3[2] ),
    .B(\brancher/rAdder_jal[2] ),
    .Y(\brancher/_0462_ ));
 sky130_fd_sc_hd__nor2b_1 \brancher/_1081_  (.A(\brancher/_0461_ ),
    .B_N(\brancher/_0462_ ),
    .Y(\brancher/_0463_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1082_  (.A(\brancher/_0460_ ),
    .B(\brancher/_0463_ ),
    .X(\brancher/_0464_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1083_  (.A(\brancher/_0463_ ),
    .B(\brancher/_0460_ ),
    .Y(\brancher/_0465_ ));
 sky130_fd_sc_hd__a32o_1 \brancher/_1084_  (.A1(\brancher/_0464_ ),
    .A2(net942),
    .A3(\brancher/_0465_ ),
    .B1(\brancher/rAlu_result[2] ),
    .B2(\brancher/_0437_ ),
    .X(\brancher/_0466_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1085_  (.A1(\brancher/_0455_ ),
    .A2(\brancher/_0457_ ),
    .A3(\brancher/_0459_ ),
    .B1(\brancher/_0466_ ),
    .X(\wPcNextCond[2] ));
 sky130_fd_sc_hd__inv_2 \brancher/_1086_  (.A(\brancher/rAdder_b[3] ),
    .Y(\brancher/_0467_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1087_  (.A(\brancher/rPc_current_reg3[3] ),
    .Y(\brancher/_0468_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1088_  (.A(\brancher/_0467_ ),
    .B(\brancher/_0468_ ),
    .Y(\brancher/_0469_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1089_  (.A(\brancher/rAdder_b[3] ),
    .B(\brancher/rPc_current_reg3[3] ),
    .Y(\brancher/_0470_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1090_  (.A(\brancher/_0469_ ),
    .B(\brancher/_0470_ ),
    .Y(\brancher/_0471_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1091_  (.A(\brancher/_0471_ ),
    .Y(\brancher/_0472_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1092_  (.A1(\brancher/_0442_ ),
    .A2(\brancher/_0449_ ),
    .B1(\brancher/_0450_ ),
    .Y(\brancher/_0473_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1093_  (.A(\brancher/_0472_ ),
    .B(\brancher/_0473_ ),
    .X(\brancher/_0474_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1094_  (.A(\brancher/_0473_ ),
    .B(\brancher/_0472_ ),
    .Y(\brancher/_0475_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1095_  (.A(net378),
    .B(net377),
    .X(\brancher/_0476_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1096_  (.A(net378),
    .B(net377),
    .Y(\brancher/_0477_ ));
 sky130_fd_sc_hd__and3_1 \brancher/_1097_  (.A(\brancher/_0476_ ),
    .B(\brancher/_0426_ ),
    .C(\brancher/_0477_ ),
    .X(\brancher/_0478_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1098_  (.A1(\brancher/_0474_ ),
    .A2(\brancher/_0428_ ),
    .A3(\brancher/_0475_ ),
    .B1(\brancher/_0478_ ),
    .X(\brancher/_0479_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1099_  (.A(net947),
    .B(net944),
    .Y(\brancher/_0480_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1100_  (.A(\brancher/rPc_current_reg3[3] ),
    .B(\brancher/rAdder_jal[3] ),
    .Y(\brancher/_0481_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1101_  (.A(\brancher/rPc_current_reg3[3] ),
    .B(\brancher/rAdder_jal[3] ),
    .Y(\brancher/_0482_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1102_  (.A(\brancher/_0482_ ),
    .Y(\brancher/_0483_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1103_  (.A(\brancher/_0481_ ),
    .B(\brancher/_0483_ ),
    .Y(\brancher/_0484_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1104_  (.A(\brancher/_0465_ ),
    .B(\brancher/_0462_ ),
    .Y(\brancher/_0485_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1105_  (.A(\brancher/_0484_ ),
    .B(\brancher/_0485_ ),
    .X(\brancher/_0486_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1106_  (.A(\brancher/_0485_ ),
    .B(\brancher/_0484_ ),
    .Y(\brancher/_0487_ ));
 sky130_fd_sc_hd__and3_1 \brancher/_1107_  (.A(\brancher/_0486_ ),
    .B(net942),
    .C(\brancher/_0487_ ),
    .X(\brancher/_0488_ ));
 sky130_fd_sc_hd__a221o_1 \brancher/_1108_  (.A1(\brancher/rAlu_result[3] ),
    .A2(\brancher/_0437_ ),
    .B1(\brancher/_0479_ ),
    .B2(\brancher/_0480_ ),
    .C1(\brancher/_0488_ ),
    .X(\wPcNextCond[3] ));
 sky130_fd_sc_hd__and2_1 \brancher/_1109_  (.A(\brancher/_0487_ ),
    .B(\brancher/_0482_ ),
    .X(\brancher/_0489_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1110_  (.A(\brancher/rPc_current_reg3[4] ),
    .B(\brancher/rAdder_jal[4] ),
    .X(\brancher/_0490_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1111_  (.A(\brancher/rPc_current_reg3[4] ),
    .B(\brancher/rAdder_jal[4] ),
    .Y(\brancher/_0491_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1112_  (.A(\brancher/_0490_ ),
    .B(\brancher/_0491_ ),
    .Y(\brancher/_0492_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1113_  (.A(\brancher/_0489_ ),
    .B(\brancher/_0492_ ),
    .Y(\brancher/_0493_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1114_  (.A(\brancher/_0492_ ),
    .B(\brancher/_0489_ ),
    .X(\brancher/_0494_ ));
 sky130_fd_sc_hd__and2_1 \brancher/_1115_  (.A(\brancher/_0475_ ),
    .B(\brancher/_0470_ ),
    .X(\brancher/_0495_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1116_  (.A(\brancher/rAdder_b[4] ),
    .Y(\brancher/_0496_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1117_  (.A(\brancher/rPc_current_reg3[4] ),
    .Y(\brancher/_0497_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1118_  (.A(\brancher/_0496_ ),
    .B(\brancher/_0497_ ),
    .Y(\brancher/_0498_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1119_  (.A(\brancher/rAdder_b[4] ),
    .B(\brancher/rPc_current_reg3[4] ),
    .Y(\brancher/_0499_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1120_  (.A(\brancher/_0498_ ),
    .B(\brancher/_0499_ ),
    .Y(\brancher/_0500_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1121_  (.A(\brancher/_0500_ ),
    .B(\brancher/_0495_ ),
    .Y(\brancher/_0501_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1122_  (.A(\brancher/_0426_ ),
    .B(\brancher/_0501_ ),
    .X(\brancher/_0502_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1123_  (.A1(\brancher/_0495_ ),
    .A2(\brancher/_0500_ ),
    .B1(\brancher/_0502_ ),
    .X(\brancher/_0503_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1124_  (.A(\brancher/_0436_ ),
    .X(\brancher/_0504_ ));
 sky130_fd_sc_hd__inv_4 \brancher/_1125_  (.A(\brancher/_0477_ ),
    .Y(\brancher/_0505_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1126_  (.A(net376),
    .B(\brancher/_0505_ ),
    .Y(\brancher/_0506_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1127_  (.A(\brancher/_0505_ ),
    .B(net376),
    .Y(\brancher/_0507_ ));
 sky130_fd_sc_hd__or3b_1 \brancher/_1128_  (.A(\brancher/_0427_ ),
    .B(\brancher/_0506_ ),
    .C_N(\brancher/_0507_ ),
    .X(\brancher/_0508_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1129_  (.A(\brancher/_0503_ ),
    .B(\brancher/_0504_ ),
    .C(\brancher/_0508_ ),
    .Y(\brancher/_0509_ ));
 sky130_fd_sc_hd__o211a_1 \brancher/_1130_  (.A1(\brancher/_0456_ ),
    .A2(\brancher/rAlu_result[4] ),
    .B1(\brancher/_0434_ ),
    .C1(\brancher/_0509_ ),
    .X(\brancher/_0510_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1131_  (.A1(net942),
    .A2(\brancher/_0493_ ),
    .A3(\brancher/_0494_ ),
    .B1(\brancher/_0510_ ),
    .X(\wPcNextCond[4] ));
 sky130_fd_sc_hd__nor2b_1 \brancher/_1132_  (.A(\brancher/_0492_ ),
    .B_N(\brancher/_0484_ ),
    .Y(\brancher/_0511_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1133_  (.A(\brancher/_0485_ ),
    .B(\brancher/_0511_ ),
    .Y(\brancher/_0512_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1134_  (.A1(\brancher/_0482_ ),
    .A2(\brancher/_0492_ ),
    .B1(\brancher/_0491_ ),
    .X(\brancher/_0513_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1135_  (.A(\brancher/_0512_ ),
    .B(\brancher/_0513_ ),
    .Y(\brancher/_0514_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1136_  (.A(\brancher/rPc_current_reg3[5] ),
    .B(\brancher/rAdder_jal[5] ),
    .Y(\brancher/_0515_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1137_  (.A(\brancher/rPc_current_reg3[5] ),
    .B(\brancher/rAdder_jal[5] ),
    .Y(\brancher/_0516_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1138_  (.A(\brancher/_0516_ ),
    .Y(\brancher/_0517_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1139_  (.A(\brancher/_0515_ ),
    .B(\brancher/_0517_ ),
    .Y(\brancher/_0518_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1140_  (.A(\brancher/_0514_ ),
    .B(\brancher/_0518_ ),
    .Y(\brancher/_0519_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1141_  (.A(\brancher/_0518_ ),
    .B(\brancher/_0514_ ),
    .X(\brancher/_0520_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1142_  (.A(net375),
    .Y(\brancher/_0521_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1143_  (.A(\brancher/_0521_ ),
    .B(\brancher/_0507_ ),
    .Y(\brancher/_0522_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1144_  (.A(\brancher/_0507_ ),
    .B(\brancher/_0521_ ),
    .Y(\brancher/_0523_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1145_  (.A(\brancher/_0523_ ),
    .B(\brancher/_0431_ ),
    .Y(\brancher/_0524_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1146_  (.A1(\brancher/_0522_ ),
    .A2(\brancher/_0524_ ),
    .B1(\brancher/_0440_ ),
    .Y(\brancher/_0525_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1147_  (.A(\brancher/rAdder_b[5] ),
    .B(\brancher/rPc_current_reg3[5] ),
    .Y(\brancher/_0526_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1148_  (.A(\brancher/rAdder_b[5] ),
    .B(\brancher/rPc_current_reg3[5] ),
    .Y(\brancher/_0527_ ));
 sky130_fd_sc_hd__and2b_1 \brancher/_1149_  (.A_N(\brancher/_0526_ ),
    .B(\brancher/_0527_ ),
    .X(\brancher/_0528_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1150_  (.A(\brancher/_0471_ ),
    .B(\brancher/_0500_ ),
    .Y(\brancher/_0529_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1151_  (.A(\brancher/_0529_ ),
    .B(\brancher/_0473_ ),
    .Y(\brancher/_0530_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1152_  (.A(\brancher/rAdder_b[4] ),
    .B(\brancher/rPc_current_reg3[4] ),
    .Y(\brancher/_0531_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1153_  (.A1(\brancher/_0470_ ),
    .A2(\brancher/_0531_ ),
    .B1(\brancher/_0499_ ),
    .X(\brancher/_0532_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1154_  (.A(\brancher/_0530_ ),
    .B(\brancher/_0532_ ),
    .Y(\brancher/_0533_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1155_  (.A(\brancher/_0528_ ),
    .B(\brancher/_0533_ ),
    .X(\brancher/_0534_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \brancher/_1156_  (.A(\brancher/_0427_ ),
    .X(\brancher/_0535_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1157_  (.A(\brancher/_0533_ ),
    .B(\brancher/_0528_ ),
    .Y(\brancher/_0536_ ));
 sky130_fd_sc_hd__and3_1 \brancher/_1158_  (.A(\brancher/_0534_ ),
    .B(\brancher/_0535_ ),
    .C(\brancher/_0536_ ),
    .X(\brancher/_0537_ ));
 sky130_fd_sc_hd__o221a_1 \brancher/_1159_  (.A1(\brancher/_0456_ ),
    .A2(\brancher/rAlu_result[5] ),
    .B1(\brancher/_0525_ ),
    .B2(\brancher/_0537_ ),
    .C1(\brancher/_0434_ ),
    .X(\brancher/_0538_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1160_  (.A1(net942),
    .A2(\brancher/_0519_ ),
    .A3(\brancher/_0520_ ),
    .B1(\brancher/_0538_ ),
    .X(\wPcNextCond[5] ));
 sky130_fd_sc_hd__or2_1 \brancher/_1161_  (.A(\brancher/rPc_current_reg3[6] ),
    .B(\brancher/rAdder_jal[6] ),
    .X(\brancher/_0539_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1162_  (.A(\brancher/rPc_current_reg3[6] ),
    .B(\brancher/rAdder_jal[6] ),
    .Y(\brancher/_0540_ ));
 sky130_fd_sc_hd__and2_1 \brancher/_1163_  (.A(\brancher/_0539_ ),
    .B(\brancher/_0540_ ),
    .X(\brancher/_0541_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1164_  (.A(\brancher/_0519_ ),
    .B(\brancher/_0516_ ),
    .Y(\brancher/_0542_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1165_  (.A(\brancher/_0541_ ),
    .B(\brancher/_0542_ ),
    .X(\brancher/_0543_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1166_  (.A(\brancher/_0542_ ),
    .B(\brancher/_0541_ ),
    .Y(\brancher/_0544_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1167_  (.A(\brancher/_0536_ ),
    .B(\brancher/_0527_ ),
    .Y(\brancher/_0545_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1168_  (.A(\brancher/rAdder_b[6] ),
    .B(\brancher/rPc_current_reg3[6] ),
    .Y(\brancher/_0546_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1169_  (.A(\brancher/rAdder_b[6] ),
    .B(\brancher/rPc_current_reg3[6] ),
    .Y(\brancher/_0547_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1170_  (.A(\brancher/_0547_ ),
    .Y(\brancher/_0548_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1171_  (.A(\brancher/_0546_ ),
    .B(\brancher/_0548_ ),
    .Y(\brancher/_0549_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1172_  (.A(\brancher/_0549_ ),
    .B(\brancher/_0545_ ),
    .X(\brancher/_0550_ ));
 sky130_fd_sc_hd__buf_2 \brancher/_1173_  (.A(\brancher/_0535_ ),
    .X(\brancher/_0551_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1174_  (.A(\brancher/_0550_ ),
    .B(\brancher/_0551_ ),
    .Y(\brancher/_0552_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1175_  (.A1(\brancher/_0545_ ),
    .A2(\brancher/_0549_ ),
    .B1(\brancher/_0552_ ),
    .X(\brancher/_0553_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1176_  (.A(net373),
    .B(\brancher/_0522_ ),
    .Y(\brancher/_0554_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1177_  (.A(\brancher/_0522_ ),
    .B(net373),
    .Y(\brancher/_0555_ ));
 sky130_fd_sc_hd__or3b_1 \brancher/_1178_  (.A(\brancher/_0535_ ),
    .B(\brancher/_0554_ ),
    .C_N(\brancher/_0555_ ),
    .X(\brancher/_0556_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1179_  (.A(\brancher/_0553_ ),
    .B(\brancher/_0457_ ),
    .C(\brancher/_0556_ ),
    .Y(\brancher/_0557_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1180_  (.A1(\brancher/rAlu_result[6] ),
    .A2(\brancher/_0456_ ),
    .B1(\brancher/_0458_ ),
    .X(\brancher/_0558_ ));
 sky130_fd_sc_hd__a32o_1 \brancher/_1181_  (.A1(net942),
    .A2(\brancher/_0543_ ),
    .A3(\brancher/_0544_ ),
    .B1(\brancher/_0557_ ),
    .B2(\brancher/_0558_ ),
    .X(\wPcNextCond[6] ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1182_  (.A(\brancher/rPc_current_reg3[7] ),
    .B(\brancher/rAdder_jal[7] ),
    .Y(\brancher/_0559_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1183_  (.A(\brancher/rPc_current_reg3[7] ),
    .B(\brancher/rAdder_jal[7] ),
    .Y(\brancher/_0560_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1184_  (.A(\brancher/_0560_ ),
    .Y(\brancher/_0561_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1185_  (.A(\brancher/_0559_ ),
    .B(\brancher/_0561_ ),
    .Y(\brancher/_0562_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1186_  (.A(\brancher/_0562_ ),
    .Y(\brancher/_0563_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1187_  (.A(\brancher/_0541_ ),
    .B(\brancher/_0518_ ),
    .Y(\brancher/_0564_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1188_  (.A(\brancher/_0514_ ),
    .Y(\brancher/_0565_ ));
 sky130_fd_sc_hd__a21bo_1 \brancher/_1189_  (.A1(\brancher/_0539_ ),
    .A2(\brancher/_0517_ ),
    .B1_N(\brancher/_0540_ ),
    .X(\brancher/_0566_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1190_  (.A(\brancher/_0566_ ),
    .Y(\brancher/_0567_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1191_  (.A1(\brancher/_0564_ ),
    .A2(\brancher/_0565_ ),
    .B1(\brancher/_0567_ ),
    .X(\brancher/_0568_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1192_  (.A(\brancher/_0563_ ),
    .B(\brancher/_0568_ ),
    .Y(\brancher/_0569_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1193_  (.A1(\brancher/_0568_ ),
    .A2(\brancher/_0563_ ),
    .B1(\brancher/_0458_ ),
    .X(\brancher/_0570_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1194_  (.A(\brancher/rAdder_b[7] ),
    .Y(\brancher/_0571_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1195_  (.A(\brancher/rPc_current_reg3[7] ),
    .Y(\brancher/_0572_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1196_  (.A(\brancher/_0571_ ),
    .B(\brancher/_0572_ ),
    .Y(\brancher/_0573_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1197_  (.A(\brancher/rAdder_b[7] ),
    .B(\brancher/rPc_current_reg3[7] ),
    .Y(\brancher/_0574_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1198_  (.A(\brancher/_0573_ ),
    .B(\brancher/_0574_ ),
    .Y(\brancher/_0575_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1199_  (.A(\brancher/_0575_ ),
    .Y(\brancher/_0576_ ));
 sky130_fd_sc_hd__and2_1 \brancher/_1200_  (.A(\brancher/_0528_ ),
    .B(\brancher/_0549_ ),
    .X(\brancher/_0577_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1201_  (.A1(\brancher/_0527_ ),
    .A2(\brancher/_0547_ ),
    .B1(\brancher/_0546_ ),
    .Y(\brancher/_0578_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1202_  (.A1(\brancher/_0533_ ),
    .A2(\brancher/_0577_ ),
    .B1(\brancher/_0578_ ),
    .X(\brancher/_0579_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1203_  (.A(\brancher/_0576_ ),
    .B(\brancher/_0579_ ),
    .X(\brancher/_0580_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1204_  (.A(\brancher/_0579_ ),
    .B(\brancher/_0576_ ),
    .Y(\brancher/_0581_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1205_  (.A(net372),
    .Y(\brancher/_0582_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1206_  (.A(\brancher/_0582_ ),
    .B(\brancher/_0555_ ),
    .Y(\brancher/_0583_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1207_  (.A(\brancher/_0427_ ),
    .B(\brancher/_0583_ ),
    .X(\brancher/_0584_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1208_  (.A1(\brancher/_0582_ ),
    .A2(\brancher/_0555_ ),
    .B1(\brancher/_0584_ ),
    .Y(\brancher/_0585_ ));
 sky130_fd_sc_hd__a311o_1 \brancher/_1209_  (.A1(\brancher/_0580_ ),
    .A2(\brancher/_0581_ ),
    .A3(\brancher/_0551_ ),
    .B1(net947),
    .C1(\brancher/_0585_ ),
    .X(\brancher/_0586_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1210_  (.A(\brancher/_0440_ ),
    .X(\brancher/_0587_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1211_  (.A(\brancher/_0433_ ),
    .X(\brancher/_0588_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1212_  (.A1(\brancher/rAlu_result[7] ),
    .A2(\brancher/_0587_ ),
    .B1(\brancher/_0588_ ),
    .X(\brancher/_0589_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1213_  (.A(\brancher/_0586_ ),
    .B(\brancher/_0589_ ),
    .Y(\brancher/_0590_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1214_  (.A1(\brancher/_0569_ ),
    .A2(\brancher/_0570_ ),
    .B1(\brancher/_0590_ ),
    .Y(\wPcNextCond[7] ));
 sky130_fd_sc_hd__or2_1 \brancher/_1215_  (.A(\brancher/rPc_current_reg3[8] ),
    .B(\brancher/rAdder_jal[8] ),
    .X(\brancher/_0591_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1216_  (.A(\brancher/rPc_current_reg3[8] ),
    .B(\brancher/rAdder_jal[8] ),
    .Y(\brancher/_0592_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1217_  (.A(\brancher/_0591_ ),
    .B(\brancher/_0592_ ),
    .Y(\brancher/_0593_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1218_  (.A(\brancher/_0561_ ),
    .B(\brancher/_0569_ ),
    .X(\brancher/_0594_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1219_  (.A(\brancher/_0593_ ),
    .B(\brancher/_0594_ ),
    .X(\brancher/_0595_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1220_  (.A(\brancher/_0594_ ),
    .B(\brancher/_0593_ ),
    .Y(\brancher/_0596_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1221_  (.A1(\brancher/_0595_ ),
    .A2(\brancher/_0596_ ),
    .B1(\brancher/_0459_ ),
    .X(\brancher/_0597_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1222_  (.A(\brancher/_0581_ ),
    .B(\brancher/_0574_ ),
    .Y(\brancher/_0598_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1223_  (.A(\brancher/rAdder_b[8] ),
    .Y(\brancher/_0599_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1224_  (.A(\brancher/rPc_current_reg3[8] ),
    .Y(\brancher/_0600_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1225_  (.A(\brancher/_0599_ ),
    .B(\brancher/_0600_ ),
    .Y(\brancher/_0601_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1226_  (.A(\brancher/rAdder_b[8] ),
    .B(\brancher/rPc_current_reg3[8] ),
    .Y(\brancher/_0602_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1227_  (.A(\brancher/_0601_ ),
    .B(\brancher/_0602_ ),
    .Y(\brancher/_0603_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1228_  (.A(\brancher/_0603_ ),
    .Y(\brancher/_0604_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1229_  (.A(\brancher/_0426_ ),
    .X(\brancher/_0605_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1230_  (.A1(\brancher/_0598_ ),
    .A2(\brancher/_0604_ ),
    .B1(\brancher/_0605_ ),
    .Y(\brancher/_0606_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1231_  (.A1(\brancher/_0598_ ),
    .A2(\brancher/_0604_ ),
    .B1(\brancher/_0606_ ),
    .Y(\brancher/_0607_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1232_  (.A(\brancher/_0440_ ),
    .X(\brancher/_0608_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1233_  (.A(net371),
    .B(\brancher/_0583_ ),
    .Y(\brancher/_0609_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1234_  (.A(\brancher/_0583_ ),
    .B(net371),
    .Y(\brancher/_0610_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1235_  (.A(\brancher/_0610_ ),
    .Y(\brancher/_0611_ ));
 sky130_fd_sc_hd__or3_1 \brancher/_1236_  (.A(\brancher/_0535_ ),
    .B(\brancher/_0609_ ),
    .C(\brancher/_0611_ ),
    .X(\brancher/_0612_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1237_  (.A1(\brancher/rAlu_result[8] ),
    .A2(\brancher/_0504_ ),
    .B1(\brancher/_0434_ ),
    .Y(\brancher/_0613_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1238_  (.A1(\brancher/_0607_ ),
    .A2(\brancher/_0608_ ),
    .A3(\brancher/_0612_ ),
    .B1(\brancher/_0613_ ),
    .X(\brancher/_0614_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1239_  (.A(\brancher/_0597_ ),
    .B(\brancher/_0614_ ),
    .Y(\wPcNextCond[8] ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1240_  (.A(\brancher/rPc_current_reg3[9] ),
    .B(\brancher/rAdder_jal[9] ),
    .Y(\brancher/_0615_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1241_  (.A(\brancher/rPc_current_reg3[9] ),
    .B(\brancher/rAdder_jal[9] ),
    .Y(\brancher/_0616_ ));
 sky130_fd_sc_hd__and2b_1 \brancher/_1242_  (.A_N(\brancher/_0615_ ),
    .B(\brancher/_0616_ ),
    .X(\brancher/_0617_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1243_  (.A(\brancher/_0593_ ),
    .B(\brancher/_0563_ ),
    .Y(\brancher/_0618_ ));
 sky130_fd_sc_hd__nor2b_1 \brancher/_1244_  (.A(\brancher/_0564_ ),
    .B_N(\brancher/_0618_ ),
    .Y(\brancher/_0619_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1245_  (.A(\brancher/_0514_ ),
    .B(\brancher/_0619_ ),
    .Y(\brancher/_0620_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1246_  (.A1(\brancher/_0560_ ),
    .A2(\brancher/_0593_ ),
    .B1(\brancher/_0592_ ),
    .Y(\brancher/_0621_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1247_  (.A1(\brancher/_0566_ ),
    .A2(\brancher/_0618_ ),
    .B1(\brancher/_0621_ ),
    .Y(\brancher/_0622_ ));
 sky130_fd_sc_hd__nand2_2 \brancher/_1248_  (.A(\brancher/_0620_ ),
    .B(\brancher/_0622_ ),
    .Y(\brancher/_0623_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1249_  (.A(\brancher/_0617_ ),
    .B(\brancher/_0623_ ),
    .X(\brancher/_0624_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1250_  (.A(\brancher/_0623_ ),
    .B(\brancher/_0617_ ),
    .Y(\brancher/_0625_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1251_  (.A(\brancher/_0576_ ),
    .B(\brancher/_0604_ ),
    .Y(\brancher/_0626_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1252_  (.A(\brancher/_0528_ ),
    .B(\brancher/_0549_ ),
    .Y(\brancher/_0627_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1253_  (.A(\brancher/_0626_ ),
    .B(\brancher/_0627_ ),
    .Y(\brancher/_0628_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1254_  (.A(\brancher/_0533_ ),
    .B(\brancher/_0628_ ),
    .Y(\brancher/_0629_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1255_  (.A(\brancher/_0575_ ),
    .B(\brancher/_0603_ ),
    .Y(\brancher/_0630_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1256_  (.A(\brancher/_0601_ ),
    .Y(\brancher/_0631_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1257_  (.A1(\brancher/_0574_ ),
    .A2(\brancher/_0631_ ),
    .B1(\brancher/_0602_ ),
    .Y(\brancher/_0632_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1258_  (.A1(\brancher/_0630_ ),
    .A2(\brancher/_0578_ ),
    .B1(\brancher/_0632_ ),
    .Y(\brancher/_0633_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1259_  (.A(\brancher/rAdder_b[9] ),
    .B(\brancher/rPc_current_reg3[9] ),
    .X(\brancher/_0634_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1260_  (.A(\brancher/rAdder_b[9] ),
    .B(\brancher/rPc_current_reg3[9] ),
    .Y(\brancher/_0635_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1261_  (.A(\brancher/_0634_ ),
    .B(\brancher/_0635_ ),
    .Y(\brancher/_0636_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1262_  (.A(\brancher/_0629_ ),
    .B(\brancher/_0633_ ),
    .Y(\brancher/_0637_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1263_  (.A(\brancher/_0637_ ),
    .B(\brancher/_0634_ ),
    .C(\brancher/_0635_ ),
    .Y(\brancher/_0638_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1264_  (.A(\brancher/_0638_ ),
    .B(\brancher/_0428_ ),
    .Y(\brancher/_0639_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1265_  (.A1(\brancher/_0629_ ),
    .A2(\brancher/_0633_ ),
    .A3(\brancher/_0636_ ),
    .B1(\brancher/_0639_ ),
    .X(\brancher/_0640_ ));
 sky130_fd_sc_hd__and4_1 \brancher/_1266_  (.A(net373),
    .B(net372),
    .C(net371),
    .D(net370),
    .X(\brancher/_0641_ ));
 sky130_fd_sc_hd__and2_1 \brancher/_1267_  (.A(\brancher/_0641_ ),
    .B(\brancher/_0522_ ),
    .X(\brancher/_0642_ ));
 sky130_fd_sc_hd__buf_6 \brancher/_1268_  (.A(\brancher/_0642_ ),
    .X(\brancher/_0643_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1269_  (.A(\brancher/_0429_ ),
    .B(\brancher/_0643_ ),
    .Y(\brancher/_0644_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1270_  (.A1(net370),
    .A2(\brancher/_0611_ ),
    .B1(\brancher/_0644_ ),
    .Y(\brancher/_0645_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1271_  (.A(\brancher/_0640_ ),
    .B(\brancher/_0457_ ),
    .C(\brancher/_0645_ ),
    .Y(\brancher/_0646_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1272_  (.A1(\brancher/rAlu_result[9] ),
    .A2(\brancher/_0456_ ),
    .B1(\brancher/_0458_ ),
    .X(\brancher/_0647_ ));
 sky130_fd_sc_hd__a32o_1 \brancher/_1273_  (.A1(net942),
    .A2(\brancher/_0624_ ),
    .A3(\brancher/_0625_ ),
    .B1(\brancher/_0646_ ),
    .B2(\brancher/_0647_ ),
    .X(\wPcNextCond[9] ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1274_  (.A1(\brancher/rAlu_result[10] ),
    .A2(\brancher/_0457_ ),
    .B1(\brancher/_0459_ ),
    .Y(\brancher/_0648_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1275_  (.A(\brancher/rAdder_b[10] ),
    .B(\brancher/rPc_current_reg3[10] ),
    .Y(\brancher/_0649_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1276_  (.A(\brancher/rAdder_b[10] ),
    .B(\brancher/rPc_current_reg3[10] ),
    .Y(\brancher/_0650_ ));
 sky130_fd_sc_hd__nand2b_1 \brancher/_1277_  (.A_N(\brancher/_0649_ ),
    .B(\brancher/_0650_ ),
    .Y(\brancher/_0651_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1278_  (.A1(\brancher/_0638_ ),
    .A2(\brancher/_0635_ ),
    .B1(\brancher/_0651_ ),
    .Y(\brancher/_0652_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1279_  (.A1(\brancher/_0638_ ),
    .A2(\brancher/_0635_ ),
    .A3(\brancher/_0651_ ),
    .B1(\brancher/_0426_ ),
    .X(\brancher/_0653_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1280_  (.A(net368),
    .B(\brancher/_0643_ ),
    .Y(\brancher/_0654_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1281_  (.A(\brancher/_0643_ ),
    .B(net368),
    .Y(\brancher/_0655_ ));
 sky130_fd_sc_hd__or3b_1 \brancher/_1282_  (.A(\brancher/_0535_ ),
    .B(\brancher/_0654_ ),
    .C_N(\brancher/_0655_ ),
    .X(\brancher/_0656_ ));
 sky130_fd_sc_hd__o211a_1 \brancher/_1283_  (.A1(\brancher/_0652_ ),
    .A2(\brancher/_0653_ ),
    .B1(\brancher/_0504_ ),
    .C1(\brancher/_0656_ ),
    .X(\brancher/_0657_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1284_  (.A(\brancher/_0625_ ),
    .B(\brancher/_0616_ ),
    .Y(\brancher/_0658_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1285_  (.A(\brancher/rPc_current_reg3[10] ),
    .B(\brancher/rAdder_jal[10] ),
    .Y(\brancher/_0659_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1286_  (.A(\brancher/rPc_current_reg3[10] ),
    .B(\brancher/rAdder_jal[10] ),
    .X(\brancher/_0660_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1287_  (.A(\brancher/_0660_ ),
    .B(\brancher/_0659_ ),
    .Y(\brancher/_0661_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1288_  (.A1(\brancher/_0625_ ),
    .A2(\brancher/_0616_ ),
    .A3(\brancher/_0661_ ),
    .B1(\brancher/_0458_ ),
    .X(\brancher/_0662_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1289_  (.A1(\brancher/_0658_ ),
    .A2(\brancher/_0659_ ),
    .A3(\brancher/_0660_ ),
    .B1(\brancher/_0662_ ),
    .X(\brancher/_0663_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1290_  (.A1(\brancher/_0648_ ),
    .A2(\brancher/_0657_ ),
    .B1(\brancher/_0663_ ),
    .Y(\wPcNextCond[10] ));
 sky130_fd_sc_hd__or2_1 \brancher/_1291_  (.A(\brancher/rPc_current_reg3[11] ),
    .B(\brancher/rAdder_jal[11] ),
    .X(\brancher/_0664_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1292_  (.A(\brancher/rPc_current_reg3[11] ),
    .B(\brancher/rAdder_jal[11] ),
    .Y(\brancher/_0665_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1293_  (.A(\brancher/_0664_ ),
    .B(\brancher/_0665_ ),
    .Y(\brancher/_0666_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1294_  (.A(\brancher/_0666_ ),
    .Y(\brancher/_0667_ ));
 sky130_fd_sc_hd__and3_1 \brancher/_1295_  (.A(\brancher/_0617_ ),
    .B(\brancher/_0659_ ),
    .C(\brancher/_0660_ ),
    .X(\brancher/_0668_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1296_  (.A(\brancher/_0623_ ),
    .B(\brancher/_0668_ ),
    .Y(\brancher/_0669_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1297_  (.A(\brancher/_0616_ ),
    .B(\brancher/_0661_ ),
    .X(\brancher/_0670_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1298_  (.A(\brancher/_0669_ ),
    .B(\brancher/_0659_ ),
    .C(\brancher/_0670_ ),
    .Y(\brancher/_0671_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1299_  (.A(\brancher/_0667_ ),
    .B(\brancher/_0671_ ),
    .X(\brancher/_0672_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1300_  (.A(\brancher/_0671_ ),
    .B(\brancher/_0667_ ),
    .Y(\brancher/_0673_ ));
 sky130_fd_sc_hd__and2_1 \brancher/_1301_  (.A(\brancher/_0673_ ),
    .B(net943),
    .X(\brancher/_0674_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1302_  (.A(\brancher/_0636_ ),
    .B(\brancher/_0651_ ),
    .Y(\brancher/_0675_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1303_  (.A(\brancher/_0637_ ),
    .B(\brancher/_0675_ ),
    .Y(\brancher/_0676_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1304_  (.A1(\brancher/_0635_ ),
    .A2(\brancher/_0650_ ),
    .B1(\brancher/_0649_ ),
    .Y(\brancher/_0677_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1305_  (.A(\brancher/_0677_ ),
    .Y(\brancher/_0678_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1306_  (.A(\brancher/rAdder_b[11] ),
    .Y(\brancher/_0679_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1307_  (.A(\brancher/rPc_current_reg3[11] ),
    .Y(\brancher/_0680_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1308_  (.A(\brancher/_0679_ ),
    .B(\brancher/_0680_ ),
    .Y(\brancher/_0681_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1309_  (.A(\brancher/rAdder_b[11] ),
    .B(\brancher/rPc_current_reg3[11] ),
    .Y(\brancher/_0682_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1310_  (.A(\brancher/_0681_ ),
    .B(\brancher/_0682_ ),
    .Y(\brancher/_0683_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1311_  (.A(\brancher/_0676_ ),
    .B(\brancher/_0678_ ),
    .Y(\brancher/_0684_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1312_  (.A(\brancher/_0684_ ),
    .B(\brancher/_0681_ ),
    .C(\brancher/_0682_ ),
    .Y(\brancher/_0685_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1313_  (.A(\brancher/_0685_ ),
    .B(\brancher/_0551_ ),
    .Y(\brancher/_0686_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1314_  (.A1(\brancher/_0676_ ),
    .A2(\brancher/_0678_ ),
    .A3(\brancher/_0683_ ),
    .B1(\brancher/_0686_ ),
    .X(\brancher/_0687_ ));
 sky130_fd_sc_hd__clkinvlp_2 \brancher/_1315_  (.A(\brancher/_0643_ ),
    .Y(\brancher/_0688_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1316_  (.A(net368),
    .B(net366),
    .Y(\brancher/_0689_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1317_  (.A1(\brancher/_0641_ ),
    .A2(net368),
    .A3(\brancher/_0522_ ),
    .B1(net367),
    .X(\brancher/_0690_ ));
 sky130_fd_sc_hd__o211a_1 \brancher/_1318_  (.A1(\brancher/_0688_ ),
    .A2(\brancher/_0689_ ),
    .B1(\brancher/_0431_ ),
    .C1(\brancher/_0690_ ),
    .X(\brancher/_0691_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1319_  (.A(net945),
    .B(\brancher/_0691_ ),
    .Y(\brancher/_0692_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1320_  (.A(\brancher/_0687_ ),
    .B(\brancher/_0692_ ),
    .Y(\brancher/_0693_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1321_  (.A1(\brancher/rAlu_result[11] ),
    .A2(\brancher/_0587_ ),
    .B1(\brancher/_0434_ ),
    .X(\brancher/_0694_ ));
 sky130_fd_sc_hd__a22o_1 \brancher/_1322_  (.A1(\brancher/_0672_ ),
    .A2(\brancher/_0674_ ),
    .B1(\brancher/_0693_ ),
    .B2(\brancher/_0694_ ),
    .X(\wPcNextCond[11] ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1323_  (.A(\brancher/rPc_current_reg3[12] ),
    .B(\brancher/rAdder_jal[12] ),
    .Y(\brancher/_0695_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1324_  (.A(\brancher/rPc_current_reg3[12] ),
    .B(\brancher/rAdder_jal[12] ),
    .Y(\brancher/_0696_ ));
 sky130_fd_sc_hd__nand2b_1 \brancher/_1325_  (.A_N(\brancher/_0695_ ),
    .B(\brancher/_0696_ ),
    .Y(\brancher/_0697_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1326_  (.A1(\brancher/_0673_ ),
    .A2(\brancher/_0665_ ),
    .B1(\brancher/_0697_ ),
    .Y(\brancher/_0698_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1327_  (.A1(\brancher/_0673_ ),
    .A2(\brancher/_0665_ ),
    .A3(\brancher/_0697_ ),
    .B1(\brancher/_0458_ ),
    .X(\brancher/_0699_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1328_  (.A1(\brancher/rAlu_result[12] ),
    .A2(\brancher/_0457_ ),
    .B1(\brancher/_0459_ ),
    .Y(\brancher/_0700_ ));
 sky130_fd_sc_hd__xnor2_1 \brancher/_1329_  (.A(\brancher/rAdder_b[12] ),
    .B(\brancher/rPc_current_reg3[12] ),
    .Y(\brancher/_0701_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1330_  (.A(\brancher/_0701_ ),
    .Y(\brancher/_0702_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1331_  (.A(\brancher/_0685_ ),
    .B(\brancher/_0682_ ),
    .Y(\brancher/_0703_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1332_  (.A(\brancher/_0702_ ),
    .B(\brancher/_0703_ ),
    .X(\brancher/_0704_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1333_  (.A(\brancher/_0428_ ),
    .X(\brancher/_0705_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1334_  (.A(\brancher/_0703_ ),
    .B(\brancher/_0702_ ),
    .Y(\brancher/_0706_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1335_  (.A(\brancher/_0689_ ),
    .B(\brancher/_0688_ ),
    .Y(\brancher/_0707_ ));
 sky130_fd_sc_hd__xnor2_1 \brancher/_1336_  (.A(net363),
    .B(\brancher/_0707_ ),
    .Y(\brancher/_0708_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1337_  (.A1(\brancher/_0429_ ),
    .A2(\brancher/_0708_ ),
    .B1(\brancher/_0587_ ),
    .Y(\brancher/_0709_ ));
 sky130_fd_sc_hd__a31oi_1 \brancher/_1338_  (.A1(\brancher/_0704_ ),
    .A2(\brancher/_0705_ ),
    .A3(\brancher/_0706_ ),
    .B1(\brancher/_0709_ ),
    .Y(\brancher/_0710_ ));
 sky130_fd_sc_hd__o22ai_1 \brancher/_1339_  (.A1(\brancher/_0698_ ),
    .A2(\brancher/_0699_ ),
    .B1(\brancher/_0700_ ),
    .B2(\brancher/_0710_ ),
    .Y(\wPcNextCond[12] ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1340_  (.A(\brancher/_0666_ ),
    .B(\brancher/_0697_ ),
    .Y(\brancher/_0711_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1341_  (.A1(\brancher/_0616_ ),
    .A2(\brancher/_0661_ ),
    .B1(\brancher/_0659_ ),
    .Y(\brancher/_0712_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1342_  (.A(\brancher/_0712_ ),
    .B(\brancher/_0711_ ),
    .Y(\brancher/_0713_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1343_  (.A1(\brancher/_0665_ ),
    .A2(\brancher/_0695_ ),
    .B1(\brancher/_0696_ ),
    .X(\brancher/_0714_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1344_  (.A(\brancher/_0713_ ),
    .B(\brancher/_0714_ ),
    .Y(\brancher/_0715_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1345_  (.A1(\brancher/_0623_ ),
    .A2(\brancher/_0668_ ),
    .A3(\brancher/_0711_ ),
    .B1(\brancher/_0715_ ),
    .X(\brancher/_0716_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1346_  (.A(\brancher/_0716_ ),
    .Y(\brancher/_0717_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1347_  (.A(\brancher/rPc_current_reg3[13] ),
    .B(\brancher/rAdder_jal[13] ),
    .X(\brancher/_0718_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1348_  (.A(\brancher/rPc_current_reg3[13] ),
    .B(\brancher/rAdder_jal[13] ),
    .Y(\brancher/_0719_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1349_  (.A(\brancher/_0718_ ),
    .B(\brancher/_0719_ ),
    .Y(\brancher/_0720_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1350_  (.A(\brancher/_0720_ ),
    .B(\brancher/_0717_ ),
    .X(\brancher/_0721_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1351_  (.A(\brancher/_0721_ ),
    .B(net941),
    .Y(\brancher/_0722_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1352_  (.A1(\brancher/_0717_ ),
    .A2(\brancher/_0720_ ),
    .B1(\brancher/_0722_ ),
    .X(\brancher/_0723_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1353_  (.A(net929),
    .B(\brancher/rPc_current_reg3[13] ),
    .Y(\brancher/_0724_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1354_  (.A(net930),
    .B(\brancher/rPc_current_reg3[13] ),
    .Y(\brancher/_0725_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1355_  (.A(\brancher/_0725_ ),
    .Y(\brancher/_0726_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1356_  (.A(\brancher/_0724_ ),
    .B(\brancher/_0726_ ),
    .Y(\brancher/_0727_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1357_  (.A(\brancher/_0683_ ),
    .B(\brancher/_0701_ ),
    .Y(\brancher/_0728_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1358_  (.A(\brancher/_0684_ ),
    .B(\brancher/_0728_ ),
    .Y(\brancher/_0729_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1359_  (.A(\brancher/rAdder_b[12] ),
    .B(\brancher/rPc_current_reg3[12] ),
    .Y(\brancher/_0730_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1360_  (.A(\brancher/rAdder_b[12] ),
    .B(\brancher/rPc_current_reg3[12] ),
    .Y(\brancher/_0731_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1361_  (.A1(\brancher/_0682_ ),
    .A2(\brancher/_0730_ ),
    .B1(\brancher/_0731_ ),
    .X(\brancher/_0732_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1362_  (.A(\brancher/_0729_ ),
    .B(\brancher/_0732_ ),
    .Y(\brancher/_0733_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1363_  (.A(\brancher/_0727_ ),
    .B(\brancher/_0733_ ),
    .X(\brancher/_0734_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1364_  (.A(\brancher/_0733_ ),
    .B(\brancher/_0727_ ),
    .Y(\brancher/_0735_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1365_  (.A(\brancher/_0689_ ),
    .Y(\brancher/_0736_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1366_  (.A1(\brancher/_0643_ ),
    .A2(net363),
    .A3(\brancher/_0736_ ),
    .B1(net362),
    .X(\brancher/_0737_ ));
 sky130_fd_sc_hd__and3_1 \brancher/_1367_  (.A(\brancher/_0736_ ),
    .B(net364),
    .C(net362),
    .X(\brancher/_0738_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1368_  (.A(\brancher/_0643_ ),
    .B(\brancher/_0738_ ),
    .Y(\brancher/_0739_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1369_  (.A1(\brancher/_0737_ ),
    .A2(\brancher/_0431_ ),
    .A3(\brancher/_0739_ ),
    .B1(net945),
    .X(\brancher/_0740_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1370_  (.A1(\brancher/_0705_ ),
    .A2(\brancher/_0734_ ),
    .A3(\brancher/_0735_ ),
    .B1(\brancher/_0740_ ),
    .X(\brancher/_0741_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1371_  (.A1(\brancher/rAlu_result[13] ),
    .A2(\brancher/_0587_ ),
    .B1(\brancher/_0445_ ),
    .X(\brancher/_0742_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1372_  (.A(\brancher/_0741_ ),
    .B(\brancher/_0742_ ),
    .Y(\brancher/_0743_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1373_  (.A(\brancher/_0723_ ),
    .B(\brancher/_0743_ ),
    .Y(\wPcNextCond[13] ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1374_  (.A(net929),
    .B(\brancher/rPc_current_reg3[14] ),
    .Y(\brancher/_0744_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1375_  (.A(net929),
    .B(\brancher/rPc_current_reg3[14] ),
    .Y(\brancher/_0745_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1376_  (.A(\brancher/_0745_ ),
    .Y(\brancher/_0746_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1377_  (.A(\brancher/_0744_ ),
    .B(\brancher/_0746_ ),
    .Y(\brancher/_0747_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1378_  (.A(\brancher/_0747_ ),
    .Y(\brancher/_0748_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1379_  (.A1(\brancher/_0735_ ),
    .A2(\brancher/_0725_ ),
    .B1(\brancher/_0748_ ),
    .X(\brancher/_0749_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1380_  (.A(\brancher/_0735_ ),
    .B(\brancher/_0725_ ),
    .C(\brancher/_0748_ ),
    .Y(\brancher/_0750_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1381_  (.A(\brancher/_0749_ ),
    .B(\brancher/_0705_ ),
    .C(\brancher/_0750_ ),
    .Y(\brancher/_0751_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1382_  (.A(net360),
    .Y(\brancher/_0752_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1383_  (.A(\brancher/_0752_ ),
    .B(\brancher/_0739_ ),
    .Y(\brancher/_0753_ ));
 sky130_fd_sc_hd__buf_6 \brancher/_1384_  (.A(\brancher/_0753_ ),
    .X(\brancher/_0754_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1385_  (.A1(\brancher/_0739_ ),
    .A2(\brancher/_0752_ ),
    .B1(\brancher/_0535_ ),
    .X(\brancher/_0755_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1386_  (.A1(\brancher/_0754_ ),
    .A2(\brancher/_0755_ ),
    .B1(\brancher/_0456_ ),
    .X(\brancher/_0756_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1387_  (.A1(\brancher/rAlu_result[14] ),
    .A2(\brancher/_0608_ ),
    .B1(\brancher/_0445_ ),
    .Y(\brancher/_0757_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1388_  (.A1(\brancher/_0751_ ),
    .A2(\brancher/_0756_ ),
    .B1(\brancher/_0757_ ),
    .X(\brancher/_0758_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1389_  (.A(\brancher/_0721_ ),
    .B(\brancher/_0719_ ),
    .Y(\brancher/_0759_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1390_  (.A(\brancher/rPc_current_reg3[14] ),
    .B(\brancher/rAdder_jal[14] ),
    .X(\brancher/_0760_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1391_  (.A(\brancher/rPc_current_reg3[14] ),
    .B(\brancher/rAdder_jal[14] ),
    .Y(\brancher/_0761_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1392_  (.A(\brancher/_0760_ ),
    .B(\brancher/_0761_ ),
    .Y(\brancher/_0762_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1393_  (.A(\brancher/_0762_ ),
    .Y(\brancher/_0763_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1394_  (.A(\brancher/_0759_ ),
    .B(\brancher/_0763_ ),
    .Y(\brancher/_0764_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1395_  (.A(\brancher/_0721_ ),
    .B(\brancher/_0719_ ),
    .C(\brancher/_0762_ ),
    .Y(\brancher/_0765_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1396_  (.A(\brancher/_0764_ ),
    .B(net943),
    .C(\brancher/_0765_ ),
    .Y(\brancher/_0766_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1397_  (.A(\brancher/_0758_ ),
    .B(\brancher/_0766_ ),
    .Y(\wPcNextCond[14] ));
 sky130_fd_sc_hd__inv_2 \brancher/_1398_  (.A(net929),
    .Y(\brancher/_0767_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1399_  (.A(\brancher/rPc_current_reg3[15] ),
    .Y(\brancher/_0768_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1400_  (.A(\brancher/_0767_ ),
    .B(\brancher/_0768_ ),
    .Y(\brancher/_0769_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1401_  (.A(net929),
    .B(\brancher/rPc_current_reg3[15] ),
    .Y(\brancher/_0770_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1402_  (.A(\brancher/_0769_ ),
    .B(\brancher/_0770_ ),
    .Y(\brancher/_0771_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1403_  (.A(\brancher/_0771_ ),
    .Y(\brancher/_0772_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1404_  (.A(\brancher/_0727_ ),
    .B(\brancher/_0747_ ),
    .Y(\brancher/_0773_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1405_  (.A(\brancher/_0773_ ),
    .Y(\brancher/_0774_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1406_  (.A(\brancher/_0733_ ),
    .B(\brancher/_0774_ ),
    .Y(\brancher/_0775_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1407_  (.A(\brancher/_0725_ ),
    .B(\brancher/_0745_ ),
    .Y(\brancher/_0776_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1408_  (.A(\brancher/_0776_ ),
    .Y(\brancher/_0777_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1409_  (.A(\brancher/_0775_ ),
    .B(\brancher/_0777_ ),
    .Y(\brancher/_0778_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1410_  (.A(\brancher/_0772_ ),
    .B(\brancher/_0778_ ),
    .X(\brancher/_0779_ ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1411_  (.A(\brancher/_0551_ ),
    .X(\brancher/_0780_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1412_  (.A(\brancher/_0778_ ),
    .B(\brancher/_0772_ ),
    .Y(\brancher/_0781_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1413_  (.A(\brancher/_0779_ ),
    .B(\brancher/_0780_ ),
    .C(\brancher/_0781_ ),
    .Y(\brancher/_0782_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1414_  (.A(net357),
    .B(\brancher/_0754_ ),
    .Y(\brancher/_0783_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1415_  (.A(\brancher/_0754_ ),
    .B(net358),
    .Y(\brancher/_0784_ ));
 sky130_fd_sc_hd__or3b_1 \brancher/_1416_  (.A(\brancher/_0428_ ),
    .B(\brancher/_0783_ ),
    .C_N(\brancher/_0784_ ),
    .X(\brancher/_0785_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1417_  (.A(\brancher/_0782_ ),
    .B(\brancher/_0457_ ),
    .C(\brancher/_0785_ ),
    .Y(\brancher/_0786_ ));
 sky130_fd_sc_hd__buf_2 \brancher/_1418_  (.A(\brancher/_0433_ ),
    .X(\brancher/_0787_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1419_  (.A1(\brancher/rAlu_result[15] ),
    .A2(\brancher/_0608_ ),
    .B1(\brancher/_0787_ ),
    .X(\brancher/_0788_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1420_  (.A(\brancher/_0786_ ),
    .B(\brancher/_0788_ ),
    .Y(\brancher/_0789_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1421_  (.A(\brancher/rPc_current_reg3[15] ),
    .B(\brancher/rAdder_jal[15] ),
    .Y(\brancher/_0790_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1422_  (.A(\brancher/rPc_current_reg3[15] ),
    .B(\brancher/rAdder_jal[15] ),
    .Y(\brancher/_0791_ ));
 sky130_fd_sc_hd__nor2b_1 \brancher/_1423_  (.A(\brancher/_0790_ ),
    .B_N(\brancher/_0791_ ),
    .Y(\brancher/_0792_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1424_  (.A(\brancher/_0720_ ),
    .B(\brancher/_0762_ ),
    .Y(\brancher/_0793_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1425_  (.A(\brancher/_0716_ ),
    .B(\brancher/_0793_ ),
    .Y(\brancher/_0794_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1426_  (.A1(\brancher/_0719_ ),
    .A2(\brancher/_0762_ ),
    .B1(\brancher/_0761_ ),
    .Y(\brancher/_0795_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1427_  (.A(\brancher/_0795_ ),
    .Y(\brancher/_0796_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1428_  (.A(\brancher/_0794_ ),
    .B(\brancher/_0796_ ),
    .Y(\brancher/_0797_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1429_  (.A(\brancher/_0792_ ),
    .B(\brancher/_0797_ ),
    .X(\brancher/_0798_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1430_  (.A(\brancher/_0797_ ),
    .B(\brancher/_0792_ ),
    .Y(\brancher/_0799_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1431_  (.A(\brancher/_0798_ ),
    .B(net941),
    .C(\brancher/_0799_ ),
    .Y(\brancher/_0800_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1432_  (.A(\brancher/_0789_ ),
    .B(\brancher/_0800_ ),
    .Y(\wPcNextCond[15] ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1433_  (.A(\brancher/_0781_ ),
    .B(\brancher/_0770_ ),
    .Y(\brancher/_0801_ ));
 sky130_fd_sc_hd__inv_4 \brancher/_1434_  (.A(\brancher/rPc_current_reg3[16] ),
    .Y(\brancher/_0802_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1435_  (.A(\brancher/_0767_ ),
    .B(\brancher/_0802_ ),
    .Y(\brancher/_0803_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1436_  (.A(net929),
    .B(\brancher/rPc_current_reg3[16] ),
    .Y(\brancher/_0804_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1437_  (.A(\brancher/_0803_ ),
    .B(\brancher/_0804_ ),
    .Y(\brancher/_0805_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1438_  (.A(\brancher/_0805_ ),
    .Y(\brancher/_0806_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1439_  (.A(\brancher/_0801_ ),
    .B(\brancher/_0806_ ),
    .Y(\brancher/_0807_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1440_  (.A(\brancher/_0781_ ),
    .B(\brancher/_0770_ ),
    .C(\brancher/_0805_ ),
    .Y(\brancher/_0808_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1441_  (.A(\brancher/_0807_ ),
    .B(\brancher/_0430_ ),
    .C(\brancher/_0808_ ),
    .Y(\brancher/_0809_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1442_  (.A(net355),
    .Y(\brancher/_0810_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1443_  (.A(\brancher/_0810_ ),
    .B(\brancher/_0784_ ),
    .Y(\brancher/_0811_ ));
 sky130_fd_sc_hd__and2_1 \brancher/_1444_  (.A(\brancher/_0784_ ),
    .B(\brancher/_0810_ ),
    .X(\brancher/_0812_ ));
 sky130_fd_sc_hd__o31a_1 \brancher/_1445_  (.A1(\brancher/_0551_ ),
    .A2(\brancher/_0811_ ),
    .A3(\brancher/_0812_ ),
    .B1(\brancher/_0504_ ),
    .X(\brancher/_0813_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1446_  (.A(\brancher/_0809_ ),
    .B(\brancher/_0813_ ),
    .Y(\brancher/_0814_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1447_  (.A1(\brancher/rAlu_result[16] ),
    .A2(\brancher/_0608_ ),
    .B1(\brancher/_0787_ ),
    .X(\brancher/_0815_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1448_  (.A(\brancher/_0814_ ),
    .B(\brancher/_0815_ ),
    .Y(\brancher/_0816_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1449_  (.A(\brancher/_0799_ ),
    .B(\brancher/_0791_ ),
    .Y(\brancher/_0817_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1450_  (.A(\brancher/rAdder_jal[16] ),
    .Y(\brancher/_0818_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1451_  (.A(\brancher/_0802_ ),
    .B(\brancher/_0818_ ),
    .Y(\brancher/_0819_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1452_  (.A(\brancher/rPc_current_reg3[16] ),
    .B(\brancher/rAdder_jal[16] ),
    .Y(\brancher/_0820_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1453_  (.A(\brancher/_0819_ ),
    .B(\brancher/_0820_ ),
    .Y(\brancher/_0821_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1454_  (.A(\brancher/_0821_ ),
    .Y(\brancher/_0822_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1455_  (.A(\brancher/_0817_ ),
    .B(\brancher/_0822_ ),
    .Y(\brancher/_0823_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1456_  (.A(\brancher/_0799_ ),
    .B(\brancher/_0791_ ),
    .C(\brancher/_0821_ ),
    .Y(\brancher/_0824_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1457_  (.A(\brancher/_0823_ ),
    .B(net941),
    .C(\brancher/_0824_ ),
    .Y(\brancher/_0825_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1458_  (.A(\brancher/_0816_ ),
    .B(\brancher/_0825_ ),
    .Y(\wPcNextCond[16] ));
 sky130_fd_sc_hd__or2_1 \brancher/_1459_  (.A(net352),
    .B(\brancher/_0811_ ),
    .X(\brancher/_0826_ ));
 sky130_fd_sc_hd__and3_1 \brancher/_1460_  (.A(net358),
    .B(net355),
    .C(net352),
    .X(\brancher/_0827_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1461_  (.A1(\brancher/_0754_ ),
    .A2(\brancher/_0827_ ),
    .B1(\brancher/_0551_ ),
    .Y(\brancher/_0828_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1462_  (.A(\brancher/_0480_ ),
    .Y(\brancher/_0829_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1463_  (.A(net930),
    .B(\brancher/rPc_current_reg3[17] ),
    .Y(\brancher/_0830_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1464_  (.A(net930),
    .B(\brancher/rPc_current_reg3[17] ),
    .Y(\brancher/_0831_ ));
 sky130_fd_sc_hd__and2b_1 \brancher/_1465_  (.A_N(\brancher/_0830_ ),
    .B(\brancher/_0831_ ),
    .X(\brancher/_0832_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1466_  (.A(\brancher/_0675_ ),
    .B(\brancher/_0728_ ),
    .Y(\brancher/_0833_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1467_  (.A(\brancher/_0771_ ),
    .B(\brancher/_0805_ ),
    .Y(\brancher/_0834_ ));
 sky130_fd_sc_hd__nor2b_1 \brancher/_1468_  (.A(\brancher/_0773_ ),
    .B_N(\brancher/_0834_ ),
    .Y(\brancher/_0835_ ));
 sky130_fd_sc_hd__nor2b_1 \brancher/_1469_  (.A(\brancher/_0833_ ),
    .B_N(\brancher/_0835_ ),
    .Y(\brancher/_0836_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1470_  (.A(\brancher/_0637_ ),
    .B(\brancher/_0836_ ),
    .Y(\brancher/_0837_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1471_  (.A(\brancher/_0728_ ),
    .B(\brancher/_0677_ ),
    .Y(\brancher/_0838_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1472_  (.A(\brancher/_0838_ ),
    .B(\brancher/_0732_ ),
    .Y(\brancher/_0839_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1473_  (.A(\brancher/_0834_ ),
    .B(\brancher/_0776_ ),
    .Y(\brancher/_0840_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1474_  (.A(\brancher/_0840_ ),
    .B(\brancher/_0770_ ),
    .C(\brancher/_0804_ ),
    .Y(\brancher/_0841_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1475_  (.A1(\brancher/_0839_ ),
    .A2(\brancher/_0835_ ),
    .B1(\brancher/_0841_ ),
    .Y(\brancher/_0842_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1476_  (.A(\brancher/_0837_ ),
    .B(\brancher/_0842_ ),
    .Y(\brancher/_0843_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1477_  (.A(\brancher/_0832_ ),
    .B(\brancher/_0843_ ),
    .X(\brancher/_0844_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1478_  (.A(\brancher/_0843_ ),
    .B(\brancher/_0832_ ),
    .Y(\brancher/_0845_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1479_  (.A(\brancher/_0844_ ),
    .B(\brancher/_0845_ ),
    .Y(\brancher/_0846_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1480_  (.A(\brancher/_0605_ ),
    .B(\brancher/_0846_ ),
    .Y(\brancher/_0847_ ));
 sky130_fd_sc_hd__a211o_1 \brancher/_1481_  (.A1(\brancher/_0826_ ),
    .A2(\brancher/_0828_ ),
    .B1(\brancher/_0829_ ),
    .C1(\brancher/_0847_ ),
    .X(\brancher/_0848_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1482_  (.A(\brancher/rPc_current_reg3[17] ),
    .B(\brancher/rAdder_jal[17] ),
    .Y(\brancher/_0849_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1483_  (.A(\brancher/rPc_current_reg3[17] ),
    .B(\brancher/rAdder_jal[17] ),
    .Y(\brancher/_0850_ ));
 sky130_fd_sc_hd__and2b_1 \brancher/_1484_  (.A_N(\brancher/_0849_ ),
    .B(\brancher/_0850_ ),
    .X(\brancher/_0851_ ));
 sky130_fd_sc_hd__and2_1 \brancher/_1485_  (.A(\brancher/_0792_ ),
    .B(\brancher/_0822_ ),
    .X(\brancher/_0852_ ));
 sky130_fd_sc_hd__and2_1 \brancher/_1486_  (.A(\brancher/_0852_ ),
    .B(\brancher/_0793_ ),
    .X(\brancher/_0853_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1487_  (.A1(\brancher/_0791_ ),
    .A2(\brancher/_0821_ ),
    .B1(\brancher/_0820_ ),
    .Y(\brancher/_0854_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1488_  (.A1(\brancher/_0795_ ),
    .A2(\brancher/_0852_ ),
    .B1(\brancher/_0854_ ),
    .X(\brancher/_0855_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1489_  (.A1(\brancher/_0715_ ),
    .A2(\brancher/_0853_ ),
    .B1(\brancher/_0855_ ),
    .Y(\brancher/_0856_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1490_  (.A(\brancher/_0668_ ),
    .B(\brancher/_0711_ ),
    .Y(\brancher/_0857_ ));
 sky130_fd_sc_hd__nor2b_1 \brancher/_1491_  (.A(\brancher/_0857_ ),
    .B_N(\brancher/_0853_ ),
    .Y(\brancher/_0858_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1492_  (.A(\brancher/_0623_ ),
    .B(\brancher/_0858_ ),
    .Y(\brancher/_0859_ ));
 sky130_fd_sc_hd__nand2_2 \brancher/_1493_  (.A(\brancher/_0856_ ),
    .B(\brancher/_0859_ ),
    .Y(\brancher/_0860_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1494_  (.A(\brancher/_0851_ ),
    .B(\brancher/_0860_ ),
    .X(\brancher/_0861_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1495_  (.A(\brancher/_0860_ ),
    .B(\brancher/_0851_ ),
    .Y(\brancher/_0862_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1496_  (.A1(\brancher/_0861_ ),
    .A2(\brancher/_0862_ ),
    .B1(\brancher/_0787_ ),
    .X(\brancher/_0863_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1497_  (.A(\brancher/rAlu_result[17] ),
    .B(\brancher/_0438_ ),
    .X(\brancher/_0864_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1498_  (.A(\brancher/_0848_ ),
    .B(\brancher/_0863_ ),
    .C(\brancher/_0864_ ),
    .Y(\brancher/_0865_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1499_  (.A(\brancher/_0865_ ),
    .Y(\wPcNextCond[17] ));
 sky130_fd_sc_hd__xor2_1 \brancher/_1500_  (.A(net931),
    .B(\brancher/rPc_current_reg3[18] ),
    .X(\brancher/_0866_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1501_  (.A(\brancher/_0845_ ),
    .B(\brancher/_0831_ ),
    .Y(\brancher/_0867_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1502_  (.A(\brancher/_0866_ ),
    .B(\brancher/_0867_ ),
    .X(\brancher/_0868_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1503_  (.A(\brancher/_0867_ ),
    .B(\brancher/_0866_ ),
    .Y(\brancher/_0869_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1504_  (.A(\brancher/_0868_ ),
    .B(\brancher/_0705_ ),
    .C(\brancher/_0869_ ),
    .Y(\brancher/_0870_ ));
 sky130_fd_sc_hd__and4_1 \brancher/_1505_  (.A(net361),
    .B(net358),
    .C(net355),
    .D(net352),
    .X(\brancher/_0871_ ));
 sky130_fd_sc_hd__and3_1 \brancher/_1506_  (.A(\brancher/_0642_ ),
    .B(\brancher/_0738_ ),
    .C(\brancher/_0871_ ),
    .X(\brancher/_0872_ ));
 sky130_fd_sc_hd__buf_2 \brancher/_1507_  (.A(\brancher/_0872_ ),
    .X(\brancher/_0873_ ));
 sky130_fd_sc_hd__xor2_1 \brancher/_1508_  (.A(net350),
    .B(\brancher/_0873_ ),
    .X(\brancher/_0874_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1509_  (.A1(\brancher/_0874_ ),
    .A2(\brancher/_0605_ ),
    .B1(net945),
    .Y(\brancher/_0875_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1510_  (.A(\brancher/_0870_ ),
    .B(\brancher/_0875_ ),
    .Y(\brancher/_0876_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1511_  (.A1(\brancher/rAlu_result[18] ),
    .A2(\brancher/_0504_ ),
    .B1(\brancher/_0434_ ),
    .X(\brancher/_0877_ ));
 sky130_fd_sc_hd__and2_1 \brancher/_1512_  (.A(\brancher/_0862_ ),
    .B(\brancher/_0850_ ),
    .X(\brancher/_0878_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1513_  (.A(\brancher/rPc_current_reg3[18] ),
    .B(\brancher/rAdder_jal[18] ),
    .Y(\brancher/_0879_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1514_  (.A(\brancher/rPc_current_reg3[18] ),
    .B(\brancher/rAdder_jal[18] ),
    .Y(\brancher/_0880_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1515_  (.A(\brancher/_0880_ ),
    .Y(\brancher/_0881_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1516_  (.A(\brancher/_0879_ ),
    .B(\brancher/_0881_ ),
    .Y(\brancher/_0882_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1517_  (.A(\brancher/_0882_ ),
    .Y(\brancher/_0883_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1518_  (.A(\brancher/_0878_ ),
    .B(\brancher/_0883_ ),
    .Y(\brancher/_0884_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1519_  (.A(\brancher/_0883_ ),
    .B(\brancher/_0878_ ),
    .Y(\brancher/_0885_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1520_  (.A(\brancher/_0459_ ),
    .B(\brancher/_0885_ ),
    .Y(\brancher/_0886_ ));
 sky130_fd_sc_hd__a22o_1 \brancher/_1521_  (.A1(\brancher/_0876_ ),
    .A2(\brancher/_0877_ ),
    .B1(\brancher/_0884_ ),
    .B2(\brancher/_0886_ ),
    .X(\wPcNextCond[18] ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1522_  (.A(net932),
    .B(\brancher/rPc_current_reg3[19] ),
    .Y(\brancher/_0887_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1523_  (.A(net932),
    .B(\brancher/rPc_current_reg3[19] ),
    .Y(\brancher/_0888_ ));
 sky130_fd_sc_hd__and2b_1 \brancher/_1524_  (.A_N(\brancher/_0887_ ),
    .B(\brancher/_0888_ ),
    .X(\brancher/_0889_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1525_  (.A(\brancher/_0832_ ),
    .B(\brancher/_0866_ ),
    .Y(\brancher/_0890_ ));
 sky130_fd_sc_hd__and2_1 \brancher/_1526_  (.A(\brancher/_0837_ ),
    .B(\brancher/_0842_ ),
    .X(\brancher/_0891_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1527_  (.A1(\brancher/rPc_current_reg3[17] ),
    .A2(\brancher/rPc_current_reg3[18] ),
    .B1(net931),
    .X(\brancher/_0892_ ));
 sky130_fd_sc_hd__o21bai_1 \brancher/_1528_  (.A1(\brancher/_0890_ ),
    .A2(\brancher/_0891_ ),
    .B1_N(\brancher/_0892_ ),
    .Y(\brancher/_0893_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1529_  (.A(\brancher/_0889_ ),
    .B(\brancher/_0893_ ),
    .X(\brancher/_0894_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1530_  (.A(\brancher/_0893_ ),
    .B(\brancher/_0889_ ),
    .Y(\brancher/_0895_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1531_  (.A(\brancher/_0894_ ),
    .B(\brancher/_0705_ ),
    .C(\brancher/_0895_ ),
    .Y(\brancher/_0896_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1532_  (.A(\brancher/_0873_ ),
    .B(net350),
    .Y(\brancher/_0897_ ));
 sky130_fd_sc_hd__xnor2_1 \brancher/_1533_  (.A(net348),
    .B(\brancher/_0897_ ),
    .Y(\brancher/_0898_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1534_  (.A1(\brancher/_0898_ ),
    .A2(\brancher/_0605_ ),
    .B1(net945),
    .Y(\brancher/_0899_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1535_  (.A1(\brancher/rAlu_result[19] ),
    .A2(\brancher/_0608_ ),
    .B1(\brancher/_0445_ ),
    .Y(\brancher/_0900_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1536_  (.A1(\brancher/_0896_ ),
    .A2(\brancher/_0899_ ),
    .B1(\brancher/_0900_ ),
    .X(\brancher/_0901_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1537_  (.A(\brancher/rPc_current_reg3[19] ),
    .B(\brancher/rAdder_jal[19] ),
    .Y(\brancher/_0902_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1538_  (.A(\brancher/rPc_current_reg3[19] ),
    .B(\brancher/rAdder_jal[19] ),
    .Y(\brancher/_0903_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1539_  (.A(\brancher/_0903_ ),
    .Y(\brancher/_0904_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1540_  (.A(\brancher/_0902_ ),
    .B(\brancher/_0904_ ),
    .Y(\brancher/_0905_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1541_  (.A(\brancher/_0851_ ),
    .B(\brancher/_0882_ ),
    .Y(\brancher/_0906_ ));
 sky130_fd_sc_hd__nand2b_1 \brancher/_1542_  (.A_N(\brancher/_0906_ ),
    .B(\brancher/_0860_ ),
    .Y(\brancher/_0907_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1543_  (.A1(\brancher/_0850_ ),
    .A2(\brancher/_0880_ ),
    .B1(\brancher/_0879_ ),
    .Y(\brancher/_0908_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1544_  (.A(\brancher/_0908_ ),
    .Y(\brancher/_0909_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1545_  (.A(\brancher/_0907_ ),
    .B(\brancher/_0909_ ),
    .Y(\brancher/_0910_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1546_  (.A(\brancher/_0905_ ),
    .B(\brancher/_0910_ ),
    .X(\brancher/_0911_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1547_  (.A(\brancher/_0910_ ),
    .B(\brancher/_0905_ ),
    .Y(\brancher/_0912_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1548_  (.A(\brancher/_0911_ ),
    .B(net941),
    .C(\brancher/_0912_ ),
    .Y(\brancher/_0913_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1549_  (.A(\brancher/_0901_ ),
    .B(\brancher/_0913_ ),
    .Y(\wPcNextCond[19] ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1550_  (.A(\brancher/rPc_current_reg3[20] ),
    .B(\brancher/rAdder_jal[20] ),
    .Y(\brancher/_0914_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1551_  (.A(\brancher/rPc_current_reg3[20] ),
    .B(\brancher/rAdder_jal[20] ),
    .Y(\brancher/_0915_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1552_  (.A(\brancher/_0915_ ),
    .Y(\brancher/_0916_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1553_  (.A(\brancher/_0914_ ),
    .B(\brancher/_0916_ ),
    .Y(\brancher/_0917_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1554_  (.A(\brancher/_0912_ ),
    .B(\brancher/_0903_ ),
    .Y(\brancher/_0918_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1555_  (.A(\brancher/_0917_ ),
    .B(\brancher/_0918_ ),
    .X(\brancher/_0919_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1556_  (.A(\brancher/_0918_ ),
    .B(\brancher/_0917_ ),
    .Y(\brancher/_0920_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1557_  (.A(\brancher/_0919_ ),
    .B(net939),
    .C(\brancher/_0920_ ),
    .Y(\brancher/_0921_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1558_  (.A(net932),
    .B(\brancher/rPc_current_reg3[20] ),
    .Y(\brancher/_0922_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1559_  (.A(net932),
    .B(\brancher/rPc_current_reg3[20] ),
    .Y(\brancher/_0923_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1560_  (.A(\brancher/_0923_ ),
    .Y(\brancher/_0924_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1561_  (.A(\brancher/_0922_ ),
    .B(\brancher/_0924_ ),
    .Y(\brancher/_0925_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1562_  (.A(\brancher/_0925_ ),
    .Y(\brancher/_0926_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1563_  (.A1(\brancher/_0895_ ),
    .A2(\brancher/_0888_ ),
    .B1(\brancher/_0926_ ),
    .Y(\brancher/_0927_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1564_  (.A(\brancher/_0895_ ),
    .B(\brancher/_0888_ ),
    .C(\brancher/_0926_ ),
    .Y(\brancher/_0928_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1565_  (.A(\brancher/_0928_ ),
    .B(\brancher/_0705_ ),
    .Y(\brancher/_0929_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1566_  (.A(net347),
    .Y(\brancher/_0930_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1567_  (.A(net351),
    .B(net348),
    .Y(\brancher/_0931_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1568_  (.A(\brancher/_0930_ ),
    .B(\brancher/_0931_ ),
    .Y(\brancher/_0932_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1569_  (.A(\brancher/_0754_ ),
    .B(\brancher/_0827_ ),
    .C(\brancher/_0932_ ),
    .Y(\brancher/_0933_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1570_  (.A(\brancher/_0933_ ),
    .B(\brancher/_0431_ ),
    .Y(\brancher/_0934_ ));
 sky130_fd_sc_hd__and3_1 \brancher/_1571_  (.A(\brancher/_0754_ ),
    .B(net351),
    .C(\brancher/_0827_ ),
    .X(\brancher/_0935_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1572_  (.A1(\brancher/_0935_ ),
    .A2(net349),
    .B1(net347),
    .Y(\brancher/_0936_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1573_  (.A1(\brancher/_0934_ ),
    .A2(\brancher/_0936_ ),
    .B1(\brancher/_0504_ ),
    .X(\brancher/_0937_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1574_  (.A1(\brancher/_0927_ ),
    .A2(\brancher/_0929_ ),
    .B1(\brancher/_0937_ ),
    .Y(\brancher/_0938_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1575_  (.A1(\brancher/rAlu_result[20] ),
    .A2(\brancher/_0587_ ),
    .B1(\brancher/_0445_ ),
    .X(\brancher/_0939_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1576_  (.A(\brancher/_0938_ ),
    .B(\brancher/_0939_ ),
    .Y(\brancher/_0940_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1577_  (.A(\brancher/_0921_ ),
    .B(\brancher/_0940_ ),
    .Y(\wPcNextCond[20] ));
 sky130_fd_sc_hd__clkbuf_2 \brancher/_1578_  (.A(\brancher/_0605_ ),
    .X(\brancher/_0941_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1579_  (.A(net932),
    .B(net958),
    .Y(\brancher/_0942_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1580_  (.A(net932),
    .B(net958),
    .Y(\brancher/_0943_ ));
 sky130_fd_sc_hd__and2b_1 \brancher/_1581_  (.A_N(\brancher/_0942_ ),
    .B(\brancher/_0943_ ),
    .X(\brancher/_0944_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1582_  (.A(\brancher/_0889_ ),
    .B(\brancher/_0925_ ),
    .Y(\brancher/_0945_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1583_  (.A(\brancher/_0945_ ),
    .B(\brancher/_0890_ ),
    .Y(\brancher/_0946_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1584_  (.A(\brancher/_0843_ ),
    .B(\brancher/_0946_ ),
    .Y(\brancher/_0947_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1585_  (.A(\brancher/_0888_ ),
    .B(\brancher/_0923_ ),
    .Y(\brancher/_0948_ ));
 sky130_fd_sc_hd__a31o_1 \brancher/_1586_  (.A1(\brancher/_0889_ ),
    .A2(\brancher/_0892_ ),
    .A3(\brancher/_0925_ ),
    .B1(\brancher/_0948_ ),
    .X(\brancher/_0949_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1587_  (.A(\brancher/_0949_ ),
    .Y(\brancher/_0950_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1588_  (.A(\brancher/_0947_ ),
    .B(\brancher/_0950_ ),
    .Y(\brancher/_0951_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1589_  (.A(\brancher/_0944_ ),
    .B(\brancher/_0951_ ),
    .X(\brancher/_0952_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1590_  (.A(\brancher/_0951_ ),
    .B(\brancher/_0944_ ),
    .Y(\brancher/_0953_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1591_  (.A(\brancher/_0952_ ),
    .B(\brancher/_0953_ ),
    .Y(\brancher/_0954_ ));
 sky130_fd_sc_hd__or2b_1 \brancher/_1592_  (.A(net345),
    .B_N(\brancher/_0933_ ),
    .X(\brancher/_0955_ ));
 sky130_fd_sc_hd__and2_1 \brancher/_1593_  (.A(\brancher/_0932_ ),
    .B(net345),
    .X(\brancher/_0956_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1594_  (.A(\brancher/_0753_ ),
    .B(\brancher/_0827_ ),
    .C(\brancher/_0956_ ),
    .Y(\brancher/_0957_ ));
 sky130_fd_sc_hd__a31oi_1 \brancher/_1595_  (.A1(\brancher/_0955_ ),
    .A2(\brancher/_0605_ ),
    .A3(\brancher/_0957_ ),
    .B1(\brancher/_0829_ ),
    .Y(\brancher/_0958_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1596_  (.A1(\brancher/_0941_ ),
    .A2(\brancher/_0954_ ),
    .B1(\brancher/_0958_ ),
    .Y(\brancher/_0959_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1597_  (.A(net958),
    .B(net948),
    .Y(\brancher/_0960_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1598_  (.A(net958),
    .B(net948),
    .Y(\brancher/_0961_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1599_  (.A(\brancher/_0961_ ),
    .Y(\brancher/_0962_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1600_  (.A(\brancher/_0960_ ),
    .B(\brancher/_0962_ ),
    .Y(\brancher/_0963_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1601_  (.A(\brancher/_0905_ ),
    .B(\brancher/_0917_ ),
    .Y(\brancher/_0964_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1602_  (.A(\brancher/_0964_ ),
    .B(\brancher/_0906_ ),
    .Y(\brancher/_0965_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1603_  (.A(\brancher/_0860_ ),
    .B(\brancher/_0965_ ),
    .Y(\brancher/_0966_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1604_  (.A(\brancher/_0917_ ),
    .B(\brancher/_0904_ ),
    .Y(\brancher/_0967_ ));
 sky130_fd_sc_hd__o211a_1 \brancher/_1605_  (.A1(\brancher/_0964_ ),
    .A2(\brancher/_0909_ ),
    .B1(\brancher/_0915_ ),
    .C1(\brancher/_0967_ ),
    .X(\brancher/_0968_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1606_  (.A(\brancher/_0966_ ),
    .B(\brancher/_0968_ ),
    .Y(\brancher/_0969_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1607_  (.A(\brancher/_0963_ ),
    .B(\brancher/_0969_ ),
    .X(\brancher/_0970_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1608_  (.A(\brancher/_0969_ ),
    .B(\brancher/_0963_ ),
    .Y(\brancher/_0971_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1609_  (.A(\brancher/_0970_ ),
    .B(\brancher/_0971_ ),
    .Y(\brancher/_0972_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1610_  (.A(\brancher/_0972_ ),
    .B(net939),
    .Y(\brancher/_0973_ ));
 sky130_fd_sc_hd__o211ai_2 \brancher/_1611_  (.A1(\brancher/rAlu_result[21] ),
    .A2(\brancher/_0438_ ),
    .B1(\brancher/_0959_ ),
    .C1(\brancher/_0973_ ),
    .Y(\brancher/_0974_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1612_  (.A(\brancher/_0974_ ),
    .Y(\wPcNextCond[21] ));
 sky130_fd_sc_hd__xor2_1 \brancher/_1613_  (.A(net933),
    .B(\brancher/rPc_current_reg3[22] ),
    .X(\brancher/_0975_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1614_  (.A(\brancher/_0953_ ),
    .B(\brancher/_0943_ ),
    .Y(\brancher/_0976_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1615_  (.A(\brancher/_0975_ ),
    .B(\brancher/_0976_ ),
    .X(\brancher/_0977_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1616_  (.A(\brancher/_0976_ ),
    .B(\brancher/_0975_ ),
    .Y(\brancher/_0978_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1617_  (.A(\brancher/_0977_ ),
    .B(\brancher/_0430_ ),
    .C(\brancher/_0978_ ),
    .Y(\brancher/_0979_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1618_  (.A(net343),
    .Y(\brancher/_0980_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1619_  (.A1(\brancher/_0957_ ),
    .A2(\brancher/_0980_ ),
    .B1(\brancher/_0429_ ),
    .Y(\brancher/_0981_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1620_  (.A(\brancher/_0980_ ),
    .B(\brancher/_0957_ ),
    .X(\brancher/_0982_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1621_  (.A1(\brancher/_0981_ ),
    .A2(\brancher/_0982_ ),
    .B1(net945),
    .Y(\brancher/_0983_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1622_  (.A(\brancher/_0979_ ),
    .B(\brancher/_0983_ ),
    .Y(\brancher/_0984_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1623_  (.A1(\brancher/rAlu_result[22] ),
    .A2(\brancher/_0608_ ),
    .B1(\brancher/_0787_ ),
    .X(\brancher/_0985_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1624_  (.A(\brancher/_0984_ ),
    .B(\brancher/_0985_ ),
    .Y(\brancher/_0986_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1625_  (.A(net948),
    .B(\brancher/rPc_current_reg3[22] ),
    .Y(\brancher/_0987_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1626_  (.A(net948),
    .B(\brancher/rPc_current_reg3[22] ),
    .Y(\brancher/_0988_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1627_  (.A(\brancher/_0988_ ),
    .Y(\brancher/_0989_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1628_  (.A(\brancher/_0987_ ),
    .B(\brancher/_0989_ ),
    .Y(\brancher/_0990_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1629_  (.A(\brancher/_0971_ ),
    .B(\brancher/_0961_ ),
    .Y(\brancher/_0991_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1630_  (.A(\brancher/_0990_ ),
    .B(\brancher/_0991_ ),
    .X(\brancher/_0992_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1631_  (.A(\brancher/_0991_ ),
    .B(\brancher/_0990_ ),
    .Y(\brancher/_0993_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1632_  (.A(\brancher/_0992_ ),
    .B(net939),
    .C(\brancher/_0993_ ),
    .Y(\brancher/_0994_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1633_  (.A(\brancher/_0986_ ),
    .B(\brancher/_0994_ ),
    .Y(\wPcNextCond[22] ));
 sky130_fd_sc_hd__xnor2_1 \brancher/_1634_  (.A(net342),
    .B(\brancher/_0982_ ),
    .Y(\brancher/_0995_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1635_  (.A1(\brancher/_0995_ ),
    .A2(\brancher/_0941_ ),
    .B1(net945),
    .Y(\brancher/_0996_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1636_  (.A(net933),
    .B(\brancher/rPc_current_reg3[23] ),
    .Y(\brancher/_0997_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1637_  (.A(net933),
    .B(\brancher/rPc_current_reg3[23] ),
    .Y(\brancher/_0998_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1638_  (.A(\brancher/_0998_ ),
    .Y(\brancher/_0999_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1639_  (.A(\brancher/_0997_ ),
    .B(\brancher/_0999_ ),
    .Y(\brancher/_1000_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1640_  (.A(\brancher/_0944_ ),
    .B(\brancher/_0975_ ),
    .Y(\brancher/_1001_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1641_  (.A(\brancher/_1001_ ),
    .Y(\brancher/_1002_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1642_  (.A(\brancher/_0951_ ),
    .B(\brancher/_1002_ ),
    .Y(\brancher/_1003_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1643_  (.A1(net958),
    .A2(\brancher/rPc_current_reg3[22] ),
    .B1(net933),
    .Y(\brancher/_1004_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1644_  (.A(\brancher/_1003_ ),
    .B(\brancher/_1004_ ),
    .Y(\brancher/_1005_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1645_  (.A(\brancher/_1000_ ),
    .B(\brancher/_1005_ ),
    .X(\brancher/_1006_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1646_  (.A(\brancher/_1005_ ),
    .B(\brancher/_1000_ ),
    .Y(\brancher/_1007_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1647_  (.A(\brancher/_1006_ ),
    .B(\brancher/_0780_ ),
    .C(\brancher/_1007_ ),
    .Y(\brancher/_1008_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1648_  (.A(\brancher/_0996_ ),
    .B(\brancher/_1008_ ),
    .Y(\brancher/_1009_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \brancher/_1649_  (.A(\brancher/_0440_ ),
    .X(\brancher/_0096_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1650_  (.A1(\brancher/rAlu_result[23] ),
    .A2(\brancher/_0096_ ),
    .B1(\brancher/_0787_ ),
    .X(\brancher/_0097_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1651_  (.A(\brancher/_1009_ ),
    .B(\brancher/_0097_ ),
    .Y(\brancher/_0098_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1652_  (.A(net948),
    .B(\brancher/rPc_current_reg3[23] ),
    .Y(\brancher/_0099_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1653_  (.A(net948),
    .B(\brancher/rPc_current_reg3[23] ),
    .Y(\brancher/_0100_ ));
 sky130_fd_sc_hd__and2b_1 \brancher/_1654_  (.A_N(\brancher/_0099_ ),
    .B(\brancher/_0100_ ),
    .X(\brancher/_0101_ ));
 sky130_fd_sc_hd__and2_1 \brancher/_1655_  (.A(\brancher/_0963_ ),
    .B(\brancher/_0990_ ),
    .X(\brancher/_0102_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1656_  (.A(\brancher/_0969_ ),
    .B(\brancher/_0102_ ),
    .Y(\brancher/_0103_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1657_  (.A(\brancher/_0962_ ),
    .B(\brancher/_0989_ ),
    .Y(\brancher/_0104_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1658_  (.A(\brancher/_0103_ ),
    .B(\brancher/_0104_ ),
    .Y(\brancher/_0105_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1659_  (.A(\brancher/_0101_ ),
    .B(\brancher/_0105_ ),
    .X(\brancher/_0106_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1660_  (.A(\brancher/_0105_ ),
    .B(\brancher/_0101_ ),
    .Y(\brancher/_0107_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1661_  (.A(\brancher/_0106_ ),
    .B(net939),
    .C(\brancher/_0107_ ),
    .Y(\brancher/_0108_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1662_  (.A(\brancher/_0098_ ),
    .B(\brancher/_0108_ ),
    .Y(\wPcNextCond[23] ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1663_  (.A(\brancher/_1007_ ),
    .B(\brancher/_0998_ ),
    .Y(\brancher/_0109_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1664_  (.A(net933),
    .B(\brancher/rPc_current_reg3[24] ),
    .Y(\brancher/_0110_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1665_  (.A(net933),
    .B(\brancher/rPc_current_reg3[24] ),
    .Y(\brancher/_0111_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1666_  (.A(\brancher/_0111_ ),
    .Y(\brancher/_0112_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1667_  (.A(\brancher/_0110_ ),
    .B(\brancher/_0112_ ),
    .Y(\brancher/_0113_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1668_  (.A(\brancher/_0109_ ),
    .B(\brancher/_0113_ ),
    .Y(\brancher/_0114_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1669_  (.A(\brancher/_0113_ ),
    .Y(\brancher/_0115_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1670_  (.A(\brancher/_1007_ ),
    .B(\brancher/_0998_ ),
    .C(\brancher/_0115_ ),
    .Y(\brancher/_0116_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1671_  (.A(\brancher/_0114_ ),
    .B(\brancher/_0430_ ),
    .C(\brancher/_0116_ ),
    .Y(\brancher/_0117_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1672_  (.A(net340),
    .Y(\brancher/_0118_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1673_  (.A(net344),
    .B(net342),
    .Y(\brancher/_0119_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1674_  (.A(\brancher/_0119_ ),
    .Y(\brancher/_0120_ ));
 sky130_fd_sc_hd__nand3_2 \brancher/_1675_  (.A(\brancher/_0873_ ),
    .B(\brancher/_0956_ ),
    .C(\brancher/_0120_ ),
    .Y(\brancher/_0121_ ));
 sky130_fd_sc_hd__xor2_1 \brancher/_1676_  (.A(\brancher/_0118_ ),
    .B(\brancher/_0121_ ),
    .X(\brancher/_0122_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1677_  (.A1(\brancher/_0122_ ),
    .A2(\brancher/_0432_ ),
    .B1(net946),
    .Y(\brancher/_0123_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1678_  (.A(\brancher/_0117_ ),
    .B(\brancher/_0123_ ),
    .Y(\brancher/_0124_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1679_  (.A1(\brancher/rAlu_result[24] ),
    .A2(\brancher/_0096_ ),
    .B1(\brancher/_0588_ ),
    .X(\brancher/_0125_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1680_  (.A(\brancher/_0124_ ),
    .B(\brancher/_0125_ ),
    .Y(\brancher/_0126_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1681_  (.A(\brancher/_0107_ ),
    .B(\brancher/_0100_ ),
    .Y(\brancher/_0127_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1682_  (.A(net949),
    .B(\brancher/rPc_current_reg3[24] ),
    .Y(\brancher/_0128_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1683_  (.A(net949),
    .B(\brancher/rPc_current_reg3[24] ),
    .Y(\brancher/_0129_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1684_  (.A(\brancher/_0129_ ),
    .Y(\brancher/_0130_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1685_  (.A(\brancher/_0128_ ),
    .B(\brancher/_0130_ ),
    .Y(\brancher/_0131_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1686_  (.A(\brancher/_0127_ ),
    .B(\brancher/_0131_ ),
    .Y(\brancher/_0132_ ));
 sky130_fd_sc_hd__nand3b_1 \brancher/_1687_  (.A_N(\brancher/_0131_ ),
    .B(\brancher/_0107_ ),
    .C(\brancher/_0100_ ),
    .Y(\brancher/_0133_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1688_  (.A(\brancher/_0132_ ),
    .B(\brancher/_0133_ ),
    .C(net939),
    .Y(\brancher/_0134_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1689_  (.A(\brancher/_0126_ ),
    .B(\brancher/_0134_ ),
    .Y(\wPcNextCond[24] ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1690_  (.A(net949),
    .B(net957),
    .Y(\brancher/_0135_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1691_  (.A(net949),
    .B(net957),
    .Y(\brancher/_0136_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1692_  (.A(\brancher/_0136_ ),
    .Y(\brancher/_0137_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1693_  (.A(\brancher/_0135_ ),
    .B(\brancher/_0137_ ),
    .Y(\brancher/_0138_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1694_  (.A(\brancher/_0102_ ),
    .B(\brancher/_0101_ ),
    .C(\brancher/_0131_ ),
    .Y(\brancher/_0139_ ));
 sky130_fd_sc_hd__o41a_1 \brancher/_1695_  (.A1(\brancher/rPc_current_reg3[21] ),
    .A2(\brancher/rPc_current_reg3[22] ),
    .A3(\brancher/rPc_current_reg3[23] ),
    .A4(\brancher/rPc_current_reg3[24] ),
    .B1(net950),
    .X(\brancher/_0140_ ));
 sky130_fd_sc_hd__o21ba_1 \brancher/_1696_  (.A1(\brancher/_0968_ ),
    .A2(\brancher/_0139_ ),
    .B1_N(\brancher/_0140_ ),
    .X(\brancher/_0141_ ));
 sky130_fd_sc_hd__and2b_1 \brancher/_1697_  (.A_N(\brancher/_0139_ ),
    .B(\brancher/_0965_ ),
    .X(\brancher/_0142_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1698_  (.A(\brancher/_0860_ ),
    .B(\brancher/_0142_ ),
    .Y(\brancher/_0143_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1699_  (.A(\brancher/_0141_ ),
    .B(\brancher/_0143_ ),
    .Y(\brancher/_0144_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1700_  (.A(\brancher/_0138_ ),
    .B(\brancher/_0144_ ),
    .X(\brancher/_0145_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1701_  (.A(\brancher/_0144_ ),
    .B(\brancher/_0138_ ),
    .Y(\brancher/_0146_ ));
 sky130_fd_sc_hd__a21o_1 \brancher/_1702_  (.A1(\brancher/_0145_ ),
    .A2(\brancher/_0146_ ),
    .B1(\brancher/_0787_ ),
    .X(\brancher/_0147_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1703_  (.A(net934),
    .B(net957),
    .Y(\brancher/_0148_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1704_  (.A(net934),
    .B(net957),
    .Y(\brancher/_0149_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1705_  (.A(\brancher/_0149_ ),
    .Y(\brancher/_0150_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1706_  (.A(\brancher/_0148_ ),
    .B(\brancher/_0150_ ),
    .Y(\brancher/_0151_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1707_  (.A(\brancher/_1000_ ),
    .B(\brancher/_0113_ ),
    .Y(\brancher/_0152_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1708_  (.A(\brancher/_0152_ ),
    .B(\brancher/_1001_ ),
    .Y(\brancher/_0153_ ));
 sky130_fd_sc_hd__and2_1 \brancher/_1709_  (.A(\brancher/_0946_ ),
    .B(\brancher/_0153_ ),
    .X(\brancher/_0154_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1710_  (.A(\brancher/_0843_ ),
    .B(\brancher/_0154_ ),
    .Y(\brancher/_0155_ ));
 sky130_fd_sc_hd__or3b_1 \brancher/_1711_  (.A(\brancher/_0999_ ),
    .B(\brancher/_0112_ ),
    .C_N(\brancher/_1004_ ),
    .X(\brancher/_0156_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1712_  (.A1(\brancher/_0949_ ),
    .A2(\brancher/_0153_ ),
    .B1(\brancher/_0156_ ),
    .Y(\brancher/_0157_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1713_  (.A(\brancher/_0155_ ),
    .B(\brancher/_0157_ ),
    .Y(\brancher/_0158_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1714_  (.A(\brancher/_0151_ ),
    .B(\brancher/_0158_ ),
    .X(\brancher/_0159_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1715_  (.A(\brancher/_0158_ ),
    .B(\brancher/_0151_ ),
    .Y(\brancher/_0160_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1716_  (.A(\brancher/_0159_ ),
    .B(\brancher/_0160_ ),
    .Y(\brancher/_0161_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1717_  (.A(\brancher/_0121_ ),
    .Y(\brancher/_0162_ ));
 sky130_fd_sc_hd__nand3b_1 \brancher/_1718_  (.A_N(net339),
    .B(\brancher/_0162_ ),
    .C(net341),
    .Y(\brancher/_0163_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1719_  (.A1(\brancher/_0118_ ),
    .A2(\brancher/_0121_ ),
    .B1(net339),
    .Y(\brancher/_0164_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1720_  (.A(\brancher/_0163_ ),
    .B(\brancher/_0164_ ),
    .Y(\brancher/_0165_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1721_  (.A1(\brancher/_0165_ ),
    .A2(\brancher/_0941_ ),
    .B1(\brancher/_0829_ ),
    .Y(\brancher/_0166_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1722_  (.A1(\brancher/_0941_ ),
    .A2(\brancher/_0161_ ),
    .B1(\brancher/_0166_ ),
    .Y(\brancher/_0167_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1723_  (.A(\brancher/rAlu_result[25] ),
    .B(\brancher/_0438_ ),
    .X(\brancher/_0168_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1724_  (.A(\brancher/_0147_ ),
    .B(\brancher/_0167_ ),
    .C(\brancher/_0168_ ),
    .Y(\brancher/_0169_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1725_  (.A(\brancher/_0169_ ),
    .Y(\wPcNextCond[25] ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1726_  (.A(net934),
    .B(net956),
    .Y(\brancher/_0170_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1727_  (.A(net934),
    .B(net956),
    .Y(\brancher/_0171_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1728_  (.A(\brancher/_0171_ ),
    .Y(\brancher/_0172_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1729_  (.A(\brancher/_0170_ ),
    .B(\brancher/_0172_ ),
    .Y(\brancher/_0173_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1730_  (.A(\brancher/_0160_ ),
    .B(\brancher/_0149_ ),
    .Y(\brancher/_0174_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1731_  (.A(\brancher/_0173_ ),
    .B(\brancher/_0174_ ),
    .X(\brancher/_0175_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1732_  (.A(\brancher/_0174_ ),
    .B(\brancher/_0173_ ),
    .Y(\brancher/_0176_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1733_  (.A(\brancher/_0175_ ),
    .B(\brancher/_0430_ ),
    .C(\brancher/_0176_ ),
    .Y(\brancher/_0177_ ));
 sky130_fd_sc_hd__and4_1 \brancher/_1734_  (.A(\brancher/_0956_ ),
    .B(net341),
    .C(net339),
    .D(\brancher/_0120_ ),
    .X(\brancher/_0178_ ));
 sky130_fd_sc_hd__and2_1 \brancher/_1735_  (.A(\brancher/_0873_ ),
    .B(\brancher/_0178_ ),
    .X(\brancher/_0179_ ));
 sky130_fd_sc_hd__xor2_1 \brancher/_1736_  (.A(net336),
    .B(\brancher/_0179_ ),
    .X(\brancher/_0180_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1737_  (.A1(\brancher/_0180_ ),
    .A2(\brancher/_0432_ ),
    .B1(net946),
    .Y(\brancher/_0181_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1738_  (.A(\brancher/_0177_ ),
    .B(\brancher/_0181_ ),
    .Y(\brancher/_0182_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1739_  (.A1(\brancher/rAlu_result[26] ),
    .A2(\brancher/_0096_ ),
    .B1(\brancher/_0588_ ),
    .X(\brancher/_0183_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1740_  (.A(\brancher/_0182_ ),
    .B(\brancher/_0183_ ),
    .Y(\brancher/_0184_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1741_  (.A(net951),
    .B(net956),
    .Y(\brancher/_0185_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1742_  (.A(net951),
    .B(net956),
    .Y(\brancher/_0186_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1743_  (.A(\brancher/_0186_ ),
    .Y(\brancher/_0187_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1744_  (.A(\brancher/_0185_ ),
    .B(\brancher/_0187_ ),
    .Y(\brancher/_0188_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1745_  (.A(\brancher/_0146_ ),
    .B(\brancher/_0136_ ),
    .Y(\brancher/_0189_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1746_  (.A(\brancher/_0188_ ),
    .B(\brancher/_0189_ ),
    .X(\brancher/_0190_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1747_  (.A(\brancher/_0189_ ),
    .B(\brancher/_0188_ ),
    .Y(\brancher/_0191_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1748_  (.A(\brancher/_0190_ ),
    .B(net939),
    .C(\brancher/_0191_ ),
    .Y(\brancher/_0192_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1749_  (.A(\brancher/_0184_ ),
    .B(\brancher/_0192_ ),
    .Y(\wPcNextCond[26] ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1750_  (.A(net951),
    .B(net955),
    .Y(\brancher/_0193_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1751_  (.A(net951),
    .B(net955),
    .Y(\brancher/_0194_ ));
 sky130_fd_sc_hd__and2b_1 \brancher/_1752_  (.A_N(\brancher/_0193_ ),
    .B(\brancher/_0194_ ),
    .X(\brancher/_0195_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1753_  (.A(\brancher/_0138_ ),
    .B(\brancher/_0188_ ),
    .Y(\brancher/_0196_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1754_  (.A(\brancher/_0196_ ),
    .Y(\brancher/_0197_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1755_  (.A(\brancher/_0144_ ),
    .B(\brancher/_0197_ ),
    .Y(\brancher/_0198_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1756_  (.A(\brancher/_0137_ ),
    .B(\brancher/_0187_ ),
    .Y(\brancher/_0199_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1757_  (.A(\brancher/_0198_ ),
    .B(\brancher/_0199_ ),
    .Y(\brancher/_0200_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1758_  (.A(\brancher/_0195_ ),
    .B(\brancher/_0200_ ),
    .X(\brancher/_0201_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1759_  (.A(\brancher/_0200_ ),
    .B(\brancher/_0195_ ),
    .Y(\brancher/_0202_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1760_  (.A(\brancher/_0201_ ),
    .B(\brancher/_0202_ ),
    .Y(\brancher/_0203_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1761_  (.A(\brancher/_0179_ ),
    .B(net336),
    .Y(\brancher/_0204_ ));
 sky130_fd_sc_hd__xnor2_1 \brancher/_1762_  (.A(net335),
    .B(\brancher/_0204_ ),
    .Y(\brancher/_0205_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1763_  (.A1(\brancher/_0205_ ),
    .A2(\brancher/_0941_ ),
    .B1(net946),
    .Y(\brancher/_0206_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1764_  (.A(net935),
    .B(\brancher/rPc_current_reg3[27] ),
    .Y(\brancher/_0207_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1765_  (.A(net935),
    .B(net955),
    .Y(\brancher/_0208_ ));
 sky130_fd_sc_hd__and2b_1 \brancher/_1766_  (.A_N(\brancher/_0207_ ),
    .B(\brancher/_0208_ ),
    .X(\brancher/_0209_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1767_  (.A(\brancher/_0151_ ),
    .B(\brancher/_0173_ ),
    .Y(\brancher/_0210_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1768_  (.A(\brancher/_0210_ ),
    .Y(\brancher/_0211_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1769_  (.A(\brancher/_0158_ ),
    .B(\brancher/_0211_ ),
    .Y(\brancher/_0212_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1770_  (.A(\brancher/_0150_ ),
    .B(\brancher/_0172_ ),
    .Y(\brancher/_0213_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1771_  (.A(\brancher/_0212_ ),
    .B(\brancher/_0213_ ),
    .Y(\brancher/_0214_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1772_  (.A(\brancher/_0209_ ),
    .B(\brancher/_0214_ ),
    .X(\brancher/_0215_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1773_  (.A(\brancher/_0214_ ),
    .B(\brancher/_0209_ ),
    .Y(\brancher/_0216_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1774_  (.A(\brancher/_0215_ ),
    .B(\brancher/_0780_ ),
    .C(\brancher/_0216_ ),
    .Y(\brancher/_0217_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1775_  (.A(\brancher/_0206_ ),
    .B(\brancher/_0217_ ),
    .Y(\brancher/_0218_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1776_  (.A1(\brancher/rAlu_result[27] ),
    .A2(\brancher/_0587_ ),
    .B1(\brancher/_0445_ ),
    .X(\brancher/_0219_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1777_  (.A(\brancher/_0218_ ),
    .B(\brancher/_0219_ ),
    .Y(\brancher/_0220_ ));
 sky130_fd_sc_hd__o21ai_1 \brancher/_1778_  (.A1(\brancher/_0459_ ),
    .A2(\brancher/_0203_ ),
    .B1(\brancher/_0220_ ),
    .Y(\wPcNextCond[27] ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1779_  (.A(\brancher/_0216_ ),
    .B(\brancher/_0208_ ),
    .Y(\brancher/_0221_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1780_  (.A(net935),
    .B(net954),
    .Y(\brancher/_0222_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1781_  (.A(net935),
    .B(net954),
    .Y(\brancher/_0223_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1782_  (.A(\brancher/_0223_ ),
    .Y(\brancher/_0224_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1783_  (.A(\brancher/_0222_ ),
    .B(\brancher/_0224_ ),
    .Y(\brancher/_0225_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1784_  (.A(\brancher/_0221_ ),
    .B(\brancher/_0225_ ),
    .Y(\brancher/_0226_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1785_  (.A(\brancher/_0225_ ),
    .Y(\brancher/_0227_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1786_  (.A(\brancher/_0216_ ),
    .B(\brancher/_0208_ ),
    .C(\brancher/_0227_ ),
    .Y(\brancher/_0228_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1787_  (.A(\brancher/_0226_ ),
    .B(\brancher/_0780_ ),
    .C(\brancher/_0228_ ),
    .Y(\brancher/_0229_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1788_  (.A(net333),
    .Y(\brancher/_0230_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1789_  (.A(net337),
    .B(net335),
    .Y(\brancher/_0231_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1790_  (.A(\brancher/_0231_ ),
    .Y(\brancher/_0232_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1791_  (.A(\brancher/_0873_ ),
    .B(\brancher/_0178_ ),
    .C(\brancher/_0232_ ),
    .Y(\brancher/_0233_ ));
 sky130_fd_sc_hd__xor2_1 \brancher/_1792_  (.A(\brancher/_0230_ ),
    .B(\brancher/_0233_ ),
    .X(\brancher/_0234_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1793_  (.A1(\brancher/_0234_ ),
    .A2(\brancher/_0432_ ),
    .B1(net946),
    .Y(\brancher/_0235_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1794_  (.A(\brancher/_0229_ ),
    .B(\brancher/_0235_ ),
    .Y(\brancher/_0236_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1795_  (.A1(\brancher/rAlu_result[28] ),
    .A2(\brancher/_0096_ ),
    .B1(\brancher/_0588_ ),
    .X(\brancher/_0237_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1796_  (.A(\brancher/_0236_ ),
    .B(\brancher/_0237_ ),
    .Y(\brancher/_0238_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1797_  (.A(\brancher/_0202_ ),
    .B(\brancher/_0194_ ),
    .Y(\brancher/_0239_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1798_  (.A(net951),
    .B(net954),
    .Y(\brancher/_0240_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1799_  (.A(net951),
    .B(\brancher/rPc_current_reg3[28] ),
    .Y(\brancher/_0241_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1800_  (.A(\brancher/_0241_ ),
    .Y(\brancher/_0242_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1801_  (.A(\brancher/_0240_ ),
    .B(\brancher/_0242_ ),
    .Y(\brancher/_0243_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1802_  (.A(\brancher/_0239_ ),
    .B(\brancher/_0243_ ),
    .Y(\brancher/_0244_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1803_  (.A(\brancher/_0243_ ),
    .Y(\brancher/_0245_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1804_  (.A(\brancher/_0202_ ),
    .B(\brancher/_0194_ ),
    .C(\brancher/_0245_ ),
    .Y(\brancher/_0246_ ));
 sky130_fd_sc_hd__nand3_2 \brancher/_1805_  (.A(\brancher/_0244_ ),
    .B(net940),
    .C(\brancher/_0246_ ),
    .Y(\brancher/_0247_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1806_  (.A(\brancher/_0238_ ),
    .B(\brancher/_0247_ ),
    .Y(\wPcNextCond[28] ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1807_  (.A(\brancher/_0230_ ),
    .B(\brancher/_0233_ ),
    .Y(\brancher/_0248_ ));
 sky130_fd_sc_hd__xor2_1 \brancher/_1808_  (.A(net332),
    .B(\brancher/_0248_ ),
    .X(\brancher/_0249_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1809_  (.A1(\brancher/_0249_ ),
    .A2(\brancher/_0941_ ),
    .B1(\brancher/_0829_ ),
    .Y(\brancher/_0250_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1810_  (.A(net936),
    .B(\brancher/rPc_current_reg3[29] ),
    .Y(\brancher/_0251_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1811_  (.A(net935),
    .B(\brancher/rPc_current_reg3[29] ),
    .Y(\brancher/_0252_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1812_  (.A(\brancher/_0252_ ),
    .Y(\brancher/_0253_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1813_  (.A(\brancher/_0251_ ),
    .B(\brancher/_0253_ ),
    .Y(\brancher/_0254_ ));
 sky130_fd_sc_hd__and3_1 \brancher/_1814_  (.A(\brancher/_0211_ ),
    .B(\brancher/_0209_ ),
    .C(\brancher/_0225_ ),
    .X(\brancher/_0255_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1815_  (.A(\brancher/_0158_ ),
    .B(\brancher/_0255_ ),
    .Y(\brancher/_0256_ ));
 sky130_fd_sc_hd__o41a_1 \brancher/_1816_  (.A1(net957),
    .A2(net956),
    .A3(net955),
    .A4(net954),
    .B1(net935),
    .X(\brancher/_0257_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1817_  (.A(\brancher/_0257_ ),
    .Y(\brancher/_0258_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1818_  (.A(\brancher/_0256_ ),
    .B(\brancher/_0258_ ),
    .Y(\brancher/_0259_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1819_  (.A(\brancher/_0254_ ),
    .B(\brancher/_0259_ ),
    .X(\brancher/_0260_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1820_  (.A(\brancher/_0259_ ),
    .B(\brancher/_0254_ ),
    .Y(\brancher/_0261_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1821_  (.A(\brancher/_0260_ ),
    .B(\brancher/_0430_ ),
    .C(\brancher/_0261_ ),
    .Y(\brancher/_0262_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1822_  (.A(\brancher/_0250_ ),
    .B(\brancher/_0262_ ),
    .Y(\brancher/_0263_ ));
 sky130_fd_sc_hd__and3_1 \brancher/_1823_  (.A(\brancher/_0197_ ),
    .B(\brancher/_0195_ ),
    .C(\brancher/_0243_ ),
    .X(\brancher/_0264_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1824_  (.A(\brancher/_0144_ ),
    .B(\brancher/_0264_ ),
    .Y(\brancher/_0265_ ));
 sky130_fd_sc_hd__o41a_1 \brancher/_1825_  (.A1(\brancher/rPc_current_reg3[25] ),
    .A2(\brancher/rPc_current_reg3[26] ),
    .A3(net955),
    .A4(net954),
    .B1(net952),
    .X(\brancher/_0266_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1826_  (.A(\brancher/_0266_ ),
    .Y(\brancher/_0267_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1827_  (.A(\brancher/_0265_ ),
    .B(\brancher/_0267_ ),
    .Y(\brancher/_0268_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1828_  (.A(net952),
    .B(\brancher/rPc_current_reg3[29] ),
    .Y(\brancher/_0269_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1829_  (.A(net952),
    .B(\brancher/rPc_current_reg3[29] ),
    .Y(\brancher/_0270_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1830_  (.A(\brancher/_0270_ ),
    .Y(\brancher/_0271_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1831_  (.A(\brancher/_0269_ ),
    .B(\brancher/_0271_ ),
    .Y(\brancher/_0272_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1832_  (.A(\brancher/_0272_ ),
    .Y(\brancher/_0273_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1833_  (.A(\brancher/_0268_ ),
    .B(\brancher/_0273_ ),
    .Y(\brancher/_0274_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1834_  (.A(\brancher/_0265_ ),
    .B(\brancher/_0267_ ),
    .C(\brancher/_0272_ ),
    .Y(\brancher/_0275_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1835_  (.A(\brancher/_0274_ ),
    .B(net940),
    .C(\brancher/_0275_ ),
    .Y(\brancher/_0276_ ));
 sky130_fd_sc_hd__or2_1 \brancher/_1836_  (.A(\brancher/rAlu_result[29] ),
    .B(\brancher/_0438_ ),
    .X(\brancher/_0277_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1837_  (.A(\brancher/_0263_ ),
    .B(\brancher/_0276_ ),
    .C(\brancher/_0277_ ),
    .Y(\brancher/_0278_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1838_  (.A(\brancher/_0278_ ),
    .Y(\wPcNextCond[29] ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1839_  (.A(\brancher/_0261_ ),
    .B(\brancher/_0252_ ),
    .Y(\brancher/_0279_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1840_  (.A(net936),
    .B(\brancher/rPc_current_reg3[30] ),
    .Y(\brancher/_0280_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1841_  (.A(net936),
    .B(\brancher/rPc_current_reg3[30] ),
    .Y(\brancher/_0281_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1842_  (.A(\brancher/_0281_ ),
    .Y(\brancher/_0282_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1843_  (.A(\brancher/_0280_ ),
    .B(\brancher/_0282_ ),
    .Y(\brancher/_0283_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1844_  (.A(\brancher/_0279_ ),
    .B(\brancher/_0283_ ),
    .Y(\brancher/_0284_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1845_  (.A(\brancher/_0283_ ),
    .Y(\brancher/_0285_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1846_  (.A(\brancher/_0261_ ),
    .B(\brancher/_0252_ ),
    .C(\brancher/_0285_ ),
    .Y(\brancher/_0286_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1847_  (.A(\brancher/_0284_ ),
    .B(\brancher/_0780_ ),
    .C(\brancher/_0286_ ),
    .Y(\brancher/_0287_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1848_  (.A(net330),
    .Y(\brancher/_0288_ ));
 sky130_fd_sc_hd__and3_1 \brancher/_1849_  (.A(\brancher/_0232_ ),
    .B(net333),
    .C(net332),
    .X(\brancher/_0289_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1850_  (.A(\brancher/_0873_ ),
    .B(\brancher/_0178_ ),
    .C(\brancher/_0289_ ),
    .Y(\brancher/_0290_ ));
 sky130_fd_sc_hd__xor2_1 \brancher/_1851_  (.A(\brancher/_0288_ ),
    .B(\brancher/_0290_ ),
    .X(\brancher/_0291_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1852_  (.A1(\brancher/_0291_ ),
    .A2(\brancher/_0432_ ),
    .B1(\brancher/rOp_jalr ),
    .Y(\brancher/_0292_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1853_  (.A(\brancher/_0287_ ),
    .B(\brancher/_0292_ ),
    .Y(\brancher/_0293_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1854_  (.A1(\brancher/rAlu_result[30] ),
    .A2(\brancher/_0096_ ),
    .B1(\brancher/_0588_ ),
    .X(\brancher/_0294_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1855_  (.A(\brancher/_0293_ ),
    .B(\brancher/_0294_ ),
    .Y(\brancher/_0295_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1856_  (.A(\brancher/_0268_ ),
    .B(\brancher/_0272_ ),
    .Y(\brancher/_0296_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1857_  (.A(\brancher/_0296_ ),
    .B(\brancher/_0270_ ),
    .Y(\brancher/_0297_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1858_  (.A(net952),
    .B(\brancher/rPc_current_reg3[30] ),
    .Y(\brancher/_0298_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1859_  (.A(net952),
    .B(\brancher/rPc_current_reg3[30] ),
    .Y(\brancher/_0299_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1860_  (.A(\brancher/_0299_ ),
    .Y(\brancher/_0300_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1861_  (.A(\brancher/_0298_ ),
    .B(\brancher/_0300_ ),
    .Y(\brancher/_0301_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1862_  (.A(\brancher/_0297_ ),
    .B(\brancher/_0301_ ),
    .Y(\brancher/_0302_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1863_  (.A(\brancher/_0301_ ),
    .Y(\brancher/_0303_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1864_  (.A(\brancher/_0296_ ),
    .B(\brancher/_0270_ ),
    .C(\brancher/_0303_ ),
    .Y(\brancher/_0304_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1865_  (.A(\brancher/_0302_ ),
    .B(net940),
    .C(\brancher/_0304_ ),
    .Y(\brancher/_0305_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1866_  (.A(\brancher/_0295_ ),
    .B(\brancher/_0305_ ),
    .Y(\wPcNextCond[30] ));
 sky130_fd_sc_hd__and2_1 \brancher/_1867_  (.A(\brancher/_0254_ ),
    .B(\brancher/_0283_ ),
    .X(\brancher/_0306_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1868_  (.A(\brancher/_0259_ ),
    .B(\brancher/_0306_ ),
    .Y(\brancher/_0307_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1869_  (.A(\brancher/_0253_ ),
    .B(\brancher/_0282_ ),
    .Y(\brancher/_0308_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1870_  (.A(\brancher/_0307_ ),
    .B(\brancher/_0308_ ),
    .Y(\brancher/_0309_ ));
 sky130_fd_sc_hd__xnor2_1 \brancher/_1871_  (.A(net938),
    .B(\brancher/rPc_current_reg3[31] ),
    .Y(\brancher/_0310_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1872_  (.A(\brancher/_0310_ ),
    .Y(\brancher/_0311_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1873_  (.A(\brancher/_0309_ ),
    .B(\brancher/_0311_ ),
    .Y(\brancher/_0312_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1874_  (.A(\brancher/_0307_ ),
    .B(\brancher/_0308_ ),
    .C(\brancher/_0310_ ),
    .Y(\brancher/_0313_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1875_  (.A(\brancher/_0312_ ),
    .B(\brancher/_0780_ ),
    .C(\brancher/_0313_ ),
    .Y(\brancher/_0314_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1876_  (.A(\brancher/_0288_ ),
    .B(\brancher/_0290_ ),
    .Y(\brancher/_0315_ ));
 sky130_fd_sc_hd__xor2_1 \brancher/_1877_  (.A(net329),
    .B(\brancher/_0315_ ),
    .X(\brancher/_0316_ ));
 sky130_fd_sc_hd__a21oi_1 \brancher/_1878_  (.A1(\brancher/_0316_ ),
    .A2(\brancher/_0432_ ),
    .B1(net947),
    .Y(\brancher/_0317_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1879_  (.A(\brancher/_0314_ ),
    .B(\brancher/_0317_ ),
    .Y(\brancher/_0318_ ));
 sky130_fd_sc_hd__o21a_1 \brancher/_1880_  (.A1(\brancher/rAlu_result[31] ),
    .A2(\brancher/_0096_ ),
    .B1(\brancher/_0588_ ),
    .X(\brancher/_0319_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1881_  (.A(\brancher/_0318_ ),
    .B(\brancher/_0319_ ),
    .Y(\brancher/_0320_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1882_  (.A(\brancher/_0273_ ),
    .B(\brancher/_0303_ ),
    .Y(\brancher/_0321_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1883_  (.A(\brancher/_0268_ ),
    .B(\brancher/_0321_ ),
    .Y(\brancher/_0322_ ));
 sky130_fd_sc_hd__nor2_1 \brancher/_1884_  (.A(\brancher/_0271_ ),
    .B(\brancher/_0300_ ),
    .Y(\brancher/_0323_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1885_  (.A(\brancher/_0322_ ),
    .B(\brancher/_0323_ ),
    .Y(\brancher/_0324_ ));
 sky130_fd_sc_hd__xnor2_1 \brancher/_1886_  (.A(net952),
    .B(\brancher/rPc_current_reg3[31] ),
    .Y(\brancher/_0325_ ));
 sky130_fd_sc_hd__inv_2 \brancher/_1887_  (.A(\brancher/_0325_ ),
    .Y(\brancher/_0326_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1888_  (.A(\brancher/_0324_ ),
    .B(\brancher/_0326_ ),
    .Y(\brancher/_0327_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1889_  (.A(\brancher/_0322_ ),
    .B(\brancher/_0323_ ),
    .C(\brancher/_0325_ ),
    .Y(\brancher/_0328_ ));
 sky130_fd_sc_hd__nand3_1 \brancher/_1890_  (.A(\brancher/_0327_ ),
    .B(net940),
    .C(\brancher/_0328_ ),
    .Y(\brancher/_0329_ ));
 sky130_fd_sc_hd__nand2_1 \brancher/_1891_  (.A(\brancher/_0320_ ),
    .B(\brancher/_0329_ ),
    .Y(\wPcNextCond[31] ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1892_  (.A0(net2138),
    .A1(\brancher/rPc_current_reg3[0] ),
    .S(net274),
    .X(\brancher/_0330_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1893_  (.A(\brancher/_0330_ ),
    .X(\brancher/_0000_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1894_  (.A0(net2147),
    .A1(\brancher/rPc_current_reg3[1] ),
    .S(net274),
    .X(\brancher/_0331_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1895_  (.A(\brancher/_0331_ ),
    .X(\brancher/_0001_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1896_  (.A0(net2132),
    .A1(\brancher/rPc_current_reg3[2] ),
    .S(net272),
    .X(\brancher/_0332_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1897_  (.A(\brancher/_0332_ ),
    .X(\brancher/_0002_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1898_  (.A0(net2149),
    .A1(\brancher/rPc_current_reg3[3] ),
    .S(net269),
    .X(\brancher/_0333_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1899_  (.A(\brancher/_0333_ ),
    .X(\brancher/_0003_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1900_  (.A0(net2121),
    .A1(\brancher/rPc_current_reg3[4] ),
    .S(net269),
    .X(\brancher/_0334_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1901_  (.A(\brancher/_0334_ ),
    .X(\brancher/_0004_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1902_  (.A0(net2118),
    .A1(\brancher/rPc_current_reg3[5] ),
    .S(net268),
    .X(\brancher/_0335_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1903_  (.A(\brancher/_0335_ ),
    .X(\brancher/_0005_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1904_  (.A0(net2113),
    .A1(\brancher/rPc_current_reg3[6] ),
    .S(net266),
    .X(\brancher/_0336_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1905_  (.A(\brancher/_0336_ ),
    .X(\brancher/_0006_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1906_  (.A0(net2095),
    .A1(\brancher/rPc_current_reg3[7] ),
    .S(net276),
    .X(\brancher/_0337_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1907_  (.A(\brancher/_0337_ ),
    .X(\brancher/_0007_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1908_  (.A0(net2112),
    .A1(\brancher/rPc_current_reg3[8] ),
    .S(net271),
    .X(\brancher/_0338_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1909_  (.A(\brancher/_0338_ ),
    .X(\brancher/_0008_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1910_  (.A0(\brancher/rPc_current_reg2[9] ),
    .A1(\brancher/rPc_current_reg3[9] ),
    .S(net264),
    .X(\brancher/_0339_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1911_  (.A(\brancher/_0339_ ),
    .X(\brancher/_0009_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1912_  (.A0(\brancher/rPc_current_reg2[10] ),
    .A1(\brancher/rPc_current_reg3[10] ),
    .S(net263),
    .X(\brancher/_0340_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1913_  (.A(\brancher/_0340_ ),
    .X(\brancher/_0010_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1914_  (.A0(net2120),
    .A1(\brancher/rPc_current_reg3[11] ),
    .S(net263),
    .X(\brancher/_0341_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1915_  (.A(\brancher/_0341_ ),
    .X(\brancher/_0011_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1916_  (.A0(net2099),
    .A1(\brancher/rPc_current_reg3[12] ),
    .S(net239),
    .X(\brancher/_0342_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1917_  (.A(\brancher/_0342_ ),
    .X(\brancher/_0012_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1918_  (.A0(net2083),
    .A1(\brancher/rPc_current_reg3[13] ),
    .S(net241),
    .X(\brancher/_0343_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1919_  (.A(\brancher/_0343_ ),
    .X(\brancher/_0013_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1920_  (.A0(net2043),
    .A1(\brancher/rPc_current_reg3[14] ),
    .S(net239),
    .X(\brancher/_0344_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1921_  (.A(\brancher/_0344_ ),
    .X(\brancher/_0014_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1922_  (.A0(net2115),
    .A1(\brancher/rPc_current_reg3[15] ),
    .S(net249),
    .X(\brancher/_0345_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1923_  (.A(\brancher/_0345_ ),
    .X(\brancher/_0015_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1924_  (.A0(net2087),
    .A1(\brancher/rPc_current_reg3[16] ),
    .S(net239),
    .X(\brancher/_0346_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1925_  (.A(\brancher/_0346_ ),
    .X(\brancher/_0016_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1926_  (.A0(net2050),
    .A1(\brancher/rPc_current_reg3[17] ),
    .S(net258),
    .X(\brancher/_0347_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1927_  (.A(\brancher/_0347_ ),
    .X(\brancher/_0017_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1928_  (.A0(net2037),
    .A1(\brancher/rPc_current_reg3[18] ),
    .S(net259),
    .X(\brancher/_0348_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1929_  (.A(\brancher/_0348_ ),
    .X(\brancher/_0018_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1930_  (.A0(net2064),
    .A1(\brancher/rPc_current_reg3[19] ),
    .S(net251),
    .X(\brancher/_0349_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1931_  (.A(\brancher/_0349_ ),
    .X(\brancher/_0019_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1932_  (.A0(net2081),
    .A1(\brancher/rPc_current_reg3[20] ),
    .S(net251),
    .X(\brancher/_0350_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1933_  (.A(\brancher/_0350_ ),
    .X(\brancher/_0020_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1934_  (.A0(net2055),
    .A1(net958),
    .S(net252),
    .X(\brancher/_0351_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1935_  (.A(\brancher/_0351_ ),
    .X(\brancher/_0021_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1936_  (.A0(net1975),
    .A1(\brancher/rPc_current_reg3[22] ),
    .S(net252),
    .X(\brancher/_0352_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1937_  (.A(\brancher/_0352_ ),
    .X(\brancher/_0022_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1938_  (.A0(net2092),
    .A1(\brancher/rPc_current_reg3[23] ),
    .S(net254),
    .X(\brancher/_0353_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1939_  (.A(\brancher/_0353_ ),
    .X(\brancher/_0023_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1940_  (.A0(net1987),
    .A1(\brancher/rPc_current_reg3[24] ),
    .S(net254),
    .X(\brancher/_0354_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1941_  (.A(\brancher/_0354_ ),
    .X(\brancher/_0024_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1942_  (.A0(net2102),
    .A1(net957),
    .S(net255),
    .X(\brancher/_0355_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1943_  (.A(\brancher/_0355_ ),
    .X(\brancher/_0025_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1944_  (.A0(net2058),
    .A1(net956),
    .S(net254),
    .X(\brancher/_0356_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1945_  (.A(\brancher/_0356_ ),
    .X(\brancher/_0026_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1946_  (.A0(net2105),
    .A1(net955),
    .S(net256),
    .X(\brancher/_0357_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1947_  (.A(\brancher/_0357_ ),
    .X(\brancher/_0027_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1948_  (.A0(net2086),
    .A1(net954),
    .S(net255),
    .X(\brancher/_0358_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1949_  (.A(\brancher/_0358_ ),
    .X(\brancher/_0028_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1950_  (.A0(net2059),
    .A1(\brancher/rPc_current_reg3[29] ),
    .S(net256),
    .X(\brancher/_0359_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1951_  (.A(\brancher/_0359_ ),
    .X(\brancher/_0029_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1952_  (.A0(net2033),
    .A1(\brancher/rPc_current_reg3[30] ),
    .S(net256),
    .X(\brancher/_0360_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1953_  (.A(\brancher/_0360_ ),
    .X(\brancher/_0030_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1954_  (.A0(net2075),
    .A1(\brancher/rPc_current_reg3[31] ),
    .S(net258),
    .X(\brancher/_0361_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1955_  (.A(\brancher/_0361_ ),
    .X(\brancher/_0031_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1956_  (.A0(net135),
    .A1(\brancher/rPc_current_reg1[0] ),
    .S(net275),
    .X(\brancher/_0362_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1957_  (.A(\brancher/_0362_ ),
    .X(\brancher/_0032_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1958_  (.A0(net146),
    .A1(\brancher/rPc_current_reg1[1] ),
    .S(net275),
    .X(\brancher/_0363_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1959_  (.A(\brancher/_0363_ ),
    .X(\brancher/_0033_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1960_  (.A0(net379),
    .A1(\brancher/rPc_current_reg1[2] ),
    .S(net271),
    .X(\brancher/_0364_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1961_  (.A(\brancher/_0364_ ),
    .X(\brancher/_0034_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1962_  (.A0(net377),
    .A1(\brancher/rPc_current_reg1[3] ),
    .S(net275),
    .X(\brancher/_0365_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1963_  (.A(\brancher/_0365_ ),
    .X(\brancher/_0035_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1964_  (.A0(net376),
    .A1(\brancher/rPc_current_reg1[4] ),
    .S(net268),
    .X(\brancher/_0366_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1965_  (.A(\brancher/_0366_ ),
    .X(\brancher/_0036_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1966_  (.A0(net162),
    .A1(\brancher/rPc_current_reg1[5] ),
    .S(net272),
    .X(\brancher/_0367_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1967_  (.A(\brancher/_0367_ ),
    .X(\brancher/_0037_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1968_  (.A0(net374),
    .A1(\brancher/rPc_current_reg1[6] ),
    .S(net266),
    .X(\brancher/_0368_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1969_  (.A(\brancher/_0368_ ),
    .X(\brancher/_0038_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1970_  (.A0(net164),
    .A1(\brancher/rPc_current_reg1[7] ),
    .S(net276),
    .X(\brancher/_0369_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1971_  (.A(\brancher/_0369_ ),
    .X(\brancher/_0039_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1972_  (.A0(net371),
    .A1(\brancher/rPc_current_reg1[8] ),
    .S(net271),
    .X(\brancher/_0370_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1973_  (.A(\brancher/_0370_ ),
    .X(\brancher/_0040_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1974_  (.A0(net370),
    .A1(\brancher/rPc_current_reg1[9] ),
    .S(net271),
    .X(\brancher/_0371_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1975_  (.A(\brancher/_0371_ ),
    .X(\brancher/_0041_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1976_  (.A0(net369),
    .A1(\brancher/rPc_current_reg1[10] ),
    .S(net267),
    .X(\brancher/_0372_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1977_  (.A(\brancher/_0372_ ),
    .X(\brancher/_0042_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1978_  (.A0(net367),
    .A1(\brancher/rPc_current_reg1[11] ),
    .S(net266),
    .X(\brancher/_0373_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1979_  (.A(\brancher/_0373_ ),
    .X(\brancher/_0043_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1980_  (.A0(net363),
    .A1(\brancher/rPc_current_reg1[12] ),
    .S(net239),
    .X(\brancher/_0374_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1981_  (.A(\brancher/_0374_ ),
    .X(\brancher/_0044_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1982_  (.A0(net362),
    .A1(\brancher/rPc_current_reg1[13] ),
    .S(net251),
    .X(\brancher/_0375_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1983_  (.A(\brancher/_0375_ ),
    .X(\brancher/_0045_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1984_  (.A0(net360),
    .A1(\brancher/rPc_current_reg1[14] ),
    .S(net257),
    .X(\brancher/_0376_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1985_  (.A(\brancher/_0376_ ),
    .X(\brancher/_0046_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1986_  (.A0(net357),
    .A1(\brancher/rPc_current_reg1[15] ),
    .S(net253),
    .X(\brancher/_0377_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1987_  (.A(\brancher/_0377_ ),
    .X(\brancher/_0047_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1988_  (.A0(net354),
    .A1(\brancher/rPc_current_reg1[16] ),
    .S(net251),
    .X(\brancher/_0378_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1989_  (.A(\brancher/_0378_ ),
    .X(\brancher/_0048_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1990_  (.A0(net352),
    .A1(\brancher/rPc_current_reg1[17] ),
    .S(net253),
    .X(\brancher/_0379_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1991_  (.A(\brancher/_0379_ ),
    .X(\brancher/_0049_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1992_  (.A0(net350),
    .A1(\brancher/rPc_current_reg1[18] ),
    .S(net258),
    .X(\brancher/_0380_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1993_  (.A(\brancher/_0380_ ),
    .X(\brancher/_0050_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1994_  (.A0(net348),
    .A1(\brancher/rPc_current_reg1[19] ),
    .S(net253),
    .X(\brancher/_0381_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1995_  (.A(\brancher/_0381_ ),
    .X(\brancher/_0051_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1996_  (.A0(net346),
    .A1(\brancher/rPc_current_reg1[20] ),
    .S(net252),
    .X(\brancher/_0382_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1997_  (.A(\brancher/_0382_ ),
    .X(\brancher/_0052_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_1998_  (.A0(net148),
    .A1(\brancher/rPc_current_reg1[21] ),
    .S(net277),
    .X(\brancher/_0383_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_1999_  (.A(\brancher/_0383_ ),
    .X(\brancher/_0053_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2000_  (.A0(net344),
    .A1(\brancher/rPc_current_reg1[22] ),
    .S(net276),
    .X(\brancher/_0384_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2001_  (.A(\brancher/_0384_ ),
    .X(\brancher/_0054_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2002_  (.A0(net150),
    .A1(\brancher/rPc_current_reg1[23] ),
    .S(net276),
    .X(\brancher/_0385_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2003_  (.A(\brancher/_0385_ ),
    .X(\brancher/_0055_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2004_  (.A0(net341),
    .A1(\brancher/rPc_current_reg1[24] ),
    .S(net275),
    .X(\brancher/_0386_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2005_  (.A(\brancher/_0386_ ),
    .X(\brancher/_0056_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2006_  (.A0(net152),
    .A1(\brancher/rPc_current_reg1[25] ),
    .S(net277),
    .X(\brancher/_0387_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2007_  (.A(\brancher/_0387_ ),
    .X(\brancher/_0057_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2008_  (.A0(net338),
    .A1(\brancher/rPc_current_reg1[26] ),
    .S(net274),
    .X(\brancher/_0388_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2009_  (.A(\brancher/_0388_ ),
    .X(\brancher/_0058_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2010_  (.A0(net154),
    .A1(\brancher/rPc_current_reg1[27] ),
    .S(net274),
    .X(\brancher/_0389_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2011_  (.A(\brancher/_0389_ ),
    .X(\brancher/_0059_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2012_  (.A0(net334),
    .A1(\brancher/rPc_current_reg1[28] ),
    .S(net277),
    .X(\brancher/_0390_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2013_  (.A(\brancher/_0390_ ),
    .X(\brancher/_0060_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2014_  (.A0(net156),
    .A1(\brancher/rPc_current_reg1[29] ),
    .S(net274),
    .X(\brancher/_0391_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2015_  (.A(\brancher/_0391_ ),
    .X(\brancher/_0061_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2016_  (.A0(net331),
    .A1(\brancher/rPc_current_reg1[30] ),
    .S(net277),
    .X(\brancher/_0392_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2017_  (.A(\brancher/_0392_ ),
    .X(\brancher/_0062_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2018_  (.A0(net329),
    .A1(\brancher/rPc_current_reg1[31] ),
    .S(net277),
    .X(\brancher/_0393_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2019_  (.A(\brancher/_0393_ ),
    .X(\brancher/_0063_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2020_  (.A0(\brancher/rPc_current_reg1[0] ),
    .A1(net2138),
    .S(net274),
    .X(\brancher/_0394_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2021_  (.A(\brancher/_0394_ ),
    .X(\brancher/_0064_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2022_  (.A0(\brancher/rPc_current_reg1[1] ),
    .A1(net2147),
    .S(net275),
    .X(\brancher/_0395_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2023_  (.A(\brancher/_0395_ ),
    .X(\brancher/_0065_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2024_  (.A0(\brancher/rPc_current_reg1[2] ),
    .A1(net2132),
    .S(net272),
    .X(\brancher/_0396_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2025_  (.A(\brancher/_0396_ ),
    .X(\brancher/_0066_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2026_  (.A0(\brancher/rPc_current_reg1[3] ),
    .A1(net2149),
    .S(net269),
    .X(\brancher/_0397_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2027_  (.A(\brancher/_0397_ ),
    .X(\brancher/_0067_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2028_  (.A0(\brancher/rPc_current_reg1[4] ),
    .A1(net2121),
    .S(net269),
    .X(\brancher/_0398_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2029_  (.A(\brancher/_0398_ ),
    .X(\brancher/_0068_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2030_  (.A0(\brancher/rPc_current_reg1[5] ),
    .A1(net2118),
    .S(net266),
    .X(\brancher/_0399_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2031_  (.A(\brancher/_0399_ ),
    .X(\brancher/_0069_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2032_  (.A0(\brancher/rPc_current_reg1[6] ),
    .A1(net2113),
    .S(net267),
    .X(\brancher/_0400_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2033_  (.A(\brancher/_0400_ ),
    .X(\brancher/_0070_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2034_  (.A0(\brancher/rPc_current_reg1[7] ),
    .A1(net2095),
    .S(net276),
    .X(\brancher/_0401_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2035_  (.A(\brancher/_0401_ ),
    .X(\brancher/_0071_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2036_  (.A0(\brancher/rPc_current_reg1[8] ),
    .A1(net2112),
    .S(net271),
    .X(\brancher/_0402_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2037_  (.A(\brancher/_0402_ ),
    .X(\brancher/_0072_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2038_  (.A0(\brancher/rPc_current_reg1[9] ),
    .A1(\brancher/rPc_current_reg2[9] ),
    .S(net271),
    .X(\brancher/_0403_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2039_  (.A(\brancher/_0403_ ),
    .X(\brancher/_0073_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2040_  (.A0(\brancher/rPc_current_reg1[10] ),
    .A1(\brancher/rPc_current_reg2[10] ),
    .S(net267),
    .X(\brancher/_0404_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2041_  (.A(\brancher/_0404_ ),
    .X(\brancher/_0074_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2042_  (.A0(\brancher/rPc_current_reg1[11] ),
    .A1(net2120),
    .S(net263),
    .X(\brancher/_0405_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2043_  (.A(\brancher/_0405_ ),
    .X(\brancher/_0075_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2044_  (.A0(\brancher/rPc_current_reg1[12] ),
    .A1(net2099),
    .S(net239),
    .X(\brancher/_0406_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2045_  (.A(\brancher/_0406_ ),
    .X(\brancher/_0076_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2046_  (.A0(\brancher/rPc_current_reg1[13] ),
    .A1(net2083),
    .S(net251),
    .X(\brancher/_0407_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2047_  (.A(\brancher/_0407_ ),
    .X(\brancher/_0077_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2048_  (.A0(\brancher/rPc_current_reg1[14] ),
    .A1(net2043),
    .S(net257),
    .X(\brancher/_0408_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2049_  (.A(\brancher/_0408_ ),
    .X(\brancher/_0078_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2050_  (.A0(\brancher/rPc_current_reg1[15] ),
    .A1(net2115),
    .S(net240),
    .X(\brancher/_0409_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2051_  (.A(\brancher/_0409_ ),
    .X(\brancher/_0079_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2052_  (.A0(\brancher/rPc_current_reg1[16] ),
    .A1(net2087),
    .S(net241),
    .X(\brancher/_0410_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2053_  (.A(\brancher/_0410_ ),
    .X(\brancher/_0080_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2054_  (.A0(\brancher/rPc_current_reg1[17] ),
    .A1(net2050),
    .S(net253),
    .X(\brancher/_0411_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2055_  (.A(\brancher/_0411_ ),
    .X(\brancher/_0081_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2056_  (.A0(\brancher/rPc_current_reg1[18] ),
    .A1(net2037),
    .S(net258),
    .X(\brancher/_0412_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2057_  (.A(\brancher/_0412_ ),
    .X(\brancher/_0082_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2058_  (.A0(\brancher/rPc_current_reg1[19] ),
    .A1(net2064),
    .S(net252),
    .X(\brancher/_0413_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2059_  (.A(\brancher/_0413_ ),
    .X(\brancher/_0083_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2060_  (.A0(\brancher/rPc_current_reg1[20] ),
    .A1(net2081),
    .S(net252),
    .X(\brancher/_0414_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2061_  (.A(\brancher/_0414_ ),
    .X(\brancher/_0084_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2062_  (.A0(\brancher/rPc_current_reg1[21] ),
    .A1(net2055),
    .S(net252),
    .X(\brancher/_0415_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2063_  (.A(\brancher/_0415_ ),
    .X(\brancher/_0085_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2064_  (.A0(\brancher/rPc_current_reg1[22] ),
    .A1(net1975),
    .S(net254),
    .X(\brancher/_0416_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2065_  (.A(\brancher/_0416_ ),
    .X(\brancher/_0086_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2066_  (.A0(\brancher/rPc_current_reg1[23] ),
    .A1(net2092),
    .S(net255),
    .X(\brancher/_0417_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2067_  (.A(\brancher/_0417_ ),
    .X(\brancher/_0087_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2068_  (.A0(\brancher/rPc_current_reg1[24] ),
    .A1(net1987),
    .S(net254),
    .X(\brancher/_0418_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2069_  (.A(\brancher/_0418_ ),
    .X(\brancher/_0088_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2070_  (.A0(\brancher/rPc_current_reg1[25] ),
    .A1(net2102),
    .S(net256),
    .X(\brancher/_0419_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2071_  (.A(\brancher/_0419_ ),
    .X(\brancher/_0089_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2072_  (.A0(\brancher/rPc_current_reg1[26] ),
    .A1(net2058),
    .S(net254),
    .X(\brancher/_0420_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2073_  (.A(\brancher/_0420_ ),
    .X(\brancher/_0090_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2074_  (.A0(\brancher/rPc_current_reg1[27] ),
    .A1(net2105),
    .S(net255),
    .X(\brancher/_0421_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2075_  (.A(\brancher/_0421_ ),
    .X(\brancher/_0091_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2076_  (.A0(\brancher/rPc_current_reg1[28] ),
    .A1(net2086),
    .S(net255),
    .X(\brancher/_0422_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2077_  (.A(\brancher/_0422_ ),
    .X(\brancher/_0092_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2078_  (.A0(\brancher/rPc_current_reg1[29] ),
    .A1(net2059),
    .S(net256),
    .X(\brancher/_0423_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2079_  (.A(\brancher/_0423_ ),
    .X(\brancher/_0093_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2080_  (.A0(\brancher/rPc_current_reg1[30] ),
    .A1(net2033),
    .S(net257),
    .X(\brancher/_0424_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2081_  (.A(\brancher/_0424_ ),
    .X(\brancher/_0094_ ));
 sky130_fd_sc_hd__mux2_1 \brancher/_2082_  (.A0(\brancher/rPc_current_reg1[31] ),
    .A1(net2075),
    .S(net258),
    .X(\brancher/_0425_ ));
 sky130_fd_sc_hd__clkbuf_1 \brancher/_2083_  (.A(\brancher/_0425_ ),
    .X(\brancher/_0095_ ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2084_  (.CLK(clknet_leaf_53_clk),
    .D(\brancher/_0000_ ),
    .Q(\brancher/rPc_current_reg3[0] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2085_  (.CLK(clknet_leaf_53_clk),
    .D(\brancher/_0001_ ),
    .Q(\brancher/rPc_current_reg3[1] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2086_  (.CLK(clknet_leaf_56_clk),
    .D(\brancher/_0002_ ),
    .Q(\brancher/rPc_current_reg3[2] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2087_  (.CLK(clknet_leaf_62_clk),
    .D(\brancher/_0003_ ),
    .Q(\brancher/rPc_current_reg3[3] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2088_  (.CLK(clknet_leaf_62_clk),
    .D(\brancher/_0004_ ),
    .Q(\brancher/rPc_current_reg3[4] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2089_  (.CLK(clknet_leaf_57_clk),
    .D(\brancher/_0005_ ),
    .Q(\brancher/rPc_current_reg3[5] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2090_  (.CLK(clknet_leaf_57_clk),
    .D(\brancher/_0006_ ),
    .Q(\brancher/rPc_current_reg3[6] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2091_  (.CLK(clknet_leaf_52_clk),
    .D(\brancher/_0007_ ),
    .Q(\brancher/rPc_current_reg3[7] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2092_  (.CLK(clknet_leaf_57_clk),
    .D(\brancher/_0008_ ),
    .Q(\brancher/rPc_current_reg3[8] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2093_  (.CLK(clknet_leaf_62_clk),
    .D(\brancher/_0009_ ),
    .Q(\brancher/rPc_current_reg3[9] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2094_  (.CLK(clknet_leaf_63_clk),
    .D(\brancher/_0010_ ),
    .Q(\brancher/rPc_current_reg3[10] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2095_  (.CLK(clknet_leaf_63_clk),
    .D(\brancher/_0011_ ),
    .Q(\brancher/rPc_current_reg3[11] ));
 sky130_fd_sc_hd__dfxtp_2 \brancher/_2096_  (.CLK(clknet_leaf_25_clk),
    .D(\brancher/_0012_ ),
    .Q(\brancher/rPc_current_reg3[12] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2097_  (.CLK(clknet_leaf_31_clk),
    .D(\brancher/_0013_ ),
    .Q(\brancher/rPc_current_reg3[13] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2098_  (.CLK(clknet_leaf_26_clk),
    .D(\brancher/_0014_ ),
    .Q(\brancher/rPc_current_reg3[14] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2099_  (.CLK(clknet_leaf_41_clk),
    .D(\brancher/_0015_ ),
    .Q(\brancher/rPc_current_reg3[15] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2100_  (.CLK(clknet_leaf_26_clk),
    .D(\brancher/_0016_ ),
    .Q(\brancher/rPc_current_reg3[16] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2101_  (.CLK(clknet_leaf_40_clk),
    .D(\brancher/_0017_ ),
    .Q(\brancher/rPc_current_reg3[17] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2102_  (.CLK(clknet_leaf_40_clk),
    .D(\brancher/_0018_ ),
    .Q(\brancher/rPc_current_reg3[18] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2103_  (.CLK(clknet_leaf_32_clk),
    .D(\brancher/_0019_ ),
    .Q(\brancher/rPc_current_reg3[19] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2104_  (.CLK(clknet_leaf_32_clk),
    .D(\brancher/_0020_ ),
    .Q(\brancher/rPc_current_reg3[20] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2105_  (.CLK(clknet_leaf_33_clk),
    .D(\brancher/_0021_ ),
    .Q(\brancher/rPc_current_reg3[21] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2106_  (.CLK(clknet_leaf_32_clk),
    .D(\brancher/_0022_ ),
    .Q(\brancher/rPc_current_reg3[22] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2107_  (.CLK(clknet_leaf_33_clk),
    .D(\brancher/_0023_ ),
    .Q(\brancher/rPc_current_reg3[23] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2108_  (.CLK(clknet_leaf_34_clk),
    .D(\brancher/_0024_ ),
    .Q(\brancher/rPc_current_reg3[24] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2109_  (.CLK(clknet_leaf_34_clk),
    .D(\brancher/_0025_ ),
    .Q(\brancher/rPc_current_reg3[25] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2110_  (.CLK(clknet_leaf_33_clk),
    .D(\brancher/_0026_ ),
    .Q(\brancher/rPc_current_reg3[26] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2111_  (.CLK(clknet_leaf_34_clk),
    .D(\brancher/_0027_ ),
    .Q(\brancher/rPc_current_reg3[27] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2112_  (.CLK(clknet_leaf_34_clk),
    .D(\brancher/_0028_ ),
    .Q(\brancher/rPc_current_reg3[28] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2113_  (.CLK(clknet_leaf_37_clk),
    .D(\brancher/_0029_ ),
    .Q(\brancher/rPc_current_reg3[29] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2114_  (.CLK(clknet_leaf_34_clk),
    .D(\brancher/_0030_ ),
    .Q(\brancher/rPc_current_reg3[30] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2115_  (.CLK(clknet_leaf_37_clk),
    .D(\brancher/_0031_ ),
    .Q(\brancher/rPc_current_reg3[31] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2116_  (.CLK(clknet_leaf_51_clk),
    .D(net1075),
    .Q(\brancher/rAdder_jal[1] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2117_  (.CLK(clknet_leaf_47_clk),
    .D(net1401),
    .Q(\brancher/rAdder_jal[2] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2118_  (.CLK(clknet_leaf_62_clk),
    .D(net1152),
    .Q(\brancher/rAdder_jal[3] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2119_  (.CLK(clknet_leaf_62_clk),
    .D(net1162),
    .Q(\brancher/rAdder_jal[4] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2120_  (.CLK(clknet_leaf_62_clk),
    .D(net1171),
    .Q(\brancher/rAdder_jal[5] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2121_  (.CLK(clknet_leaf_61_clk),
    .D(\imm21_j[5] ),
    .Q(\brancher/rAdder_jal[6] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2122_  (.CLK(clknet_leaf_56_clk),
    .D(\imm21_j[6] ),
    .Q(\brancher/rAdder_jal[7] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2123_  (.CLK(clknet_leaf_57_clk),
    .D(\imm21_j[7] ),
    .Q(\brancher/rAdder_jal[8] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2124_  (.CLK(clknet_leaf_46_clk),
    .D(\imm21_j[8] ),
    .Q(\brancher/rAdder_jal[9] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2125_  (.CLK(clknet_leaf_46_clk),
    .D(\imm21_j[9] ),
    .Q(\brancher/rAdder_jal[10] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2126_  (.CLK(clknet_leaf_45_clk),
    .D(\imm21_j[10] ),
    .Q(\brancher/rAdder_jal[11] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2127_  (.CLK(clknet_leaf_46_clk),
    .D(net1138),
    .Q(\brancher/rAdder_jal[12] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2128_  (.CLK(clknet_leaf_43_clk),
    .D(net1191),
    .Q(\brancher/rAdder_jal[13] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2129_  (.CLK(clknet_leaf_43_clk),
    .D(net1189),
    .Q(\brancher/rAdder_jal[14] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2130_  (.CLK(clknet_leaf_41_clk),
    .D(net1157),
    .Q(\brancher/rAdder_jal[15] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2131_  (.CLK(clknet_leaf_41_clk),
    .D(net1134),
    .Q(\brancher/rAdder_jal[16] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2132_  (.CLK(clknet_leaf_40_clk),
    .D(net1153),
    .Q(\brancher/rAdder_jal[17] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2133_  (.CLK(clknet_leaf_43_clk),
    .D(net1149),
    .Q(\brancher/rAdder_jal[18] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2134_  (.CLK(clknet_leaf_32_clk),
    .D(net1141),
    .Q(\brancher/rAdder_jal[19] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2135_  (.CLK(clknet_leaf_32_clk),
    .D(net1148),
    .Q(\brancher/rAdder_jal[20] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2136_  (.CLK(clknet_leaf_32_clk),
    .D(\imm21_j[20] ),
    .Q(\brancher/rAdder_jal[21] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2137_  (.CLK(clknet_leaf_48_clk),
    .D(net899),
    .Q(\brancher/rOp_jalr ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2138_  (.CLK(clknet_leaf_54_clk),
    .D(\wAluOut[1] ),
    .Q(\brancher/rAlu_result[1] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2139_  (.CLK(clknet_leaf_56_clk),
    .D(\wAluOut[2] ),
    .Q(\brancher/rAlu_result[2] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2140_  (.CLK(clknet_leaf_55_clk),
    .D(\wAluOut[3] ),
    .Q(\brancher/rAlu_result[3] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2141_  (.CLK(clknet_leaf_58_clk),
    .D(\wAluOut[4] ),
    .Q(\brancher/rAlu_result[4] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2142_  (.CLK(clknet_leaf_58_clk),
    .D(\wAluOut[5] ),
    .Q(\brancher/rAlu_result[5] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2143_  (.CLK(clknet_leaf_88_clk),
    .D(\wAluOut[6] ),
    .Q(\brancher/rAlu_result[6] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2144_  (.CLK(clknet_leaf_56_clk),
    .D(\wAluOut[7] ),
    .Q(\brancher/rAlu_result[7] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2145_  (.CLK(clknet_leaf_55_clk),
    .D(\wAluOut[8] ),
    .Q(\brancher/rAlu_result[8] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2146_  (.CLK(clknet_leaf_57_clk),
    .D(\wAluOut[9] ),
    .Q(\brancher/rAlu_result[9] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2147_  (.CLK(clknet_leaf_58_clk),
    .D(\wAluOut[10] ),
    .Q(\brancher/rAlu_result[10] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2148_  (.CLK(clknet_leaf_58_clk),
    .D(\wAluOut[11] ),
    .Q(\brancher/rAlu_result[11] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2149_  (.CLK(clknet_leaf_57_clk),
    .D(\wAluOut[12] ),
    .Q(\brancher/rAlu_result[12] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2150_  (.CLK(clknet_leaf_58_clk),
    .D(\wAluOut[13] ),
    .Q(\brancher/rAlu_result[13] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2151_  (.CLK(clknet_leaf_89_clk),
    .D(\wAluOut[14] ),
    .Q(\brancher/rAlu_result[14] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2152_  (.CLK(clknet_leaf_58_clk),
    .D(\wAluOut[15] ),
    .Q(\brancher/rAlu_result[15] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2153_  (.CLK(clknet_leaf_57_clk),
    .D(\wAluOut[16] ),
    .Q(\brancher/rAlu_result[16] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2154_  (.CLK(clknet_leaf_56_clk),
    .D(\wAluOut[17] ),
    .Q(\brancher/rAlu_result[17] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2155_  (.CLK(clknet_leaf_56_clk),
    .D(\wAluOut[18] ),
    .Q(\brancher/rAlu_result[18] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2156_  (.CLK(clknet_leaf_56_clk),
    .D(\wAluOut[19] ),
    .Q(\brancher/rAlu_result[19] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2157_  (.CLK(clknet_leaf_56_clk),
    .D(\wAluOut[20] ),
    .Q(\brancher/rAlu_result[20] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2158_  (.CLK(clknet_leaf_56_clk),
    .D(\wAluOut[21] ),
    .Q(\brancher/rAlu_result[21] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2159_  (.CLK(clknet_leaf_56_clk),
    .D(\wAluOut[22] ),
    .Q(\brancher/rAlu_result[22] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2160_  (.CLK(clknet_leaf_52_clk),
    .D(\wAluOut[23] ),
    .Q(\brancher/rAlu_result[23] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2161_  (.CLK(clknet_leaf_52_clk),
    .D(\wAluOut[24] ),
    .Q(\brancher/rAlu_result[24] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2162_  (.CLK(clknet_leaf_52_clk),
    .D(\wAluOut[25] ),
    .Q(\brancher/rAlu_result[25] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2163_  (.CLK(clknet_leaf_53_clk),
    .D(\wAluOut[26] ),
    .Q(\brancher/rAlu_result[26] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2164_  (.CLK(clknet_leaf_52_clk),
    .D(\wAluOut[27] ),
    .Q(\brancher/rAlu_result[27] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2165_  (.CLK(clknet_leaf_52_clk),
    .D(\wAluOut[28] ),
    .Q(\brancher/rAlu_result[28] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2166_  (.CLK(clknet_leaf_53_clk),
    .D(\wAluOut[29] ),
    .Q(\brancher/rAlu_result[29] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2167_  (.CLK(clknet_leaf_52_clk),
    .D(\wAluOut[30] ),
    .Q(\brancher/rAlu_result[30] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2168_  (.CLK(clknet_leaf_53_clk),
    .D(\wAluOut[31] ),
    .Q(\brancher/rAlu_result[31] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2169_  (.CLK(clknet_leaf_25_clk),
    .D(net320),
    .Q(\brancher/rOp_jal ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2170_  (.CLK(clknet_leaf_60_clk),
    .D(net896),
    .Q(\brancher/rOp_b_type ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2171_  (.CLK(clknet_leaf_47_clk),
    .D(net1074),
    .Q(\brancher/rAdder_b[1] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2172_  (.CLK(clknet_leaf_63_clk),
    .D(net1151),
    .Q(\brancher/rAdder_b[2] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2173_  (.CLK(clknet_leaf_63_clk),
    .D(net1144),
    .Q(\brancher/rAdder_b[3] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2174_  (.CLK(clknet_leaf_63_clk),
    .D(net1147),
    .Q(\brancher/rAdder_b[4] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2175_  (.CLK(clknet_leaf_63_clk),
    .D(net1139),
    .Q(\brancher/rAdder_b[5] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2176_  (.CLK(clknet_leaf_61_clk),
    .D(\imm13_b[5] ),
    .Q(\brancher/rAdder_b[6] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2177_  (.CLK(clknet_leaf_52_clk),
    .D(\imm13_b[6] ),
    .Q(\brancher/rAdder_b[7] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2178_  (.CLK(clknet_leaf_57_clk),
    .D(\imm13_b[7] ),
    .Q(\brancher/rAdder_b[8] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2179_  (.CLK(clknet_leaf_46_clk),
    .D(\imm13_b[8] ),
    .Q(\brancher/rAdder_b[9] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2180_  (.CLK(clknet_leaf_46_clk),
    .D(\imm13_b[9] ),
    .Q(\brancher/rAdder_b[10] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2181_  (.CLK(clknet_leaf_45_clk),
    .D(\imm13_b[10] ),
    .Q(\brancher/rAdder_b[11] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2182_  (.CLK(clknet_leaf_45_clk),
    .D(net1135),
    .Q(\brancher/rAdder_b[12] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2183_  (.CLK(clknet_leaf_26_clk),
    .D(\imm13_b[12] ),
    .Q(\brancher/rAdder_b[13] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2184_  (.CLK(clknet_leaf_54_clk),
    .D(\brancher/_0032_ ),
    .Q(\brancher/rPc_current_reg1[0] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2185_  (.CLK(clknet_leaf_54_clk),
    .D(\brancher/_0033_ ),
    .Q(\brancher/rPc_current_reg1[1] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2186_  (.CLK(clknet_leaf_56_clk),
    .D(\brancher/_0034_ ),
    .Q(\brancher/rPc_current_reg1[2] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2187_  (.CLK(clknet_leaf_54_clk),
    .D(\brancher/_0035_ ),
    .Q(\brancher/rPc_current_reg1[3] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2188_  (.CLK(clknet_leaf_61_clk),
    .D(\brancher/_0036_ ),
    .Q(\brancher/rPc_current_reg1[4] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2189_  (.CLK(clknet_leaf_56_clk),
    .D(\brancher/_0037_ ),
    .Q(\brancher/rPc_current_reg1[5] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2190_  (.CLK(clknet_leaf_58_clk),
    .D(\brancher/_0038_ ),
    .Q(\brancher/rPc_current_reg1[6] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2191_  (.CLK(clknet_leaf_54_clk),
    .D(\brancher/_0039_ ),
    .Q(\brancher/rPc_current_reg1[7] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2192_  (.CLK(clknet_leaf_56_clk),
    .D(\brancher/_0040_ ),
    .Q(\brancher/rPc_current_reg1[8] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2193_  (.CLK(clknet_leaf_56_clk),
    .D(\brancher/_0041_ ),
    .Q(\brancher/rPc_current_reg1[9] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2194_  (.CLK(clknet_leaf_59_clk),
    .D(\brancher/_0042_ ),
    .Q(\brancher/rPc_current_reg1[10] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2195_  (.CLK(clknet_leaf_58_clk),
    .D(\brancher/_0043_ ),
    .Q(\brancher/rPc_current_reg1[11] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2196_  (.CLK(clknet_leaf_25_clk),
    .D(\brancher/_0044_ ),
    .Q(\brancher/rPc_current_reg1[12] ));
 sky130_fd_sc_hd__dfxtp_2 \brancher/_2197_  (.CLK(clknet_leaf_31_clk),
    .D(\brancher/_0045_ ),
    .Q(\brancher/rPc_current_reg1[13] ));
 sky130_fd_sc_hd__dfxtp_2 \brancher/_2198_  (.CLK(clknet_leaf_36_clk),
    .D(\brancher/_0046_ ),
    .Q(\brancher/rPc_current_reg1[14] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2199_  (.CLK(clknet_leaf_41_clk),
    .D(\brancher/_0047_ ),
    .Q(\brancher/rPc_current_reg1[15] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2200_  (.CLK(clknet_leaf_31_clk),
    .D(\brancher/_0048_ ),
    .Q(\brancher/rPc_current_reg1[16] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2201_  (.CLK(clknet_leaf_41_clk),
    .D(\brancher/_0049_ ),
    .Q(\brancher/rPc_current_reg1[17] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2202_  (.CLK(clknet_leaf_40_clk),
    .D(\brancher/_0050_ ),
    .Q(\brancher/rPc_current_reg1[18] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2203_  (.CLK(clknet_leaf_36_clk),
    .D(\brancher/_0051_ ),
    .Q(\brancher/rPc_current_reg1[19] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2204_  (.CLK(clknet_leaf_32_clk),
    .D(\brancher/_0052_ ),
    .Q(\brancher/rPc_current_reg1[20] ));
 sky130_fd_sc_hd__dfxtp_2 \brancher/_2205_  (.CLK(clknet_leaf_52_clk),
    .D(\brancher/_0053_ ),
    .Q(\brancher/rPc_current_reg1[21] ));
 sky130_fd_sc_hd__dfxtp_2 \brancher/_2206_  (.CLK(clknet_leaf_52_clk),
    .D(\brancher/_0054_ ),
    .Q(\brancher/rPc_current_reg1[22] ));
 sky130_fd_sc_hd__dfxtp_2 \brancher/_2207_  (.CLK(clknet_leaf_53_clk),
    .D(\brancher/_0055_ ),
    .Q(\brancher/rPc_current_reg1[23] ));
 sky130_fd_sc_hd__dfxtp_2 \brancher/_2208_  (.CLK(clknet_leaf_53_clk),
    .D(\brancher/_0056_ ),
    .Q(\brancher/rPc_current_reg1[24] ));
 sky130_fd_sc_hd__dfxtp_2 \brancher/_2209_  (.CLK(clknet_leaf_53_clk),
    .D(\brancher/_0057_ ),
    .Q(\brancher/rPc_current_reg1[25] ));
 sky130_fd_sc_hd__dfxtp_2 \brancher/_2210_  (.CLK(clknet_leaf_53_clk),
    .D(\brancher/_0058_ ),
    .Q(\brancher/rPc_current_reg1[26] ));
 sky130_fd_sc_hd__dfxtp_2 \brancher/_2211_  (.CLK(clknet_leaf_54_clk),
    .D(\brancher/_0059_ ),
    .Q(\brancher/rPc_current_reg1[27] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2212_  (.CLK(clknet_leaf_53_clk),
    .D(\brancher/_0060_ ),
    .Q(\brancher/rPc_current_reg1[28] ));
 sky130_fd_sc_hd__dfxtp_2 \brancher/_2213_  (.CLK(clknet_leaf_53_clk),
    .D(\brancher/_0061_ ),
    .Q(\brancher/rPc_current_reg1[29] ));
 sky130_fd_sc_hd__dfxtp_2 \brancher/_2214_  (.CLK(clknet_leaf_53_clk),
    .D(\brancher/_0062_ ),
    .Q(\brancher/rPc_current_reg1[30] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2215_  (.CLK(clknet_leaf_53_clk),
    .D(\brancher/_0063_ ),
    .Q(\brancher/rPc_current_reg1[31] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2216_  (.CLK(clknet_leaf_53_clk),
    .D(\brancher/_0064_ ),
    .Q(\brancher/rPc_current_reg2[0] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2217_  (.CLK(clknet_leaf_53_clk),
    .D(\brancher/_0065_ ),
    .Q(\brancher/rPc_current_reg2[1] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2218_  (.CLK(clknet_leaf_56_clk),
    .D(\brancher/_0066_ ),
    .Q(\brancher/rPc_current_reg2[2] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2219_  (.CLK(clknet_leaf_60_clk),
    .D(\brancher/_0067_ ),
    .Q(\brancher/rPc_current_reg2[3] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2220_  (.CLK(clknet_leaf_60_clk),
    .D(\brancher/_0068_ ),
    .Q(\brancher/rPc_current_reg2[4] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2221_  (.CLK(clknet_leaf_57_clk),
    .D(\brancher/_0069_ ),
    .Q(\brancher/rPc_current_reg2[5] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2222_  (.CLK(clknet_leaf_58_clk),
    .D(\brancher/_0070_ ),
    .Q(\brancher/rPc_current_reg2[6] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2223_  (.CLK(clknet_leaf_54_clk),
    .D(\brancher/_0071_ ),
    .Q(\brancher/rPc_current_reg2[7] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2224_  (.CLK(clknet_leaf_57_clk),
    .D(\brancher/_0072_ ),
    .Q(\brancher/rPc_current_reg2[8] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2225_  (.CLK(clknet_leaf_56_clk),
    .D(\brancher/_0073_ ),
    .Q(\brancher/rPc_current_reg2[9] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2226_  (.CLK(clknet_leaf_60_clk),
    .D(\brancher/_0074_ ),
    .Q(\brancher/rPc_current_reg2[10] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2227_  (.CLK(clknet_leaf_63_clk),
    .D(\brancher/_0075_ ),
    .Q(\brancher/rPc_current_reg2[11] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2228_  (.CLK(clknet_leaf_25_clk),
    .D(\brancher/_0076_ ),
    .Q(\brancher/rPc_current_reg2[12] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2229_  (.CLK(clknet_leaf_31_clk),
    .D(\brancher/_0077_ ),
    .Q(\brancher/rPc_current_reg2[13] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2230_  (.CLK(clknet_leaf_26_clk),
    .D(\brancher/_0078_ ),
    .Q(\brancher/rPc_current_reg2[14] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2231_  (.CLK(clknet_leaf_25_clk),
    .D(\brancher/_0079_ ),
    .Q(\brancher/rPc_current_reg2[15] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2232_  (.CLK(clknet_leaf_26_clk),
    .D(\brancher/_0080_ ),
    .Q(\brancher/rPc_current_reg2[16] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2233_  (.CLK(clknet_leaf_41_clk),
    .D(\brancher/_0081_ ),
    .Q(\brancher/rPc_current_reg2[17] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2234_  (.CLK(clknet_leaf_40_clk),
    .D(\brancher/_0082_ ),
    .Q(\brancher/rPc_current_reg2[18] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2235_  (.CLK(clknet_leaf_32_clk),
    .D(\brancher/_0083_ ),
    .Q(\brancher/rPc_current_reg2[19] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2236_  (.CLK(clknet_leaf_32_clk),
    .D(\brancher/_0084_ ),
    .Q(\brancher/rPc_current_reg2[20] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2237_  (.CLK(clknet_leaf_33_clk),
    .D(\brancher/_0085_ ),
    .Q(\brancher/rPc_current_reg2[21] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2238_  (.CLK(clknet_leaf_35_clk),
    .D(\brancher/_0086_ ),
    .Q(\brancher/rPc_current_reg2[22] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2239_  (.CLK(clknet_leaf_33_clk),
    .D(\brancher/_0087_ ),
    .Q(\brancher/rPc_current_reg2[23] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2240_  (.CLK(clknet_leaf_35_clk),
    .D(\brancher/_0088_ ),
    .Q(\brancher/rPc_current_reg2[24] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2241_  (.CLK(clknet_leaf_34_clk),
    .D(\brancher/_0089_ ),
    .Q(\brancher/rPc_current_reg2[25] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2242_  (.CLK(clknet_leaf_33_clk),
    .D(\brancher/_0090_ ),
    .Q(\brancher/rPc_current_reg2[26] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2243_  (.CLK(clknet_leaf_34_clk),
    .D(\brancher/_0091_ ),
    .Q(\brancher/rPc_current_reg2[27] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2244_  (.CLK(clknet_leaf_34_clk),
    .D(\brancher/_0092_ ),
    .Q(\brancher/rPc_current_reg2[28] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2245_  (.CLK(clknet_leaf_37_clk),
    .D(\brancher/_0093_ ),
    .Q(\brancher/rPc_current_reg2[29] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2246_  (.CLK(clknet_leaf_37_clk),
    .D(\brancher/_0094_ ),
    .Q(\brancher/rPc_current_reg2[30] ));
 sky130_fd_sc_hd__dfxtp_1 \brancher/_2247_  (.CLK(clknet_leaf_37_clk),
    .D(\brancher/_0095_ ),
    .Q(\brancher/rPc_current_reg2[31] ));
 sky130_fd_sc_hd__inv_8 \dec/_301_  (.A(net886),
    .Y(\dec/_061_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_302_  (.A(\dec/_061_ ),
    .X(\dec/_062_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_303_  (.A(\dec/_062_ ),
    .X(\dec/_063_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_304_  (.A1(net889),
    .A2(\dec/rInstrustion2[20] ),
    .B1(net882),
    .X(\dec/_064_ ));
 sky130_fd_sc_hd__inv_4 \dec/_305_  (.A(net888),
    .Y(\dec/_065_ ));
 sky130_fd_sc_hd__buf_6 \dec/_306_  (.A(\dec/_065_ ),
    .X(\dec/_066_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_307_  (.A(\dec/_066_ ),
    .X(\dec/_067_ ));
 sky130_fd_sc_hd__and3_1 \dec/_308_  (.A(\dec/_067_ ),
    .B(net1069),
    .C(net46),
    .X(\dec/_068_ ));
 sky130_fd_sc_hd__o221a_2 \dec/_309_  (.A1(\dec/_063_ ),
    .A2(\dec/rInstrustion1[20] ),
    .B1(\dec/_064_ ),
    .B2(\dec/_068_ ),
    .C1(net1015),
    .X(\dec/_069_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_310_  (.A(wJumping),
    .B(net240),
    .Y(\dec/_070_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_311_  (.A(\dec/_070_ ),
    .X(\dec/_071_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_312_  (.A(\dec/_071_ ),
    .X(\dec/_072_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_313_  (.A1(\reg_s2[0] ),
    .A2(net243),
    .B1(\dec/_069_ ),
    .B2(\dec/_072_ ),
    .X(\wReg_s2_out[0] ));
 sky130_fd_sc_hd__a21o_1 \dec/_314_  (.A1(net889),
    .A2(\dec/rInstrustion2[21] ),
    .B1(net882),
    .X(\dec/_073_ ));
 sky130_fd_sc_hd__and3_1 \dec/_315_  (.A(\dec/_067_ ),
    .B(net1069),
    .C(net47),
    .X(\dec/_074_ ));
 sky130_fd_sc_hd__o221a_2 \dec/_316_  (.A1(\dec/_063_ ),
    .A2(\dec/rInstrustion1[21] ),
    .B1(\dec/_073_ ),
    .B2(\dec/_074_ ),
    .C1(net1015),
    .X(\dec/_075_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_317_  (.A(\dec/_071_ ),
    .X(\dec/_076_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_318_  (.A1(net260),
    .A2(\reg_s2[1] ),
    .B1(\dec/_075_ ),
    .B2(\dec/_076_ ),
    .X(\wReg_s2_out[1] ));
 sky130_fd_sc_hd__a21o_1 \dec/_319_  (.A1(net889),
    .A2(\dec/rInstrustion2[22] ),
    .B1(net882),
    .X(\dec/_077_ ));
 sky130_fd_sc_hd__and3_1 \dec/_320_  (.A(\dec/_067_ ),
    .B(net1069),
    .C(net48),
    .X(\dec/_078_ ));
 sky130_fd_sc_hd__o221a_2 \dec/_321_  (.A1(\dec/_063_ ),
    .A2(\dec/rInstrustion1[22] ),
    .B1(\dec/_077_ ),
    .B2(\dec/_078_ ),
    .C1(net1015),
    .X(\dec/_079_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_322_  (.A1(net260),
    .A2(\reg_s2[2] ),
    .B1(\dec/_079_ ),
    .B2(\dec/_076_ ),
    .X(\wReg_s2_out[2] ));
 sky130_fd_sc_hd__a21o_1 \dec/_323_  (.A1(net889),
    .A2(\dec/rInstrustion2[23] ),
    .B1(net882),
    .X(\dec/_080_ ));
 sky130_fd_sc_hd__and3_1 \dec/_324_  (.A(\dec/_067_ ),
    .B(net1069),
    .C(net49),
    .X(\dec/_081_ ));
 sky130_fd_sc_hd__o221a_2 \dec/_325_  (.A1(\dec/_063_ ),
    .A2(\dec/rInstrustion1[23] ),
    .B1(\dec/_080_ ),
    .B2(\dec/_081_ ),
    .C1(net1016),
    .X(\dec/_082_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_326_  (.A1(net260),
    .A2(\reg_s2[3] ),
    .B1(\dec/_082_ ),
    .B2(\dec/_076_ ),
    .X(\wReg_s2_out[3] ));
 sky130_fd_sc_hd__a21o_1 \dec/_327_  (.A1(net889),
    .A2(\dec/rInstrustion2[24] ),
    .B1(net882),
    .X(\dec/_083_ ));
 sky130_fd_sc_hd__and3_1 \dec/_328_  (.A(\dec/_067_ ),
    .B(net1069),
    .C(net50),
    .X(\dec/_084_ ));
 sky130_fd_sc_hd__o221a_2 \dec/_329_  (.A1(\dec/_063_ ),
    .A2(\dec/rInstrustion1[24] ),
    .B1(\dec/_083_ ),
    .B2(\dec/_084_ ),
    .C1(net1015),
    .X(\dec/_085_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_330_  (.A1(net260),
    .A2(\reg_s2[4] ),
    .B1(\dec/_085_ ),
    .B2(\dec/_076_ ),
    .X(\wReg_s2_out[4] ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_331_  (.A(\dec/_062_ ),
    .X(\dec/_086_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_332_  (.A(\dec/_086_ ),
    .X(\dec/_087_ ));
 sky130_fd_sc_hd__inv_2 \dec/_333_  (.A(net1071),
    .Y(\dec/_088_ ));
 sky130_fd_sc_hd__nor2_2 \dec/_334_  (.A(net892),
    .B(\dec/_088_ ),
    .Y(\dec/_089_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_335_  (.A(\dec/_089_ ),
    .X(\dec/_090_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_336_  (.A(\dec/_090_ ),
    .X(\dec/_091_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_337_  (.A(\dec/_091_ ),
    .B(net40),
    .Y(\dec/_092_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_338_  (.A(net893),
    .B(\dec/rInstrustion2[15] ),
    .Y(\dec/_093_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_339_  (.A(\dec/_063_ ),
    .X(\dec/_094_ ));
 sky130_fd_sc_hd__inv_2 \dec/_340_  (.A(net1017),
    .Y(\dec/_095_ ));
 sky130_fd_sc_hd__inv_2 \dec/_341_  (.A(\dec/_070_ ),
    .Y(\dec/_096_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_342_  (.A(\dec/_095_ ),
    .B(\dec/_096_ ),
    .Y(\dec/_097_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \dec/_343_  (.A(\dec/_097_ ),
    .X(\dec/_098_ ));
 sky130_fd_sc_hd__o21ai_1 \dec/_344_  (.A1(\dec/_094_ ),
    .A2(\dec/rInstrustion1[15] ),
    .B1(\dec/_098_ ),
    .Y(\dec/_099_ ));
 sky130_fd_sc_hd__a31o_1 \dec/_345_  (.A1(\dec/_087_ ),
    .A2(\dec/_092_ ),
    .A3(\dec/_093_ ),
    .B1(\dec/_099_ ),
    .X(\dec/_100_ ));
 sky130_fd_sc_hd__a21bo_1 \dec/_346_  (.A1(net243),
    .A2(\reg_s1[0] ),
    .B1_N(\dec/_100_ ),
    .X(\wReg_s1_out[0] ));
 sky130_fd_sc_hd__nand2_1 \dec/_347_  (.A(\dec/_091_ ),
    .B(net41),
    .Y(\dec/_101_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_348_  (.A(net888),
    .B(\dec/rInstrustion2[16] ),
    .Y(\dec/_102_ ));
 sky130_fd_sc_hd__o21ai_1 \dec/_349_  (.A1(\dec/_094_ ),
    .A2(\dec/rInstrustion1[16] ),
    .B1(\dec/_098_ ),
    .Y(\dec/_103_ ));
 sky130_fd_sc_hd__a31o_1 \dec/_350_  (.A1(\dec/_087_ ),
    .A2(\dec/_101_ ),
    .A3(\dec/_102_ ),
    .B1(\dec/_103_ ),
    .X(\dec/_104_ ));
 sky130_fd_sc_hd__a21bo_1 \dec/_351_  (.A1(net260),
    .A2(\reg_s1[1] ),
    .B1_N(\dec/_104_ ),
    .X(\wReg_s1_out[1] ));
 sky130_fd_sc_hd__nand2_1 \dec/_352_  (.A(\dec/_091_ ),
    .B(net42),
    .Y(\dec/_105_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_353_  (.A(net892),
    .B(\dec/rInstrustion2[17] ),
    .Y(\dec/_106_ ));
 sky130_fd_sc_hd__o21ai_1 \dec/_354_  (.A1(\dec/_094_ ),
    .A2(\dec/rInstrustion1[17] ),
    .B1(\dec/_098_ ),
    .Y(\dec/_107_ ));
 sky130_fd_sc_hd__a31o_1 \dec/_355_  (.A1(\dec/_087_ ),
    .A2(\dec/_105_ ),
    .A3(\dec/_106_ ),
    .B1(\dec/_107_ ),
    .X(\dec/_108_ ));
 sky130_fd_sc_hd__a21bo_1 \dec/_356_  (.A1(net243),
    .A2(\reg_s1[2] ),
    .B1_N(\dec/_108_ ),
    .X(\wReg_s1_out[2] ));
 sky130_fd_sc_hd__nand2_1 \dec/_357_  (.A(\dec/_091_ ),
    .B(net43),
    .Y(\dec/_109_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_358_  (.A(net888),
    .B(\dec/rInstrustion2[18] ),
    .Y(\dec/_110_ ));
 sky130_fd_sc_hd__o21ai_1 \dec/_359_  (.A1(\dec/_094_ ),
    .A2(\dec/rInstrustion1[18] ),
    .B1(\dec/_098_ ),
    .Y(\dec/_111_ ));
 sky130_fd_sc_hd__a31o_1 \dec/_360_  (.A1(\dec/_087_ ),
    .A2(\dec/_109_ ),
    .A3(\dec/_110_ ),
    .B1(\dec/_111_ ),
    .X(\dec/_112_ ));
 sky130_fd_sc_hd__a21bo_1 \dec/_361_  (.A1(net243),
    .A2(net2155),
    .B1_N(\dec/_112_ ),
    .X(\wReg_s1_out[3] ));
 sky130_fd_sc_hd__nand2_1 \dec/_362_  (.A(\dec/_091_ ),
    .B(net44),
    .Y(\dec/_113_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_363_  (.A(net895),
    .B(\dec/rInstrustion2[19] ),
    .Y(\dec/_114_ ));
 sky130_fd_sc_hd__o21ai_1 \dec/_364_  (.A1(\dec/_094_ ),
    .A2(\dec/rInstrustion1[19] ),
    .B1(\dec/_097_ ),
    .Y(\dec/_115_ ));
 sky130_fd_sc_hd__a31o_1 \dec/_365_  (.A1(\dec/_087_ ),
    .A2(\dec/_113_ ),
    .A3(\dec/_114_ ),
    .B1(\dec/_115_ ),
    .X(\dec/_116_ ));
 sky130_fd_sc_hd__a21bo_1 \dec/_366_  (.A1(net262),
    .A2(\reg_s1[4] ),
    .B1_N(\dec/_116_ ),
    .X(\wReg_s1_out[4] ));
 sky130_fd_sc_hd__nand2_1 \dec/_367_  (.A(net889),
    .B(\dec/rInstrustion2[0] ),
    .Y(\dec/_117_ ));
 sky130_fd_sc_hd__buf_6 \dec/_368_  (.A(\dec/_061_ ),
    .X(\dec/_118_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_369_  (.A(\dec/_117_ ),
    .B(\dec/_118_ ),
    .Y(\dec/_119_ ));
 sky130_fd_sc_hd__inv_2 \dec/_370_  (.A(\dec/_119_ ),
    .Y(\dec/_120_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_371_  (.A(\dec/_067_ ),
    .B(net1069),
    .C(net34),
    .Y(\dec/_121_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_372_  (.A(\dec/_120_ ),
    .B(\dec/_121_ ),
    .Y(\dec/_122_ ));
 sky130_fd_sc_hd__o21ai_1 \dec/_373_  (.A1(\dec/rInstrustion1[0] ),
    .A2(\dec/_118_ ),
    .B1(net1017),
    .Y(\dec/_123_ ));
 sky130_fd_sc_hd__inv_2 \dec/_374_  (.A(\dec/_123_ ),
    .Y(\dec/_124_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_375_  (.A(\dec/_122_ ),
    .B(\dec/_124_ ),
    .Y(\dec/_125_ ));
 sky130_fd_sc_hd__a21oi_1 \dec/_376_  (.A1(net890),
    .A2(\dec/rInstrustion2[1] ),
    .B1(net882),
    .Y(\dec/_126_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_377_  (.A(\dec/_066_ ),
    .B(net1070),
    .C(net45),
    .Y(\dec/_127_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_378_  (.A(\dec/_126_ ),
    .B(\dec/_127_ ),
    .Y(\dec/_128_ ));
 sky130_fd_sc_hd__o21ai_1 \dec/_379_  (.A1(\dec/rInstrustion1[1] ),
    .A2(\dec/_118_ ),
    .B1(net1017),
    .Y(\dec/_129_ ));
 sky130_fd_sc_hd__clkinvlp_2 \dec/_380_  (.A(\dec/_129_ ),
    .Y(\dec/_130_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_381_  (.A(\dec/_128_ ),
    .B(\dec/_130_ ),
    .Y(\dec/_131_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_382_  (.A(\dec/_125_ ),
    .B(\dec/_131_ ),
    .Y(\dec/_132_ ));
 sky130_fd_sc_hd__a21oi_1 \dec/_383_  (.A1(net894),
    .A2(\dec/rInstrustion2[2] ),
    .B1(net887),
    .Y(\dec/_133_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_384_  (.A(\dec/_066_ ),
    .B(net1071),
    .C(net56),
    .Y(\dec/_134_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_385_  (.A(\dec/_133_ ),
    .B(\dec/_134_ ),
    .Y(\dec/_135_ ));
 sky130_fd_sc_hd__o21a_1 \dec/_386_  (.A1(\dec/rInstrustion1[2] ),
    .A2(\dec/_061_ ),
    .B1(net1017),
    .X(\dec/_136_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_387_  (.A(\dec/_135_ ),
    .B(\dec/_136_ ),
    .Y(\dec/_137_ ));
 sky130_fd_sc_hd__inv_2 \dec/_388_  (.A(\dec/_137_ ),
    .Y(\dec/_138_ ));
 sky130_fd_sc_hd__a21oi_1 \dec/_389_  (.A1(net890),
    .A2(\dec/rInstrustion2[3] ),
    .B1(net887),
    .Y(\dec/_139_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_390_  (.A(\dec/_065_ ),
    .B(net1070),
    .C(net59),
    .Y(\dec/_140_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_391_  (.A(\dec/_139_ ),
    .B(\dec/_140_ ),
    .Y(\dec/_141_ ));
 sky130_fd_sc_hd__o21a_1 \dec/_392_  (.A1(\dec/rInstrustion1[3] ),
    .A2(\dec/_061_ ),
    .B1(net1017),
    .X(\dec/_142_ ));
 sky130_fd_sc_hd__nand2_2 \dec/_393_  (.A(\dec/_141_ ),
    .B(\dec/_142_ ),
    .Y(\dec/_143_ ));
 sky130_fd_sc_hd__inv_2 \dec/_394_  (.A(\dec/_143_ ),
    .Y(\dec/_144_ ));
 sky130_fd_sc_hd__and4_1 \dec/_395_  (.A(\dec/_132_ ),
    .B(\dec/_138_ ),
    .C(\dec/_144_ ),
    .D(\dec/_070_ ),
    .X(\dec/_145_ ));
 sky130_fd_sc_hd__a21oi_1 \dec/_396_  (.A1(net894),
    .A2(\dec/rInstrustion2[6] ),
    .B1(net886),
    .Y(\dec/_146_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_397_  (.A(\dec/_066_ ),
    .B(net1071),
    .C(net62),
    .Y(\dec/_147_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_398_  (.A(\dec/_146_ ),
    .B(\dec/_147_ ),
    .Y(\dec/_148_ ));
 sky130_fd_sc_hd__o21a_1 \dec/_399_  (.A1(\dec/rInstrustion1[6] ),
    .A2(\dec/_061_ ),
    .B1(net1017),
    .X(\dec/_149_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_400_  (.A(\dec/_148_ ),
    .B(\dec/_149_ ),
    .Y(\dec/_150_ ));
 sky130_fd_sc_hd__inv_2 \dec/_401_  (.A(\dec/_150_ ),
    .Y(\dec/_151_ ));
 sky130_fd_sc_hd__a21oi_1 \dec/_402_  (.A1(net894),
    .A2(\dec/rInstrustion2[5] ),
    .B1(net886),
    .Y(\dec/_152_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_403_  (.A(\dec/_066_ ),
    .B(net1071),
    .C(net61),
    .Y(\dec/_153_ ));
 sky130_fd_sc_hd__o21ai_1 \dec/_404_  (.A1(\dec/rInstrustion1[5] ),
    .A2(\dec/_118_ ),
    .B1(net1018),
    .Y(\dec/_154_ ));
 sky130_fd_sc_hd__a21oi_2 \dec/_405_  (.A1(\dec/_152_ ),
    .A2(\dec/_153_ ),
    .B1(\dec/_154_ ),
    .Y(\dec/_155_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_406_  (.A(\dec/_066_ ),
    .B(net1072),
    .C(net60),
    .Y(\dec/_156_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_407_  (.A(net894),
    .B(\dec/rInstrustion2[4] ),
    .Y(\dec/_157_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_408_  (.A(\dec/_156_ ),
    .B(\dec/_062_ ),
    .C(\dec/_157_ ),
    .Y(\dec/_158_ ));
 sky130_fd_sc_hd__o21ai_1 \dec/_409_  (.A1(\dec/rInstrustion1[4] ),
    .A2(\dec/_118_ ),
    .B1(net1018),
    .Y(\dec/_159_ ));
 sky130_fd_sc_hd__inv_2 \dec/_410_  (.A(\dec/_159_ ),
    .Y(\dec/_160_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_411_  (.A(\dec/_158_ ),
    .B(\dec/_160_ ),
    .Y(\dec/_161_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_412_  (.A(\dec/_151_ ),
    .B(\dec/_155_ ),
    .C(\dec/_161_ ),
    .Y(\dec/_162_ ));
 sky130_fd_sc_hd__inv_2 \dec/_413_  (.A(\dec/_162_ ),
    .Y(\dec/_163_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_414_  (.A1(net240),
    .A2(net1203),
    .B1(\dec/_145_ ),
    .B2(\dec/_163_ ),
    .X(\dec/_000_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_415_  (.A(net1070),
    .B(net34),
    .Y(\dec/_164_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_416_  (.A(net890),
    .B(\dec/_164_ ),
    .Y(\dec/_165_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_417_  (.A(\dec/_119_ ),
    .B(\dec/_165_ ),
    .Y(\dec/_166_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_418_  (.A(\dec/_123_ ),
    .B(\dec/_166_ ),
    .Y(\dec/_167_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_419_  (.A1(net242),
    .A2(net1183),
    .B1(\dec/_167_ ),
    .B2(\dec/_076_ ),
    .X(\dec/_001_ ));
 sky130_fd_sc_hd__a21oi_1 \dec/_420_  (.A1(\dec/_126_ ),
    .A2(\dec/_127_ ),
    .B1(\dec/_129_ ),
    .Y(\dec/_168_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_421_  (.A1(net242),
    .A2(net1180),
    .B1(\dec/_168_ ),
    .B2(\dec/_076_ ),
    .X(\dec/_002_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_422_  (.A(\dec/_071_ ),
    .X(\dec/_169_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_423_  (.A1(net242),
    .A2(net1184),
    .B1(\dec/_138_ ),
    .B2(\dec/_169_ ),
    .X(\dec/_003_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_424_  (.A1(net242),
    .A2(net1182),
    .B1(\dec/_144_ ),
    .B2(\dec/_169_ ),
    .X(\dec/_004_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_425_  (.A(\dec/_157_ ),
    .B(\dec/_118_ ),
    .Y(\dec/_170_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_426_  (.A(net1072),
    .B(net60),
    .Y(\dec/_171_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_427_  (.A(net894),
    .B(\dec/_171_ ),
    .Y(\dec/_172_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_428_  (.A(\dec/_170_ ),
    .B(\dec/_172_ ),
    .Y(\dec/_173_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_429_  (.A(\dec/_159_ ),
    .B(\dec/_173_ ),
    .Y(\dec/_174_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_430_  (.A1(net238),
    .A2(net1174),
    .B1(\dec/_174_ ),
    .B2(\dec/_169_ ),
    .X(\dec/_005_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_431_  (.A1(net238),
    .A2(net1173),
    .B1(\dec/_155_ ),
    .B2(\dec/_169_ ),
    .X(\dec/_006_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_432_  (.A1(net238),
    .A2(net1172),
    .B1(\dec/_151_ ),
    .B2(\dec/_169_ ),
    .X(\dec/_007_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_433_  (.A(\dec/_152_ ),
    .B(\dec/_153_ ),
    .Y(\dec/_175_ ));
 sky130_fd_sc_hd__inv_2 \dec/_434_  (.A(\dec/_154_ ),
    .Y(\dec/_176_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_435_  (.A(\dec/_175_ ),
    .B(\dec/_176_ ),
    .Y(\dec/_177_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_436_  (.A(\dec/_161_ ),
    .B(\dec/_177_ ),
    .Y(\dec/_178_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_437_  (.A(\dec/_151_ ),
    .B(\dec/_178_ ),
    .Y(\dec/_179_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_438_  (.A(\dec/_137_ ),
    .B(\dec/_143_ ),
    .Y(\dec/_180_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_439_  (.A(\dec/_179_ ),
    .B(\dec/_132_ ),
    .C(\dec/_180_ ),
    .Y(\dec/_181_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_440_  (.A(\dec/_168_ ),
    .B(\dec/_167_ ),
    .Y(\dec/_182_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_441_  (.A(\dec/_138_ ),
    .B(\dec/_143_ ),
    .Y(\dec/_183_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_442_  (.A(\dec/_182_ ),
    .B(\dec/_183_ ),
    .Y(\dec/_184_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_443_  (.A(\dec/_163_ ),
    .B(\dec/_184_ ),
    .Y(\dec/_185_ ));
 sky130_fd_sc_hd__nand2_2 \dec/_444_  (.A(\dec/_181_ ),
    .B(\dec/_185_ ),
    .Y(\dec/_186_ ));
 sky130_fd_sc_hd__buf_6 \dec/_445_  (.A(\dec/_186_ ),
    .X(\dec/_187_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_446_  (.A(\dec/_137_ ),
    .B(\dec/_143_ ),
    .Y(\dec/_188_ ));
 sky130_fd_sc_hd__nor2_2 \dec/_447_  (.A(\dec/_188_ ),
    .B(\dec/_182_ ),
    .Y(\dec/_189_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_448_  (.A(\dec/_155_ ),
    .B(\dec/_174_ ),
    .Y(\dec/_190_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_449_  (.A(\dec/_150_ ),
    .B(\dec/_190_ ),
    .Y(\dec/_191_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_450_  (.A(\dec/_189_ ),
    .B(\dec/_191_ ),
    .Y(\dec/_192_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_451_  (.A(\dec/_174_ ),
    .B(\dec/_150_ ),
    .Y(\dec/_193_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_452_  (.A(\dec/_155_ ),
    .B(\dec/_193_ ),
    .Y(\dec/_194_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_453_  (.A(\dec/_189_ ),
    .B(\dec/_194_ ),
    .Y(\dec/_195_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_454_  (.A(\dec/_189_ ),
    .B(\dec/_179_ ),
    .Y(\dec/_196_ ));
 sky130_fd_sc_hd__nand3_2 \dec/_455_  (.A(\dec/_192_ ),
    .B(\dec/_195_ ),
    .C(\dec/_196_ ),
    .Y(\dec/_197_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_456_  (.A(\dec/_187_ ),
    .B(\dec/_197_ ),
    .Y(\dec/_198_ ));
 sky130_fd_sc_hd__o2bb2ai_1 \dec/_457_  (.A1_N(net245),
    .A2_N(net1160),
    .B1(\dec/_096_ ),
    .B2(\dec/_198_ ),
    .Y(\dec/_008_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_458_  (.A(\dec/_177_ ),
    .B(\dec/_193_ ),
    .Y(\dec/_199_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_459_  (.A(\dec/_070_ ),
    .X(\dec/_200_ ));
 sky130_fd_sc_hd__a32o_1 \dec/_460_  (.A1(\dec/_189_ ),
    .A2(\dec/_199_ ),
    .A3(\dec/_200_ ),
    .B1(net246),
    .B2(net2066),
    .X(\dec/_009_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_461_  (.A(\dec/_132_ ),
    .B(\dec/_138_ ),
    .C(\dec/_143_ ),
    .Y(\dec/_201_ ));
 sky130_fd_sc_hd__or2_1 \dec/_462_  (.A(\dec/_096_ ),
    .B(\dec/_193_ ),
    .X(\dec/_202_ ));
 sky130_fd_sc_hd__a2bb2o_1 \dec/_463_  (.A1_N(\dec/_201_ ),
    .A2_N(\dec/_202_ ),
    .B1(net238),
    .B2(net1170),
    .X(\dec/_010_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_464_  (.A1(net888),
    .A2(\dec/rInstrustion2[8] ),
    .B1(net883),
    .X(\dec/_203_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_465_  (.A1(net64),
    .A2(\dec/_090_ ),
    .B1(\dec/_203_ ),
    .X(\dec/_204_ ));
 sky130_fd_sc_hd__o211a_1 \dec/_466_  (.A1(\dec/_086_ ),
    .A2(\dec/rInstrustion1[8] ),
    .B1(net1019),
    .C1(\dec/_204_ ),
    .X(\dec/_205_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_467_  (.A1(net245),
    .A2(net1151),
    .B1(\dec/_205_ ),
    .B2(\dec/_169_ ),
    .X(\dec/_011_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_468_  (.A1(net888),
    .A2(\dec/rInstrustion2[9] ),
    .B1(net883),
    .X(\dec/_206_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_469_  (.A1(net65),
    .A2(\dec/_090_ ),
    .B1(\dec/_206_ ),
    .X(\dec/_207_ ));
 sky130_fd_sc_hd__o211a_1 \dec/_470_  (.A1(\dec/_086_ ),
    .A2(\dec/rInstrustion1[9] ),
    .B1(net1015),
    .C1(\dec/_207_ ),
    .X(\dec/_208_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_471_  (.A(\dec/_071_ ),
    .X(\dec/_209_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_472_  (.A1(net243),
    .A2(net1144),
    .B1(\dec/_208_ ),
    .B2(\dec/_209_ ),
    .X(\dec/_012_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_473_  (.A1(net891),
    .A2(\dec/rInstrustion2[10] ),
    .B1(net883),
    .X(\dec/_210_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_474_  (.A1(net35),
    .A2(\dec/_090_ ),
    .B1(\dec/_210_ ),
    .X(\dec/_211_ ));
 sky130_fd_sc_hd__o211a_1 \dec/_475_  (.A1(\dec/_086_ ),
    .A2(\dec/rInstrustion1[10] ),
    .B1(net1019),
    .C1(\dec/_211_ ),
    .X(\dec/_212_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_476_  (.A1(net243),
    .A2(net1147),
    .B1(\dec/_212_ ),
    .B2(\dec/_209_ ),
    .X(\dec/_013_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_477_  (.A1(net888),
    .A2(\dec/rInstrustion2[11] ),
    .B1(net883),
    .X(\dec/_213_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_478_  (.A1(net36),
    .A2(\dec/_090_ ),
    .B1(\dec/_213_ ),
    .X(\dec/_214_ ));
 sky130_fd_sc_hd__o211a_1 \dec/_479_  (.A1(\dec/_086_ ),
    .A2(\dec/rInstrustion1[11] ),
    .B1(net1015),
    .C1(\dec/_214_ ),
    .X(\dec/_215_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_480_  (.A1(net244),
    .A2(net1139),
    .B1(\dec/_215_ ),
    .B2(\dec/_209_ ),
    .X(\dec/_014_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_481_  (.A1(net891),
    .A2(\dec/rInstrustion2[7] ),
    .B1(net883),
    .X(\dec/_216_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_482_  (.A1(net63),
    .A2(\dec/_089_ ),
    .B1(\dec/_216_ ),
    .X(\dec/_217_ ));
 sky130_fd_sc_hd__o211a_1 \dec/_483_  (.A1(\dec/_086_ ),
    .A2(\dec/rInstrustion1[7] ),
    .B1(net1019),
    .C1(\dec/_217_ ),
    .X(\dec/_218_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_484_  (.A1(net244),
    .A2(net1135),
    .B1(\dec/_218_ ),
    .B2(\dec/_209_ ),
    .X(\dec/_015_ ));
 sky130_fd_sc_hd__o21bai_1 \dec/_485_  (.A1(\dec/_187_ ),
    .A2(\dec/_197_ ),
    .B1_N(\dec/_069_ ),
    .Y(\dec/_219_ ));
 sky130_fd_sc_hd__inv_2 \dec/_486_  (.A(\dec/_195_ ),
    .Y(\dec/_220_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_487_  (.A(\dec/_192_ ),
    .B(\dec/_196_ ),
    .Y(\dec/_221_ ));
 sky130_fd_sc_hd__nor2_2 \dec/_488_  (.A(\dec/_220_ ),
    .B(\dec/_221_ ),
    .Y(\dec/_222_ ));
 sky130_fd_sc_hd__inv_4 \dec/_489_  (.A(\dec/_186_ ),
    .Y(\dec/_223_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_490_  (.A(\dec/_155_ ),
    .B(\dec/_161_ ),
    .Y(\dec/_224_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_491_  (.A(\dec/_151_ ),
    .B(\dec/_224_ ),
    .Y(\dec/_225_ ));
 sky130_fd_sc_hd__and2_1 \dec/_492_  (.A(\dec/_189_ ),
    .B(\dec/_225_ ),
    .X(\dec/_226_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_493_  (.A(\dec/_226_ ),
    .X(\dec/_227_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_494_  (.A(\dec/_227_ ),
    .B(\dec/_218_ ),
    .Y(\dec/_228_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_495_  (.A(\dec/_222_ ),
    .B(\dec/_223_ ),
    .C(\dec/_228_ ),
    .Y(\dec/_229_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_496_  (.A(\dec/_219_ ),
    .B(\dec/_229_ ),
    .C(\dec/_072_ ),
    .Y(\dec/_230_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_497_  (.A(net261),
    .B(net2191),
    .Y(\dec/_231_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_498_  (.A(\dec/_230_ ),
    .B(\dec/_231_ ),
    .Y(\dec/_016_ ));
 sky130_fd_sc_hd__o21bai_1 \dec/_499_  (.A1(\dec/_187_ ),
    .A2(\dec/_197_ ),
    .B1_N(\dec/_075_ ),
    .Y(\dec/_232_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_500_  (.A(\dec/_227_ ),
    .B(\dec/_205_ ),
    .Y(\dec/_233_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_501_  (.A(\dec/_222_ ),
    .B(\dec/_223_ ),
    .C(\dec/_233_ ),
    .Y(\dec/_234_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_502_  (.A(\dec/_232_ ),
    .B(\dec/_234_ ),
    .C(\dec/_072_ ),
    .Y(\dec/_235_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_503_  (.A(net244),
    .B(net2221),
    .Y(\dec/_236_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_504_  (.A(\dec/_235_ ),
    .B(\dec/_236_ ),
    .Y(\dec/_017_ ));
 sky130_fd_sc_hd__o21bai_1 \dec/_505_  (.A1(\dec/_187_ ),
    .A2(\dec/_197_ ),
    .B1_N(\dec/_079_ ),
    .Y(\dec/_237_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_506_  (.A(\dec/_227_ ),
    .B(\dec/_208_ ),
    .Y(\dec/_238_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_507_  (.A(\dec/_222_ ),
    .B(\dec/_223_ ),
    .C(\dec/_238_ ),
    .Y(\dec/_239_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_508_  (.A(\dec/_237_ ),
    .B(\dec/_239_ ),
    .C(\dec/_072_ ),
    .Y(\dec/_240_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_509_  (.A(net244),
    .B(\imm12_i_s[2] ),
    .Y(\dec/_241_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_510_  (.A(\dec/_240_ ),
    .B(\dec/_241_ ),
    .Y(\dec/_018_ ));
 sky130_fd_sc_hd__o21bai_1 \dec/_511_  (.A1(\dec/_187_ ),
    .A2(\dec/_197_ ),
    .B1_N(\dec/_082_ ),
    .Y(\dec/_242_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_512_  (.A(\dec/_227_ ),
    .B(\dec/_212_ ),
    .Y(\dec/_243_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_513_  (.A(\dec/_222_ ),
    .B(\dec/_223_ ),
    .C(\dec/_243_ ),
    .Y(\dec/_244_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_514_  (.A(\dec/_242_ ),
    .B(\dec/_244_ ),
    .C(\dec/_072_ ),
    .Y(\dec/_245_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_515_  (.A(net244),
    .B(\imm12_i_s[3] ),
    .Y(\dec/_246_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_516_  (.A(\dec/_245_ ),
    .B(\dec/_246_ ),
    .Y(\dec/_019_ ));
 sky130_fd_sc_hd__o21bai_1 \dec/_517_  (.A1(\dec/_187_ ),
    .A2(\dec/_197_ ),
    .B1_N(\dec/_085_ ),
    .Y(\dec/_247_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_518_  (.A(\dec/_227_ ),
    .B(\dec/_215_ ),
    .Y(\dec/_248_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_519_  (.A(\dec/_222_ ),
    .B(\dec/_223_ ),
    .C(\dec/_248_ ),
    .Y(\dec/_249_ ));
 sky130_fd_sc_hd__nand3_1 \dec/_520_  (.A(\dec/_247_ ),
    .B(\dec/_249_ ),
    .C(\dec/_072_ ),
    .Y(\dec/_250_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_521_  (.A(net260),
    .B(net2211),
    .Y(\dec/_251_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_522_  (.A(\dec/_250_ ),
    .B(\dec/_251_ ),
    .Y(\dec/_020_ ));
 sky130_fd_sc_hd__nand3b_2 \dec/_523_  (.A_N(\dec/_226_ ),
    .B(\dec/_222_ ),
    .C(\dec/_223_ ),
    .Y(\dec/_252_ ));
 sky130_fd_sc_hd__buf_6 \dec/_524_  (.A(\dec/_252_ ),
    .X(\dec/_253_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \dec/_525_  (.A(\dec/_062_ ),
    .X(\dec/_254_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_526_  (.A(\dec/_097_ ),
    .X(\dec/_255_ ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_527_  (.A(\dec/_089_ ),
    .X(\dec/_256_ ));
 sky130_fd_sc_hd__a221o_1 \dec/_528_  (.A1(net893),
    .A2(\dec/rInstrustion2[25] ),
    .B1(\dec/_256_ ),
    .B2(net51),
    .C1(net884),
    .X(\dec/_257_ ));
 sky130_fd_sc_hd__o211a_2 \dec/_529_  (.A1(\dec/_254_ ),
    .A2(\dec/rInstrustion1[25] ),
    .B1(\dec/_255_ ),
    .C1(\dec/_257_ ),
    .X(\dec/_258_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_530_  (.A(\dec/_253_ ),
    .B(\dec/_258_ ),
    .Y(\dec/_259_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_531_  (.A(net267),
    .B(net2135),
    .Y(\dec/_260_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_532_  (.A(\dec/_259_ ),
    .B(\dec/_260_ ),
    .Y(\dec/_021_ ));
 sky130_fd_sc_hd__a221o_1 \dec/_533_  (.A1(net893),
    .A2(\dec/rInstrustion2[26] ),
    .B1(\dec/_256_ ),
    .B2(net52),
    .C1(net885),
    .X(\dec/_261_ ));
 sky130_fd_sc_hd__o211a_2 \dec/_534_  (.A1(\dec/_254_ ),
    .A2(\dec/rInstrustion1[26] ),
    .B1(\dec/_255_ ),
    .C1(\dec/_261_ ),
    .X(\dec/_262_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_535_  (.A(\dec/_253_ ),
    .B(\dec/_262_ ),
    .Y(\dec/_263_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_536_  (.A(net266),
    .B(\imm12_i_s[6] ),
    .Y(\dec/_264_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_537_  (.A(\dec/_263_ ),
    .B(\dec/_264_ ),
    .Y(\dec/_022_ ));
 sky130_fd_sc_hd__a221o_1 \dec/_538_  (.A1(net892),
    .A2(\dec/rInstrustion2[27] ),
    .B1(\dec/_256_ ),
    .B2(net53),
    .C1(net884),
    .X(\dec/_265_ ));
 sky130_fd_sc_hd__o211a_2 \dec/_539_  (.A1(\dec/_254_ ),
    .A2(\dec/rInstrustion1[27] ),
    .B1(\dec/_255_ ),
    .C1(\dec/_265_ ),
    .X(\dec/_266_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_540_  (.A(\dec/_253_ ),
    .B(\dec/_266_ ),
    .Y(\dec/_267_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_541_  (.A(net265),
    .B(net2142),
    .Y(\dec/_268_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_542_  (.A(\dec/_267_ ),
    .B(\dec/_268_ ),
    .Y(\dec/_023_ ));
 sky130_fd_sc_hd__a221o_1 \dec/_543_  (.A1(net893),
    .A2(\dec/rInstrustion2[28] ),
    .B1(\dec/_256_ ),
    .B2(net54),
    .C1(net885),
    .X(\dec/_269_ ));
 sky130_fd_sc_hd__o211a_2 \dec/_544_  (.A1(\dec/_254_ ),
    .A2(\dec/rInstrustion1[28] ),
    .B1(\dec/_255_ ),
    .C1(\dec/_269_ ),
    .X(\dec/_270_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_545_  (.A(\dec/_253_ ),
    .B(\dec/_270_ ),
    .Y(\dec/_271_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_546_  (.A(net266),
    .B(\imm12_i_s[8] ),
    .Y(\dec/_272_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_547_  (.A(\dec/_271_ ),
    .B(\dec/_272_ ),
    .Y(\dec/_024_ ));
 sky130_fd_sc_hd__a221o_1 \dec/_548_  (.A1(net893),
    .A2(\dec/rInstrustion2[29] ),
    .B1(\dec/_256_ ),
    .B2(net55),
    .C1(net885),
    .X(\dec/_273_ ));
 sky130_fd_sc_hd__o211a_2 \dec/_549_  (.A1(\dec/_254_ ),
    .A2(\dec/rInstrustion1[29] ),
    .B1(\dec/_255_ ),
    .C1(\dec/_273_ ),
    .X(\dec/_274_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_550_  (.A(\dec/_253_ ),
    .B(\dec/_274_ ),
    .Y(\dec/_275_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_551_  (.A(net267),
    .B(net2098),
    .Y(\dec/_276_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_552_  (.A(\dec/_275_ ),
    .B(\dec/_276_ ),
    .Y(\dec/_025_ ));
 sky130_fd_sc_hd__a221o_1 \dec/_553_  (.A1(net892),
    .A2(\dec/rInstrustion2[30] ),
    .B1(\dec/_256_ ),
    .B2(net57),
    .C1(net884),
    .X(\dec/_277_ ));
 sky130_fd_sc_hd__o211a_2 \dec/_554_  (.A1(\dec/_254_ ),
    .A2(\dec/rInstrustion1[30] ),
    .B1(\dec/_098_ ),
    .C1(\dec/_277_ ),
    .X(\dec/_278_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_555_  (.A(\dec/_253_ ),
    .B(\dec/_278_ ),
    .Y(\dec/_279_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_556_  (.A(net265),
    .B(net2106),
    .Y(\dec/_280_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_557_  (.A(\dec/_279_ ),
    .B(\dec/_280_ ),
    .Y(\dec/_026_ ));
 sky130_fd_sc_hd__a221o_1 \dec/_558_  (.A1(net892),
    .A2(\dec/rInstrustion2[31] ),
    .B1(\dec/_090_ ),
    .B2(net58),
    .C1(net884),
    .X(\dec/_281_ ));
 sky130_fd_sc_hd__o211a_2 \dec/_559_  (.A1(\dec/_094_ ),
    .A2(\dec/rInstrustion1[31] ),
    .B1(\dec/_098_ ),
    .C1(\dec/_281_ ),
    .X(\dec/_282_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_560_  (.A(\dec/_252_ ),
    .B(\dec/_282_ ),
    .Y(\dec/_283_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_561_  (.A(net263),
    .B(net2165),
    .Y(\dec/_284_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_562_  (.A(\dec/_283_ ),
    .B(\dec/_284_ ),
    .Y(\dec/_027_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_563_  (.A1(net261),
    .A2(\imm21_j[1] ),
    .B1(\dec/_075_ ),
    .B2(\dec/_209_ ),
    .X(\dec/_028_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_564_  (.A1(net261),
    .A2(net1152),
    .B1(\dec/_079_ ),
    .B2(\dec/_209_ ),
    .X(\dec/_029_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_565_  (.A1(net261),
    .A2(net1162),
    .B1(\dec/_082_ ),
    .B2(\dec/_200_ ),
    .X(\dec/_030_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_566_  (.A1(net261),
    .A2(\imm21_j[4] ),
    .B1(\dec/_085_ ),
    .B2(\dec/_200_ ),
    .X(\dec/_031_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_567_  (.A1(net265),
    .A2(net1981),
    .B1(\dec/_258_ ),
    .X(\dec/_032_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_568_  (.A1(net265),
    .A2(\funct7[1] ),
    .B1(\dec/_262_ ),
    .X(\dec/_033_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_569_  (.A1(net265),
    .A2(\funct7[2] ),
    .B1(\dec/_266_ ),
    .X(\dec/_034_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_570_  (.A1(net268),
    .A2(net1866),
    .B1(\dec/_270_ ),
    .X(\dec/_035_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_571_  (.A1(net265),
    .A2(net2073),
    .B1(\dec/_274_ ),
    .X(\dec/_036_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_572_  (.A1(net263),
    .A2(net2053),
    .B1(\dec/_278_ ),
    .X(\dec/_037_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_573_  (.A1(net248),
    .A2(net1138),
    .B1(\dec/_069_ ),
    .B2(\dec/_200_ ),
    .X(\dec/_038_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_574_  (.A(wJumping),
    .B(\dec/_095_ ),
    .Y(\dec/_285_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_575_  (.A1(net894),
    .A2(\dec/rInstrustion2[12] ),
    .B1(net887),
    .X(\dec/_286_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_576_  (.A1(net37),
    .A2(\dec/_089_ ),
    .B1(\dec/_286_ ),
    .X(\dec/_287_ ));
 sky130_fd_sc_hd__o211ai_2 \dec/_577_  (.A1(\dec/_062_ ),
    .A2(\dec/rInstrustion1[12] ),
    .B1(\dec/_285_ ),
    .C1(\dec/_287_ ),
    .Y(\dec/_288_ ));
 sky130_fd_sc_hd__or2_1 \dec/_578_  (.A(net247),
    .B(\dec/_288_ ),
    .X(\dec/_289_ ));
 sky130_fd_sc_hd__a21bo_1 \dec/_579_  (.A1(net247),
    .A2(\imm21_j[12] ),
    .B1_N(\dec/_289_ ),
    .X(\dec/_039_ ));
 sky130_fd_sc_hd__o21ai_1 \dec/_580_  (.A1(\dec/_062_ ),
    .A2(\dec/rInstrustion1[13] ),
    .B1(\dec/_285_ ),
    .Y(\dec/_290_ ));
 sky130_fd_sc_hd__a221oi_1 \dec/_581_  (.A1(net892),
    .A2(\dec/rInstrustion2[13] ),
    .B1(\dec/_089_ ),
    .B2(net38),
    .C1(net884),
    .Y(\dec/_291_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_582_  (.A(\dec/_290_ ),
    .B(\dec/_291_ ),
    .Y(\dec/_292_ ));
 sky130_fd_sc_hd__or2b_1 \dec/_583_  (.A(net248),
    .B_N(\dec/_292_ ),
    .X(\dec/_293_ ));
 sky130_fd_sc_hd__a21bo_1 \dec/_584_  (.A1(net264),
    .A2(net2226),
    .B1_N(\dec/_293_ ),
    .X(\dec/_040_ ));
 sky130_fd_sc_hd__a221o_1 \dec/_585_  (.A1(\dec/rInstrustion2[14] ),
    .A2(net893),
    .B1(\dec/_091_ ),
    .B2(net39),
    .C1(net884),
    .X(\dec/_294_ ));
 sky130_fd_sc_hd__o21a_1 \dec/_586_  (.A1(\dec/rInstrustion1[14] ),
    .A2(\dec/_087_ ),
    .B1(\dec/_255_ ),
    .X(\dec/_295_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_587_  (.A1(net241),
    .A2(net1157),
    .B1(\dec/_294_ ),
    .B2(\dec/_295_ ),
    .X(\dec/_041_ ));
 sky130_fd_sc_hd__a21bo_1 \dec/_588_  (.A1(net249),
    .A2(net1134),
    .B1_N(\dec/_100_ ),
    .X(\dec/_042_ ));
 sky130_fd_sc_hd__a21bo_1 \dec/_589_  (.A1(net246),
    .A2(net1153),
    .B1_N(\dec/_104_ ),
    .X(\dec/_043_ ));
 sky130_fd_sc_hd__a21bo_1 \dec/_590_  (.A1(net247),
    .A2(net1149),
    .B1_N(\dec/_108_ ),
    .X(\dec/_044_ ));
 sky130_fd_sc_hd__a21bo_1 \dec/_591_  (.A1(net241),
    .A2(net1141),
    .B1_N(\dec/_112_ ),
    .X(\dec/_045_ ));
 sky130_fd_sc_hd__a21bo_1 \dec/_592_  (.A1(net239),
    .A2(net1148),
    .B1_N(\dec/_116_ ),
    .X(\dec/_046_ ));
 sky130_fd_sc_hd__a21o_1 \dec/_593_  (.A1(net251),
    .A2(\funct7[6] ),
    .B1(\dec/_282_ ),
    .X(\dec/_047_ ));
 sky130_fd_sc_hd__a32o_1 \dec/_594_  (.A1(\dec/_184_ ),
    .A2(\dec/_199_ ),
    .A3(\dec/_200_ ),
    .B1(net246),
    .B2(net2151),
    .X(\dec/_048_ ));
 sky130_fd_sc_hd__a32o_1 \dec/_595_  (.A1(\dec/_184_ ),
    .A2(\dec/_194_ ),
    .A3(\dec/_071_ ),
    .B1(net246),
    .B2(net921),
    .X(\dec/_049_ ));
 sky130_fd_sc_hd__a21bo_1 \dec/_596_  (.A1(net248),
    .A2(net2179),
    .B1_N(\dec/_289_ ),
    .X(\dec/_050_ ));
 sky130_fd_sc_hd__a21bo_1 \dec/_597_  (.A1(net273),
    .A2(net2146),
    .B1_N(\dec/_293_ ),
    .X(\dec/_051_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_598_  (.A1(net241),
    .A2(net67),
    .B1(\dec/_294_ ),
    .B2(\dec/_295_ ),
    .X(\dec/_052_ ));
 sky130_fd_sc_hd__a2bb2o_1 \dec/_599_  (.A1_N(\dec/_096_ ),
    .A2_N(\dec/_185_ ),
    .B1(net238),
    .B2(net898),
    .X(\dec/_053_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_600_  (.A(\dec/_189_ ),
    .B(\dec/_071_ ),
    .Y(\dec/_296_ ));
 sky130_fd_sc_hd__a2bb2o_1 \dec/_601_  (.A1_N(\dec/_162_ ),
    .A2_N(\dec/_296_ ),
    .B1(net246),
    .B2(net897),
    .X(\dec/_054_ ));
 sky130_fd_sc_hd__a2bb2o_1 \dec/_602_  (.A1_N(\dec/_096_ ),
    .A2_N(\dec/_196_ ),
    .B1(net245),
    .B2(op_memLd),
    .X(\dec/_055_ ));
 sky130_fd_sc_hd__inv_2 \dec/_603_  (.A(\dec/_194_ ),
    .Y(\dec/_297_ ));
 sky130_fd_sc_hd__nor2_1 \dec/_604_  (.A(\dec/_288_ ),
    .B(\dec/_292_ ),
    .Y(\dec/_298_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_605_  (.A(net247),
    .B(net1557),
    .Y(\dec/_299_ ));
 sky130_fd_sc_hd__o31ai_1 \dec/_606_  (.A1(\dec/_297_ ),
    .A2(\dec/_296_ ),
    .A3(\dec/_298_ ),
    .B1(\dec/_299_ ),
    .Y(\dec/_056_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_607_  (.A1(net247),
    .A2(net2181),
    .B1(\dec/_227_ ),
    .B2(\dec/_200_ ),
    .X(\dec/_057_ ));
 sky130_fd_sc_hd__nand2_1 \dec/_608_  (.A(net247),
    .B(net2042),
    .Y(\dec/_300_ ));
 sky130_fd_sc_hd__o31ai_1 \dec/_609_  (.A1(\dec/_195_ ),
    .A2(\dec/_292_ ),
    .A3(\dec/_289_ ),
    .B1(\dec/_300_ ),
    .Y(\dec/_058_ ));
 sky130_fd_sc_hd__a22o_1 \dec/_610_  (.A1(net238),
    .A2(net1178),
    .B1(\dec/_145_ ),
    .B2(\dec/_179_ ),
    .X(\dec/_059_ ));
 sky130_fd_sc_hd__a2bb2o_1 \dec/_611_  (.A1_N(\dec/_096_ ),
    .A2_N(\dec/_192_ ),
    .B1(net246),
    .B2(net1168),
    .X(\dec/_060_ ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_612_  (.CLK(clknet_leaf_25_clk),
    .D(\dec/_000_ ),
    .Q(j_type));
 sky130_fd_sc_hd__dfxtp_1 \dec/_613_  (.CLK(clknet_leaf_24_clk),
    .D(\dec/_001_ ),
    .Q(\Op_code[0] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_614_  (.CLK(clknet_leaf_24_clk),
    .D(\dec/_002_ ),
    .Q(\Op_code[1] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_615_  (.CLK(clknet_leaf_27_clk),
    .D(\dec/_003_ ),
    .Q(\Op_code[2] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_616_  (.CLK(clknet_leaf_24_clk),
    .D(\dec/_004_ ),
    .Q(\Op_code[3] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_617_  (.CLK(clknet_leaf_26_clk),
    .D(\dec/_005_ ),
    .Q(\Op_code[4] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_618_  (.CLK(clknet_leaf_26_clk),
    .D(\dec/_006_ ),
    .Q(\Op_code[5] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_619_  (.CLK(clknet_leaf_25_clk),
    .D(\dec/_007_ ),
    .Q(\Op_code[6] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_620_  (.CLK(clknet_leaf_24_clk),
    .D(\dec/_008_ ),
    .Q(i_type));
 sky130_fd_sc_hd__dfxtp_2 \dec/_621_  (.CLK(clknet_leaf_24_clk),
    .D(\dec/_009_ ),
    .Q(op_intRegReg));
 sky130_fd_sc_hd__dfxtp_1 \dec/_622_  (.CLK(clknet_leaf_27_clk),
    .D(\dec/_010_ ),
    .Q(u_type));
 sky130_fd_sc_hd__dfxtp_1 \dec/_623_  (.CLK(clknet_leaf_23_clk),
    .D(\wReg_s1_out[0] ),
    .Q(\reg_s1[0] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_624_  (.CLK(clknet_leaf_20_clk),
    .D(\wReg_s1_out[1] ),
    .Q(\reg_s1[1] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_625_  (.CLK(clknet_leaf_20_clk),
    .D(\wReg_s1_out[2] ),
    .Q(\reg_s1[2] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_626_  (.CLK(clknet_leaf_20_clk),
    .D(\wReg_s1_out[3] ),
    .Q(\reg_s1[3] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_627_  (.CLK(clknet_leaf_63_clk),
    .D(\wReg_s1_out[4] ),
    .Q(\reg_s1[4] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_628_  (.CLK(clknet_leaf_23_clk),
    .D(\wReg_s2_out[0] ),
    .Q(\reg_s2[0] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_629_  (.CLK(clknet_leaf_64_clk),
    .D(\wReg_s2_out[1] ),
    .Q(\reg_s2[1] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_630_  (.CLK(clknet_leaf_19_clk),
    .D(\wReg_s2_out[2] ),
    .Q(\reg_s2[2] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_631_  (.CLK(clknet_leaf_64_clk),
    .D(\wReg_s2_out[3] ),
    .Q(\reg_s2[3] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_632_  (.CLK(clknet_leaf_64_clk),
    .D(\wReg_s2_out[4] ),
    .Q(\reg_s2[4] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_633_  (.CLK(clknet_leaf_24_clk),
    .D(\dec/_011_ ),
    .Q(\imm13_b[1] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_634_  (.CLK(clknet_leaf_20_clk),
    .D(\dec/_012_ ),
    .Q(\imm13_b[2] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_635_  (.CLK(clknet_leaf_45_clk),
    .D(\dec/_013_ ),
    .Q(\imm13_b[3] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_636_  (.CLK(clknet_leaf_23_clk),
    .D(\dec/_014_ ),
    .Q(\imm13_b[4] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_637_  (.CLK(clknet_leaf_45_clk),
    .D(\dec/_015_ ),
    .Q(\imm13_b[11] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_638_  (.CLK(clknet_leaf_45_clk),
    .D(\dec/_016_ ),
    .Q(\imm12_i_s[0] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_639_  (.CLK(clknet_leaf_44_clk),
    .D(\dec/_017_ ),
    .Q(\imm12_i_s[1] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_640_  (.CLK(clknet_leaf_44_clk),
    .D(\dec/_018_ ),
    .Q(\imm12_i_s[2] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_641_  (.CLK(clknet_leaf_44_clk),
    .D(\dec/_019_ ),
    .Q(\imm12_i_s[3] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_642_  (.CLK(clknet_leaf_63_clk),
    .D(\dec/_020_ ),
    .Q(\imm12_i_s[4] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_643_  (.CLK(clknet_leaf_60_clk),
    .D(\dec/_021_ ),
    .Q(\imm12_i_s[5] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_644_  (.CLK(clknet_leaf_57_clk),
    .D(\dec/_022_ ),
    .Q(\imm12_i_s[6] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_645_  (.CLK(clknet_leaf_60_clk),
    .D(\dec/_023_ ),
    .Q(\imm12_i_s[7] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_646_  (.CLK(clknet_leaf_57_clk),
    .D(\dec/_024_ ),
    .Q(\imm12_i_s[8] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_647_  (.CLK(clknet_leaf_61_clk),
    .D(\dec/_025_ ),
    .Q(\imm12_i_s[9] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_648_  (.CLK(clknet_leaf_60_clk),
    .D(\dec/_026_ ),
    .Q(\imm12_i_s[10] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_649_  (.CLK(clknet_leaf_45_clk),
    .D(\dec/_027_ ),
    .Q(\imm12_i_s[11] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_650_  (.CLK(clknet_leaf_63_clk),
    .D(\dec/_028_ ),
    .Q(\imm21_j[1] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_651_  (.CLK(clknet_leaf_63_clk),
    .D(\dec/_029_ ),
    .Q(\imm21_j[2] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_652_  (.CLK(clknet_leaf_63_clk),
    .D(\dec/_030_ ),
    .Q(\imm21_j[3] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_653_  (.CLK(clknet_leaf_63_clk),
    .D(\dec/_031_ ),
    .Q(\imm21_j[4] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_654_  (.CLK(clknet_leaf_62_clk),
    .D(\dec/_032_ ),
    .Q(\funct7[0] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_655_  (.CLK(clknet_leaf_61_clk),
    .D(\dec/_033_ ),
    .Q(\funct7[1] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_656_  (.CLK(clknet_leaf_61_clk),
    .D(\dec/_034_ ),
    .Q(\funct7[2] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_657_  (.CLK(clknet_leaf_61_clk),
    .D(\dec/_035_ ),
    .Q(\funct7[3] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_658_  (.CLK(clknet_leaf_60_clk),
    .D(\dec/_036_ ),
    .Q(\funct7[4] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_659_  (.CLK(clknet_leaf_45_clk),
    .D(\dec/_037_ ),
    .Q(\funct7[5] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_660_  (.CLK(clknet_leaf_45_clk),
    .D(\dec/_038_ ),
    .Q(\imm21_j[11] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_661_  (.CLK(clknet_leaf_43_clk),
    .D(\dec/_039_ ),
    .Q(\imm21_j[12] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_662_  (.CLK(clknet_leaf_62_clk),
    .D(\dec/_040_ ),
    .Q(\imm21_j[13] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_663_  (.CLK(clknet_leaf_31_clk),
    .D(\dec/_041_ ),
    .Q(\imm21_j[14] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_664_  (.CLK(clknet_leaf_25_clk),
    .D(\dec/_042_ ),
    .Q(\imm21_j[15] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_665_  (.CLK(clknet_leaf_44_clk),
    .D(\dec/_043_ ),
    .Q(\imm21_j[16] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_666_  (.CLK(clknet_leaf_44_clk),
    .D(\dec/_044_ ),
    .Q(\imm21_j[17] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_667_  (.CLK(clknet_leaf_31_clk),
    .D(\dec/_045_ ),
    .Q(\imm21_j[18] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_668_  (.CLK(clknet_leaf_26_clk),
    .D(\dec/_046_ ),
    .Q(\imm21_j[19] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_669_  (.CLK(clknet_leaf_31_clk),
    .D(\dec/_047_ ),
    .Q(\funct7[6] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_670_  (.CLK(clknet_leaf_24_clk),
    .D(\dec/_048_ ),
    .Q(op_lui));
 sky130_fd_sc_hd__dfxtp_1 \dec/_671_  (.CLK(clknet_leaf_25_clk),
    .D(\dec/_049_ ),
    .Q(op_auipc));
 sky130_fd_sc_hd__dfxtp_2 \dec/_672_  (.CLK(clknet_leaf_43_clk),
    .D(\dec/_050_ ),
    .Q(\funct3[0] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_673_  (.CLK(clknet_leaf_51_clk),
    .D(\dec/_051_ ),
    .Q(\funct3[1] ));
 sky130_fd_sc_hd__dfxtp_2 \dec/_674_  (.CLK(clknet_leaf_31_clk),
    .D(\dec/_052_ ),
    .Q(net67));
 sky130_fd_sc_hd__dfxtp_1 \dec/_675_  (.CLK(clknet_leaf_25_clk),
    .D(\dec/_053_ ),
    .Q(op_jalr));
 sky130_fd_sc_hd__dfxtp_1 \dec/_676_  (.CLK(clknet_4_4__leaf_clk),
    .D(\dec/_054_ ),
    .Q(b_type));
 sky130_fd_sc_hd__dfxtp_2 \dec/_677_  (.CLK(clknet_leaf_24_clk),
    .D(\dec/_055_ ),
    .Q(op_memLd));
 sky130_fd_sc_hd__dfxtp_1 \dec/_678_  (.CLK(clknet_leaf_44_clk),
    .D(\dec/_056_ ),
    .Q(op_intRegImm));
 sky130_fd_sc_hd__dfxtp_2 \dec/_679_  (.CLK(clknet_leaf_44_clk),
    .D(\dec/_057_ ),
    .Q(op_memSt));
 sky130_fd_sc_hd__dfxtp_2 \dec/_680_  (.CLK(clknet_leaf_44_clk),
    .D(\dec/_058_ ),
    .Q(op_consShf));
 sky130_fd_sc_hd__dfxtp_1 \dec/_681_  (.CLK(clknet_leaf_24_clk),
    .D(\dec/_059_ ),
    .Q(op_efence));
 sky130_fd_sc_hd__dfxtp_1 \dec/_682_  (.CLK(clknet_leaf_24_clk),
    .D(\dec/_060_ ),
    .Q(op_ecb));
 sky130_fd_sc_hd__dfxtp_1 \dec/_683_  (.CLK(clknet_leaf_31_clk),
    .D(net886),
    .Q(\dec/rStall2 ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_684_  (.CLK(clknet_leaf_22_clk),
    .D(net34),
    .Q(\dec/rInstrustion1[0] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_685_  (.CLK(clknet_leaf_27_clk),
    .D(net45),
    .Q(\dec/rInstrustion1[1] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_686_  (.CLK(clknet_leaf_27_clk),
    .D(net56),
    .Q(\dec/rInstrustion1[2] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_687_  (.CLK(clknet_leaf_28_clk),
    .D(net59),
    .Q(\dec/rInstrustion1[3] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_688_  (.CLK(clknet_leaf_27_clk),
    .D(net60),
    .Q(\dec/rInstrustion1[4] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_689_  (.CLK(clknet_leaf_31_clk),
    .D(net61),
    .Q(\dec/rInstrustion1[5] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_690_  (.CLK(clknet_leaf_27_clk),
    .D(net62),
    .Q(\dec/rInstrustion1[6] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_691_  (.CLK(clknet_leaf_28_clk),
    .D(net63),
    .Q(\dec/rInstrustion1[7] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_692_  (.CLK(clknet_leaf_28_clk),
    .D(net64),
    .Q(\dec/rInstrustion1[8] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_693_  (.CLK(clknet_leaf_21_clk),
    .D(net65),
    .Q(\dec/rInstrustion1[9] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_694_  (.CLK(clknet_leaf_21_clk),
    .D(net35),
    .Q(\dec/rInstrustion1[10] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_695_  (.CLK(clknet_leaf_21_clk),
    .D(net36),
    .Q(\dec/rInstrustion1[11] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_696_  (.CLK(clknet_leaf_29_clk),
    .D(net37),
    .Q(\dec/rInstrustion1[12] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_697_  (.CLK(clknet_leaf_29_clk),
    .D(net38),
    .Q(\dec/rInstrustion1[13] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_698_  (.CLK(clknet_leaf_30_clk),
    .D(net39),
    .Q(\dec/rInstrustion1[14] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_699_  (.CLK(clknet_leaf_29_clk),
    .D(net40),
    .Q(\dec/rInstrustion1[15] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_700_  (.CLK(clknet_leaf_28_clk),
    .D(net41),
    .Q(\dec/rInstrustion1[16] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_701_  (.CLK(clknet_leaf_29_clk),
    .D(net42),
    .Q(\dec/rInstrustion1[17] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_702_  (.CLK(clknet_leaf_28_clk),
    .D(net43),
    .Q(\dec/rInstrustion1[18] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_703_  (.CLK(clknet_leaf_30_clk),
    .D(net44),
    .Q(\dec/rInstrustion1[19] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_704_  (.CLK(clknet_leaf_21_clk),
    .D(net46),
    .Q(\dec/rInstrustion1[20] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_705_  (.CLK(clknet_leaf_22_clk),
    .D(net47),
    .Q(\dec/rInstrustion1[21] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_706_  (.CLK(clknet_leaf_22_clk),
    .D(net48),
    .Q(\dec/rInstrustion1[22] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_707_  (.CLK(clknet_leaf_22_clk),
    .D(net49),
    .Q(\dec/rInstrustion1[23] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_708_  (.CLK(clknet_leaf_21_clk),
    .D(net50),
    .Q(\dec/rInstrustion1[24] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_709_  (.CLK(clknet_leaf_29_clk),
    .D(net51),
    .Q(\dec/rInstrustion1[25] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_710_  (.CLK(clknet_leaf_29_clk),
    .D(net52),
    .Q(\dec/rInstrustion1[26] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_711_  (.CLK(clknet_leaf_29_clk),
    .D(net53),
    .Q(\dec/rInstrustion1[27] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_712_  (.CLK(clknet_leaf_30_clk),
    .D(net54),
    .Q(\dec/rInstrustion1[28] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_713_  (.CLK(clknet_leaf_30_clk),
    .D(net55),
    .Q(\dec/rInstrustion1[29] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_714_  (.CLK(clknet_leaf_29_clk),
    .D(net57),
    .Q(\dec/rInstrustion1[30] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_715_  (.CLK(clknet_leaf_28_clk),
    .D(net58),
    .Q(\dec/rInstrustion1[31] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_716_  (.CLK(clknet_leaf_22_clk),
    .D(net1107),
    .Q(\dec/rInstrustion2[0] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_717_  (.CLK(clknet_leaf_27_clk),
    .D(net1115),
    .Q(\dec/rInstrustion2[1] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_718_  (.CLK(clknet_leaf_27_clk),
    .D(net1116),
    .Q(\dec/rInstrustion2[2] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_719_  (.CLK(clknet_leaf_27_clk),
    .D(net1112),
    .Q(\dec/rInstrustion2[3] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_720_  (.CLK(clknet_leaf_27_clk),
    .D(net1128),
    .Q(\dec/rInstrustion2[4] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_721_  (.CLK(clknet_leaf_26_clk),
    .D(net1104),
    .Q(\dec/rInstrustion2[5] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_722_  (.CLK(clknet_leaf_27_clk),
    .D(net1124),
    .Q(\dec/rInstrustion2[6] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_723_  (.CLK(clknet_leaf_28_clk),
    .D(net1130),
    .Q(\dec/rInstrustion2[7] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_724_  (.CLK(clknet_leaf_28_clk),
    .D(net1106),
    .Q(\dec/rInstrustion2[8] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_725_  (.CLK(clknet_leaf_21_clk),
    .D(net1117),
    .Q(\dec/rInstrustion2[9] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_726_  (.CLK(clknet_leaf_28_clk),
    .D(net1125),
    .Q(\dec/rInstrustion2[10] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_727_  (.CLK(clknet_leaf_21_clk),
    .D(net1110),
    .Q(\dec/rInstrustion2[11] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_728_  (.CLK(clknet_leaf_31_clk),
    .D(net1143),
    .Q(\dec/rInstrustion2[12] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_729_  (.CLK(clknet_leaf_29_clk),
    .D(net1126),
    .Q(\dec/rInstrustion2[13] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_730_  (.CLK(clknet_leaf_30_clk),
    .D(net1103),
    .Q(\dec/rInstrustion2[14] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_731_  (.CLK(clknet_leaf_29_clk),
    .D(net1131),
    .Q(\dec/rInstrustion2[15] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_732_  (.CLK(clknet_leaf_27_clk),
    .D(net1101),
    .Q(\dec/rInstrustion2[16] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_733_  (.CLK(clknet_leaf_29_clk),
    .D(net1123),
    .Q(\dec/rInstrustion2[17] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_734_  (.CLK(clknet_leaf_28_clk),
    .D(net1118),
    .Q(\dec/rInstrustion2[18] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_735_  (.CLK(clknet_leaf_30_clk),
    .D(net1102),
    .Q(\dec/rInstrustion2[19] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_736_  (.CLK(clknet_leaf_22_clk),
    .D(net1119),
    .Q(\dec/rInstrustion2[20] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_737_  (.CLK(clknet_leaf_22_clk),
    .D(net1111),
    .Q(\dec/rInstrustion2[21] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_738_  (.CLK(clknet_leaf_22_clk),
    .D(net1108),
    .Q(\dec/rInstrustion2[22] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_739_  (.CLK(clknet_leaf_22_clk),
    .D(net1105),
    .Q(\dec/rInstrustion2[23] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_740_  (.CLK(clknet_leaf_21_clk),
    .D(net1121),
    .Q(\dec/rInstrustion2[24] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_741_  (.CLK(clknet_leaf_29_clk),
    .D(net1132),
    .Q(\dec/rInstrustion2[25] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_742_  (.CLK(clknet_leaf_29_clk),
    .D(net1122),
    .Q(\dec/rInstrustion2[26] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_743_  (.CLK(clknet_leaf_29_clk),
    .D(net1129),
    .Q(\dec/rInstrustion2[27] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_744_  (.CLK(clknet_leaf_30_clk),
    .D(net1109),
    .Q(\dec/rInstrustion2[28] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_745_  (.CLK(clknet_leaf_30_clk),
    .D(net1113),
    .Q(\dec/rInstrustion2[29] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_746_  (.CLK(clknet_leaf_29_clk),
    .D(net1127),
    .Q(\dec/rInstrustion2[30] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_747_  (.CLK(clknet_leaf_28_clk),
    .D(net1120),
    .Q(\dec/rInstrustion2[31] ));
 sky130_fd_sc_hd__dfxtp_1 \dec/_748_  (.CLK(clknet_leaf_31_clk),
    .D(net241),
    .Q(\dec/rStall1 ));
 sky130_fd_sc_hd__conb_1 \brancher/_2116__1075  (.LO(net1075));
 sky130_fd_sc_hd__conb_1 _1722__1076 (.LO(net1076));
 sky130_fd_sc_hd__conb_1 _1731__1078 (.LO(net1078));
 sky130_fd_sc_hd__conb_1 _1737__1080 (.LO(net1080));
 sky130_fd_sc_hd__conb_1 _1741__1082 (.LO(net1082));
 sky130_fd_sc_hd__conb_1 _1745__1084 (.LO(net1084));
 sky130_fd_sc_hd__conb_1 _1750__1086 (.LO(net1086));
 sky130_fd_sc_hd__conb_1 _1755__1088 (.LO(net1088));
 sky130_fd_sc_hd__conb_1 _1759__1090 (.LO(net1090));
 sky130_fd_sc_hd__conb_1 _1765__1092 (.LO(net1092));
 sky130_fd_sc_hd__conb_1 _1769__1094 (.LO(net1094));
 sky130_fd_sc_hd__conb_1 _1773__1096 (.LO(net1096));
 sky130_fd_sc_hd__conb_1 _1778__1098 (.LO(net1098));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkbuf_1 \dec/_763_  (.A(net1981),
    .X(\imm13_b[5] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_764_  (.A(net2069),
    .X(\imm13_b[6] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_765_  (.A(net2109),
    .X(\imm13_b[7] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_766_  (.A(net1866),
    .X(\imm13_b[8] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_767_  (.A(net2067),
    .X(\imm13_b[9] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_768_  (.A(net2048),
    .X(\imm13_b[10] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_769_  (.A(net2178),
    .X(\imm13_b[12] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_770_  (.A(net1981),
    .X(\imm21_j[5] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_771_  (.A(net2069),
    .X(\imm21_j[6] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_772_  (.A(net2109),
    .X(\imm21_j[7] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_773_  (.A(net1866),
    .X(\imm21_j[8] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_774_  (.A(net2067),
    .X(\imm21_j[9] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_775_  (.A(net2048),
    .X(\imm21_j[10] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_776_  (.A(net2178),
    .X(\imm21_j[20] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_777_  (.A(\imm21_j[12] ),
    .X(\imm32_u[12] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_778_  (.A(\imm21_j[13] ),
    .X(\imm32_u[13] ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_779_  (.A(\imm21_j[14] ),
    .X(\imm32_u[14] ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_780_  (.A(\imm21_j[15] ),
    .X(\imm32_u[15] ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_781_  (.A(\imm21_j[16] ),
    .X(\imm32_u[16] ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_782_  (.A(\imm21_j[17] ),
    .X(\imm32_u[17] ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_783_  (.A(\imm21_j[18] ),
    .X(\imm32_u[18] ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_784_  (.A(\imm21_j[19] ),
    .X(\imm32_u[19] ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_785_  (.A(\imm21_j[11] ),
    .X(\imm32_u[20] ));
 sky130_fd_sc_hd__buf_1 \dec/_786_  (.A(\imm21_j[1] ),
    .X(\imm32_u[21] ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_787_  (.A(\imm21_j[2] ),
    .X(\imm32_u[22] ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_788_  (.A(\imm21_j[3] ),
    .X(\imm32_u[23] ));
 sky130_fd_sc_hd__clkbuf_2 \dec/_789_  (.A(\imm21_j[4] ),
    .X(\imm32_u[24] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_790_  (.A(\funct7[0] ),
    .X(\imm32_u[25] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_791_  (.A(\funct7[1] ),
    .X(\imm32_u[26] ));
 sky130_fd_sc_hd__buf_1 \dec/_792_  (.A(\funct7[2] ),
    .X(\imm32_u[27] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_793_  (.A(\funct7[3] ),
    .X(\imm32_u[28] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_794_  (.A(\funct7[4] ),
    .X(\imm32_u[29] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_795_  (.A(\funct7[5] ),
    .X(\imm32_u[30] ));
 sky130_fd_sc_hd__buf_1 \dec/_796_  (.A(\funct7[6] ),
    .X(\imm32_u[31] ));
 sky130_fd_sc_hd__buf_2 \dec/_797_  (.A(net897),
    .X(op_branch));
 sky130_fd_sc_hd__clkbuf_1 \dec/_798_  (.A(j_type),
    .X(op_jal));
 sky130_fd_sc_hd__buf_1 \dec/_799_  (.A(op_intRegReg),
    .X(r_type));
 sky130_fd_sc_hd__clkbuf_1 \dec/_800_  (.A(net1135),
    .X(\reg_d[0] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_801_  (.A(net1151),
    .X(\reg_d[1] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_802_  (.A(net1144),
    .X(\reg_d[2] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_803_  (.A(net1147),
    .X(\reg_d[3] ));
 sky130_fd_sc_hd__clkbuf_1 \dec/_804_  (.A(net1139),
    .X(\reg_d[4] ));
 sky130_fd_sc_hd__buf_2 \dec/_805_  (.A(op_memSt),
    .X(s_type));
 sky130_fd_sc_hd__inv_2 \reg_module/_09760_  (.A(net593),
    .Y(\reg_module/_02489_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_09761_  (.A(\reg_module/_02489_ ),
    .X(\reg_module/_02490_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_09762_  (.A(\reg_module/_02490_ ),
    .X(\reg_module/_02491_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_09763_  (.A(\reg_module/_02491_ ),
    .X(\reg_module/_02492_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_09764_  (.A(\reg_module/_02492_ ),
    .X(\reg_module/_02493_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09765_  (.A(\reg_module/_02493_ ),
    .B(\reg_module/gprf[800] ),
    .Y(\reg_module/_02494_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09766_  (.A(\reg_module/gprf[768] ),
    .B(net530),
    .Y(\reg_module/_02495_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09767_  (.A(\reg_module/_02494_ ),
    .B(net451),
    .C(\reg_module/_02495_ ),
    .Y(\reg_module/_02496_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_09768_  (.A(\reg_module/_02489_ ),
    .X(\reg_module/_02497_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_09769_  (.A(\reg_module/_02497_ ),
    .X(\reg_module/_02498_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09770_  (.A(\reg_module/_02498_ ),
    .X(\reg_module/_02499_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09771_  (.A(\reg_module/_02499_ ),
    .B(\reg_module/gprf[864] ),
    .Y(\reg_module/_02500_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_09772_  (.A(net452),
    .Y(\reg_module/_02501_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_09773_  (.A(\reg_module/_02501_ ),
    .X(\reg_module/_02502_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_09774_  (.A(\reg_module/_02502_ ),
    .X(\reg_module/_02503_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09775_  (.A(\reg_module/_02503_ ),
    .X(\reg_module/_02504_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09776_  (.A(\reg_module/gprf[832] ),
    .B(net530),
    .Y(\reg_module/_02505_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09777_  (.A(\reg_module/_02500_ ),
    .B(\reg_module/_02504_ ),
    .C(\reg_module/_02505_ ),
    .Y(\reg_module/_02506_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09778_  (.A(\reg_module/_02496_ ),
    .B(\reg_module/_02506_ ),
    .Y(\reg_module/_02507_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09779_  (.A(\reg_module/_02507_ ),
    .B(net410),
    .Y(\reg_module/_02508_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09780_  (.A(\reg_module/_02498_ ),
    .X(\reg_module/_02509_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09781_  (.A(\reg_module/_02509_ ),
    .B(\reg_module/gprf[928] ),
    .Y(\reg_module/_02510_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09782_  (.A(\reg_module/gprf[896] ),
    .B(net523),
    .Y(\reg_module/_02511_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09783_  (.A(\reg_module/_02510_ ),
    .B(net448),
    .C(\reg_module/_02511_ ),
    .Y(\reg_module/_02512_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_09784_  (.A(\reg_module/_02490_ ),
    .X(\reg_module/_02513_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09785_  (.A(\reg_module/_02513_ ),
    .X(\reg_module/_02514_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09786_  (.A(\reg_module/_02514_ ),
    .B(\reg_module/gprf[992] ),
    .Y(\reg_module/_02515_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_09787_  (.A(\reg_module/_02501_ ),
    .X(\reg_module/_02516_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09788_  (.A(\reg_module/_02516_ ),
    .X(\reg_module/_02517_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09789_  (.A(\reg_module/gprf[960] ),
    .B(net523),
    .Y(\reg_module/_02518_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09790_  (.A(\reg_module/_02515_ ),
    .B(\reg_module/_02517_ ),
    .C(\reg_module/_02518_ ),
    .Y(\reg_module/_02519_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09791_  (.A(\reg_module/_02512_ ),
    .B(\reg_module/_02519_ ),
    .Y(\reg_module/_02520_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_09792_  (.A(net430),
    .Y(\reg_module/_02521_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_09793_  (.A(\reg_module/_02521_ ),
    .X(\reg_module/_02522_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_09794_  (.A(\reg_module/_02522_ ),
    .X(\reg_module/_02523_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09795_  (.A(\reg_module/_02523_ ),
    .X(\reg_module/_02524_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09796_  (.A(\reg_module/_02520_ ),
    .B(\reg_module/_02524_ ),
    .Y(\reg_module/_02525_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_09797_  (.A(net389),
    .Y(\reg_module/_02526_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_09798_  (.A(\reg_module/_02526_ ),
    .X(\reg_module/_02527_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09799_  (.A(\reg_module/_02527_ ),
    .X(\reg_module/_02528_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09800_  (.A(\reg_module/_02508_ ),
    .B(\reg_module/_02525_ ),
    .C(\reg_module/_02528_ ),
    .Y(\reg_module/_02529_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_09801_  (.A(\reg_module/_02491_ ),
    .X(\reg_module/_02530_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_09802_  (.A(\reg_module/_02530_ ),
    .X(\reg_module/_02531_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09803_  (.A(\reg_module/_02531_ ),
    .B(\reg_module/gprf[672] ),
    .Y(\reg_module/_02532_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09804_  (.A(\reg_module/gprf[640] ),
    .B(net521),
    .Y(\reg_module/_02533_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09805_  (.A(\reg_module/_02532_ ),
    .B(net447),
    .C(\reg_module/_02533_ ),
    .Y(\reg_module/_02534_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_09806_  (.A(\reg_module/_02497_ ),
    .X(\reg_module/_02535_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_09807_  (.A(\reg_module/_02535_ ),
    .X(\reg_module/_02536_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09808_  (.A(\reg_module/_02536_ ),
    .B(\reg_module/gprf[736] ),
    .Y(\reg_module/_02537_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_09809_  (.A(\reg_module/_02501_ ),
    .X(\reg_module/_02538_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_09810_  (.A(\reg_module/_02538_ ),
    .X(\reg_module/_02539_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09811_  (.A(\reg_module/gprf[704] ),
    .B(net521),
    .Y(\reg_module/_02540_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09812_  (.A(\reg_module/_02537_ ),
    .B(\reg_module/_02539_ ),
    .C(\reg_module/_02540_ ),
    .Y(\reg_module/_02541_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09813_  (.A(\reg_module/_02534_ ),
    .B(\reg_module/_02541_ ),
    .Y(\reg_module/_02542_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09814_  (.A(\reg_module/_02523_ ),
    .X(\reg_module/_02543_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09815_  (.A(\reg_module/_02542_ ),
    .B(\reg_module/_02543_ ),
    .Y(\reg_module/_02544_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_09816_  (.A(\reg_module/_02497_ ),
    .X(\reg_module/_02545_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09817_  (.A(\reg_module/_02545_ ),
    .X(\reg_module/_02546_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09818_  (.A(\reg_module/_02546_ ),
    .B(\reg_module/gprf[544] ),
    .Y(\reg_module/_02547_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09819_  (.A(\reg_module/gprf[512] ),
    .B(net520),
    .Y(\reg_module/_02548_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09820_  (.A(\reg_module/_02547_ ),
    .B(net447),
    .C(\reg_module/_02548_ ),
    .Y(\reg_module/_02549_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_09821_  (.A(\reg_module/_02490_ ),
    .X(\reg_module/_02550_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_09822_  (.A(\reg_module/_02550_ ),
    .X(\reg_module/_02551_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09823_  (.A(\reg_module/_02551_ ),
    .B(\reg_module/gprf[608] ),
    .Y(\reg_module/_02552_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_09824_  (.A(\reg_module/_02501_ ),
    .X(\reg_module/_02553_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09825_  (.A(\reg_module/_02553_ ),
    .X(\reg_module/_02554_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09826_  (.A(\reg_module/gprf[576] ),
    .B(net520),
    .Y(\reg_module/_02555_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09827_  (.A(\reg_module/_02552_ ),
    .B(\reg_module/_02554_ ),
    .C(\reg_module/_02555_ ),
    .Y(\reg_module/_02556_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09828_  (.A(\reg_module/_02549_ ),
    .B(\reg_module/_02556_ ),
    .Y(\reg_module/_02557_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09829_  (.A(\reg_module/_02557_ ),
    .B(net408),
    .Y(\reg_module/_02558_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09830_  (.A(\reg_module/_02544_ ),
    .B(\reg_module/_02558_ ),
    .C(net388),
    .Y(\reg_module/_02559_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09831_  (.A(\reg_module/_02529_ ),
    .B(\reg_module/_02559_ ),
    .Y(\reg_module/_02560_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_09832_  (.A(net383),
    .Y(\reg_module/_02561_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_09833_  (.A(\reg_module/_02561_ ),
    .X(\reg_module/_02562_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_09834_  (.A(\reg_module/_02562_ ),
    .X(\reg_module/_02563_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09835_  (.A(\reg_module/_02560_ ),
    .B(\reg_module/_02563_ ),
    .Y(\reg_module/_02564_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_09836_  (.A(\reg_module/_02491_ ),
    .X(\reg_module/_02565_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09837_  (.A(\reg_module/_02565_ ),
    .X(\reg_module/_02566_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09838_  (.A(\reg_module/_02566_ ),
    .B(\reg_module/gprf[288] ),
    .Y(\reg_module/_02567_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09839_  (.A(\reg_module/gprf[256] ),
    .B(net529),
    .Y(\reg_module/_02568_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09840_  (.A(\reg_module/_02567_ ),
    .B(net451),
    .C(\reg_module/_02568_ ),
    .Y(\reg_module/_02569_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_09841_  (.A(\reg_module/_02497_ ),
    .X(\reg_module/_02570_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_09842_  (.A(\reg_module/_02570_ ),
    .X(\reg_module/_02571_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09843_  (.A(\reg_module/_02571_ ),
    .B(\reg_module/gprf[352] ),
    .Y(\reg_module/_02572_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_09844_  (.A(\reg_module/_02502_ ),
    .X(\reg_module/_02573_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09845_  (.A(\reg_module/_02573_ ),
    .X(\reg_module/_02574_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09846_  (.A(\reg_module/gprf[320] ),
    .B(net529),
    .Y(\reg_module/_02575_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09847_  (.A(\reg_module/_02572_ ),
    .B(\reg_module/_02574_ ),
    .C(\reg_module/_02575_ ),
    .Y(\reg_module/_02576_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09848_  (.A(\reg_module/_02569_ ),
    .B(\reg_module/_02576_ ),
    .Y(\reg_module/_02577_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09849_  (.A(\reg_module/_02577_ ),
    .B(net407),
    .Y(\reg_module/_02578_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_09850_  (.A(\reg_module/_02497_ ),
    .X(\reg_module/_02579_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09851_  (.A(\reg_module/_02579_ ),
    .X(\reg_module/_02580_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09852_  (.A(\reg_module/_02580_ ),
    .B(\reg_module/gprf[416] ),
    .Y(\reg_module/_02581_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09853_  (.A(\reg_module/gprf[384] ),
    .B(net522),
    .Y(\reg_module/_02582_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09854_  (.A(\reg_module/_02581_ ),
    .B(net448),
    .C(\reg_module/_02582_ ),
    .Y(\reg_module/_02583_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_09855_  (.A(\reg_module/_02490_ ),
    .X(\reg_module/_02584_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09856_  (.A(\reg_module/_02584_ ),
    .X(\reg_module/_02585_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09857_  (.A(\reg_module/_02585_ ),
    .B(\reg_module/gprf[480] ),
    .Y(\reg_module/_02586_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_09858_  (.A(\reg_module/_02501_ ),
    .X(\reg_module/_02587_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_09859_  (.A(\reg_module/_02587_ ),
    .X(\reg_module/_02588_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09860_  (.A(\reg_module/gprf[448] ),
    .B(net522),
    .Y(\reg_module/_02589_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09861_  (.A(\reg_module/_02586_ ),
    .B(\reg_module/_02588_ ),
    .C(\reg_module/_02589_ ),
    .Y(\reg_module/_02590_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09862_  (.A(\reg_module/_02583_ ),
    .B(\reg_module/_02590_ ),
    .Y(\reg_module/_02591_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_09863_  (.A(\reg_module/_02521_ ),
    .X(\reg_module/_02592_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_09864_  (.A(\reg_module/_02592_ ),
    .X(\reg_module/_02593_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09865_  (.A(\reg_module/_02591_ ),
    .B(\reg_module/_02593_ ),
    .Y(\reg_module/_02594_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_09866_  (.A(\reg_module/_02526_ ),
    .X(\reg_module/_02595_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09867_  (.A(\reg_module/_02595_ ),
    .X(\reg_module/_02596_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09868_  (.A(\reg_module/_02578_ ),
    .B(\reg_module/_02594_ ),
    .C(\reg_module/_02596_ ),
    .Y(\reg_module/_02597_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09869_  (.A(\reg_module/_02571_ ),
    .B(\reg_module/gprf[32] ),
    .Y(\reg_module/_02598_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09870_  (.A(\reg_module/gprf[0] ),
    .B(net521),
    .Y(\reg_module/_02599_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09871_  (.A(\reg_module/_02598_ ),
    .B(net447),
    .C(\reg_module/_02599_ ),
    .Y(\reg_module/_02600_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_09872_  (.A(\reg_module/_02490_ ),
    .X(\reg_module/_02601_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09873_  (.A(\reg_module/_02601_ ),
    .X(\reg_module/_02602_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09874_  (.A(\reg_module/_02602_ ),
    .B(\reg_module/gprf[96] ),
    .Y(\reg_module/_02603_ ));
 sky130_fd_sc_hd__buf_8 \reg_module/_09875_  (.A(\reg_module/_02501_ ),
    .X(\reg_module/_02604_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09876_  (.A(\reg_module/_02604_ ),
    .X(\reg_module/_02605_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09877_  (.A(\reg_module/gprf[64] ),
    .B(net521),
    .Y(\reg_module/_02606_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09878_  (.A(\reg_module/_02603_ ),
    .B(\reg_module/_02605_ ),
    .C(\reg_module/_02606_ ),
    .Y(\reg_module/_02607_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09879_  (.A(\reg_module/_02600_ ),
    .B(\reg_module/_02607_ ),
    .Y(\reg_module/_02608_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09880_  (.A(\reg_module/_02608_ ),
    .B(net407),
    .Y(\reg_module/_02609_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09881_  (.A(\reg_module/_02584_ ),
    .X(\reg_module/_02610_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09882_  (.A(\reg_module/_02610_ ),
    .B(\reg_module/gprf[160] ),
    .Y(\reg_module/_02611_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09883_  (.A(\reg_module/gprf[128] ),
    .B(net519),
    .Y(\reg_module/_02612_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09884_  (.A(\reg_module/_02611_ ),
    .B(net447),
    .C(\reg_module/_02612_ ),
    .Y(\reg_module/_02613_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_09885_  (.A(\reg_module/_02490_ ),
    .X(\reg_module/_02614_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09886_  (.A(\reg_module/_02614_ ),
    .X(\reg_module/_02615_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09887_  (.A(\reg_module/_02615_ ),
    .B(\reg_module/gprf[224] ),
    .Y(\reg_module/_02616_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09888_  (.A(\reg_module/_02553_ ),
    .X(\reg_module/_02617_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09889_  (.A(\reg_module/gprf[192] ),
    .B(net519),
    .Y(\reg_module/_02618_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09890_  (.A(\reg_module/_02616_ ),
    .B(\reg_module/_02617_ ),
    .C(\reg_module/_02618_ ),
    .Y(\reg_module/_02619_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09891_  (.A(\reg_module/_02613_ ),
    .B(\reg_module/_02619_ ),
    .Y(\reg_module/_02620_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09892_  (.A(\reg_module/_02522_ ),
    .X(\reg_module/_02621_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09893_  (.A(\reg_module/_02620_ ),
    .B(\reg_module/_02621_ ),
    .Y(\reg_module/_02622_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09894_  (.A(\reg_module/_02609_ ),
    .B(\reg_module/_02622_ ),
    .C(net388),
    .Y(\reg_module/_02623_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09895_  (.A(\reg_module/_02597_ ),
    .B(\reg_module/_02623_ ),
    .Y(\reg_module/_02624_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09896_  (.A(\reg_module/_02624_ ),
    .B(net380),
    .Y(\reg_module/_02625_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_09897_  (.A(\reg_module/_02564_ ),
    .B(\reg_module/_02625_ ),
    .Y(\wRs2Data[0] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09898_  (.A(\reg_module/_02493_ ),
    .B(\reg_module/gprf[801] ),
    .Y(\reg_module/_02626_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09899_  (.A(\reg_module/gprf[769] ),
    .B(net570),
    .Y(\reg_module/_02627_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09900_  (.A(\reg_module/_02626_ ),
    .B(net474),
    .C(\reg_module/_02627_ ),
    .Y(\reg_module/_02628_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09901_  (.A(\reg_module/_02499_ ),
    .B(\reg_module/gprf[865] ),
    .Y(\reg_module/_02629_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09902_  (.A(\reg_module/gprf[833] ),
    .B(net529),
    .Y(\reg_module/_02630_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09903_  (.A(\reg_module/_02629_ ),
    .B(\reg_module/_02504_ ),
    .C(\reg_module/_02630_ ),
    .Y(\reg_module/_02631_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09904_  (.A(\reg_module/_02628_ ),
    .B(\reg_module/_02631_ ),
    .Y(\reg_module/_02632_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09905_  (.A(\reg_module/_02632_ ),
    .B(net408),
    .Y(\reg_module/_02633_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09906_  (.A(\reg_module/_02509_ ),
    .B(\reg_module/gprf[929] ),
    .Y(\reg_module/_02634_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09907_  (.A(\reg_module/gprf[897] ),
    .B(net522),
    .Y(\reg_module/_02635_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09908_  (.A(\reg_module/_02634_ ),
    .B(net448),
    .C(\reg_module/_02635_ ),
    .Y(\reg_module/_02636_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09909_  (.A(\reg_module/_02514_ ),
    .B(\reg_module/gprf[993] ),
    .Y(\reg_module/_02637_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09910_  (.A(\reg_module/gprf[961] ),
    .B(net522),
    .Y(\reg_module/_02638_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09911_  (.A(\reg_module/_02637_ ),
    .B(\reg_module/_02517_ ),
    .C(\reg_module/_02638_ ),
    .Y(\reg_module/_02639_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09912_  (.A(\reg_module/_02636_ ),
    .B(\reg_module/_02639_ ),
    .Y(\reg_module/_02640_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09913_  (.A(\reg_module/_02640_ ),
    .B(\reg_module/_02524_ ),
    .Y(\reg_module/_02641_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09914_  (.A(\reg_module/_02633_ ),
    .B(\reg_module/_02641_ ),
    .C(\reg_module/_02528_ ),
    .Y(\reg_module/_02642_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09915_  (.A(\reg_module/_02531_ ),
    .B(\reg_module/gprf[673] ),
    .Y(\reg_module/_02643_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09916_  (.A(\reg_module/gprf[641] ),
    .B(net519),
    .Y(\reg_module/_02644_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09917_  (.A(\reg_module/_02643_ ),
    .B(net447),
    .C(\reg_module/_02644_ ),
    .Y(\reg_module/_02645_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09918_  (.A(\reg_module/_02536_ ),
    .B(\reg_module/gprf[737] ),
    .Y(\reg_module/_02646_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09919_  (.A(\reg_module/gprf[705] ),
    .B(net520),
    .Y(\reg_module/_02647_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09920_  (.A(\reg_module/_02646_ ),
    .B(\reg_module/_02539_ ),
    .C(\reg_module/_02647_ ),
    .Y(\reg_module/_02648_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09921_  (.A(\reg_module/_02645_ ),
    .B(\reg_module/_02648_ ),
    .Y(\reg_module/_02649_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09922_  (.A(\reg_module/_02649_ ),
    .B(\reg_module/_02543_ ),
    .Y(\reg_module/_02650_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09923_  (.A(\reg_module/_02546_ ),
    .B(\reg_module/gprf[545] ),
    .Y(\reg_module/_02651_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09924_  (.A(\reg_module/gprf[513] ),
    .B(net561),
    .Y(\reg_module/_02652_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09925_  (.A(\reg_module/_02651_ ),
    .B(net469),
    .C(\reg_module/_02652_ ),
    .Y(\reg_module/_02653_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09926_  (.A(\reg_module/_02551_ ),
    .B(\reg_module/gprf[609] ),
    .Y(\reg_module/_02654_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09927_  (.A(\reg_module/gprf[577] ),
    .B(net519),
    .Y(\reg_module/_02655_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09928_  (.A(\reg_module/_02654_ ),
    .B(\reg_module/_02554_ ),
    .C(\reg_module/_02655_ ),
    .Y(\reg_module/_02656_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09929_  (.A(\reg_module/_02653_ ),
    .B(\reg_module/_02656_ ),
    .Y(\reg_module/_02657_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09930_  (.A(\reg_module/_02657_ ),
    .B(net408),
    .Y(\reg_module/_02658_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09931_  (.A(\reg_module/_02650_ ),
    .B(\reg_module/_02658_ ),
    .C(net388),
    .Y(\reg_module/_02659_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09932_  (.A(\reg_module/_02642_ ),
    .B(\reg_module/_02659_ ),
    .Y(\reg_module/_02660_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09933_  (.A(\reg_module/_02660_ ),
    .B(\reg_module/_02563_ ),
    .Y(\reg_module/_02661_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09934_  (.A(\reg_module/_02566_ ),
    .B(\reg_module/gprf[289] ),
    .Y(\reg_module/_02662_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09935_  (.A(\reg_module/gprf[257] ),
    .B(net530),
    .Y(\reg_module/_02663_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09936_  (.A(\reg_module/_02662_ ),
    .B(net451),
    .C(\reg_module/_02663_ ),
    .Y(\reg_module/_02664_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09937_  (.A(\reg_module/_02570_ ),
    .X(\reg_module/_02665_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09938_  (.A(\reg_module/_02665_ ),
    .B(\reg_module/gprf[353] ),
    .Y(\reg_module/_02666_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09939_  (.A(\reg_module/gprf[321] ),
    .B(net530),
    .Y(\reg_module/_02667_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09940_  (.A(\reg_module/_02666_ ),
    .B(\reg_module/_02574_ ),
    .C(\reg_module/_02667_ ),
    .Y(\reg_module/_02668_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09941_  (.A(\reg_module/_02664_ ),
    .B(\reg_module/_02668_ ),
    .Y(\reg_module/_02669_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09942_  (.A(\reg_module/_02669_ ),
    .B(net408),
    .Y(\reg_module/_02670_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09943_  (.A(\reg_module/_02580_ ),
    .B(\reg_module/gprf[417] ),
    .Y(\reg_module/_02671_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09944_  (.A(\reg_module/gprf[385] ),
    .B(net522),
    .Y(\reg_module/_02672_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09945_  (.A(\reg_module/_02671_ ),
    .B(net448),
    .C(\reg_module/_02672_ ),
    .Y(\reg_module/_02673_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09946_  (.A(\reg_module/_02585_ ),
    .B(\reg_module/gprf[481] ),
    .Y(\reg_module/_02674_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09947_  (.A(\reg_module/gprf[449] ),
    .B(net522),
    .Y(\reg_module/_02675_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09948_  (.A(\reg_module/_02674_ ),
    .B(\reg_module/_02588_ ),
    .C(\reg_module/_02675_ ),
    .Y(\reg_module/_02676_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09949_  (.A(\reg_module/_02673_ ),
    .B(\reg_module/_02676_ ),
    .Y(\reg_module/_02677_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09950_  (.A(\reg_module/_02677_ ),
    .B(\reg_module/_02593_ ),
    .Y(\reg_module/_02678_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09951_  (.A(\reg_module/_02670_ ),
    .B(\reg_module/_02678_ ),
    .C(\reg_module/_02596_ ),
    .Y(\reg_module/_02679_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09952_  (.A(\reg_module/_02665_ ),
    .B(\reg_module/gprf[33] ),
    .Y(\reg_module/_02680_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09953_  (.A(\reg_module/gprf[1] ),
    .B(net561),
    .Y(\reg_module/_02681_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09954_  (.A(\reg_module/_02680_ ),
    .B(net469),
    .C(\reg_module/_02681_ ),
    .Y(\reg_module/_02682_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09955_  (.A(\reg_module/_02602_ ),
    .B(\reg_module/gprf[97] ),
    .Y(\reg_module/_02683_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09956_  (.A(\reg_module/gprf[65] ),
    .B(net521),
    .Y(\reg_module/_02684_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09957_  (.A(\reg_module/_02683_ ),
    .B(\reg_module/_02605_ ),
    .C(\reg_module/_02684_ ),
    .Y(\reg_module/_02685_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09958_  (.A(\reg_module/_02682_ ),
    .B(\reg_module/_02685_ ),
    .Y(\reg_module/_02686_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09959_  (.A(\reg_module/_02686_ ),
    .B(net408),
    .Y(\reg_module/_02687_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09960_  (.A(\reg_module/_02610_ ),
    .B(\reg_module/gprf[161] ),
    .Y(\reg_module/_02688_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09961_  (.A(\reg_module/gprf[129] ),
    .B(net519),
    .Y(\reg_module/_02689_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09962_  (.A(\reg_module/_02688_ ),
    .B(net447),
    .C(\reg_module/_02689_ ),
    .Y(\reg_module/_02690_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09963_  (.A(\reg_module/_02615_ ),
    .B(\reg_module/gprf[225] ),
    .Y(\reg_module/_02691_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09964_  (.A(\reg_module/gprf[193] ),
    .B(net519),
    .Y(\reg_module/_02692_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09965_  (.A(\reg_module/_02691_ ),
    .B(\reg_module/_02617_ ),
    .C(\reg_module/_02692_ ),
    .Y(\reg_module/_02693_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09966_  (.A(\reg_module/_02690_ ),
    .B(\reg_module/_02693_ ),
    .Y(\reg_module/_02694_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09967_  (.A(\reg_module/_02694_ ),
    .B(\reg_module/_02621_ ),
    .Y(\reg_module/_02695_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09968_  (.A(\reg_module/_02687_ ),
    .B(\reg_module/_02695_ ),
    .C(net388),
    .Y(\reg_module/_02696_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09969_  (.A(\reg_module/_02679_ ),
    .B(\reg_module/_02696_ ),
    .Y(\reg_module/_02697_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09970_  (.A(\reg_module/_02697_ ),
    .B(net380),
    .Y(\reg_module/_02698_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_09971_  (.A(\reg_module/_02661_ ),
    .B(\reg_module/_02698_ ),
    .Y(\wRs2Data[1] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09972_  (.A(\reg_module/_02493_ ),
    .B(\reg_module/gprf[546] ),
    .Y(\reg_module/_02699_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09973_  (.A(\reg_module/gprf[514] ),
    .B(net565),
    .Y(\reg_module/_02700_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09974_  (.A(\reg_module/_02699_ ),
    .B(net471),
    .C(\reg_module/_02700_ ),
    .Y(\reg_module/_02701_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09975_  (.A(\reg_module/_02499_ ),
    .B(\reg_module/gprf[610] ),
    .Y(\reg_module/_02702_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09976_  (.A(\reg_module/gprf[578] ),
    .B(net567),
    .Y(\reg_module/_02703_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09977_  (.A(\reg_module/_02702_ ),
    .B(\reg_module/_02504_ ),
    .C(\reg_module/_02703_ ),
    .Y(\reg_module/_02704_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09978_  (.A(\reg_module/_02701_ ),
    .B(\reg_module/_02704_ ),
    .Y(\reg_module/_02705_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09979_  (.A(\reg_module/_02705_ ),
    .B(net421),
    .Y(\reg_module/_02706_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09980_  (.A(\reg_module/_02509_ ),
    .B(\reg_module/gprf[674] ),
    .Y(\reg_module/_02707_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09981_  (.A(\reg_module/gprf[642] ),
    .B(net565),
    .Y(\reg_module/_02708_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09982_  (.A(\reg_module/_02707_ ),
    .B(net471),
    .C(\reg_module/_02708_ ),
    .Y(\reg_module/_02709_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09983_  (.A(\reg_module/_02514_ ),
    .B(\reg_module/gprf[738] ),
    .Y(\reg_module/_02710_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09984_  (.A(\reg_module/gprf[706] ),
    .B(net565),
    .Y(\reg_module/_02711_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09985_  (.A(\reg_module/_02710_ ),
    .B(\reg_module/_02517_ ),
    .C(\reg_module/_02711_ ),
    .Y(\reg_module/_02712_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09986_  (.A(\reg_module/_02709_ ),
    .B(\reg_module/_02712_ ),
    .Y(\reg_module/_02713_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_09987_  (.A(\reg_module/_02592_ ),
    .X(\reg_module/_02714_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09988_  (.A(\reg_module/_02713_ ),
    .B(\reg_module/_02714_ ),
    .Y(\reg_module/_02715_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09989_  (.A(\reg_module/_02706_ ),
    .B(\reg_module/_02715_ ),
    .C(net396),
    .Y(\reg_module/_02716_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09990_  (.A(\reg_module/_02530_ ),
    .X(\reg_module/_02717_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09991_  (.A(\reg_module/_02717_ ),
    .B(\reg_module/gprf[802] ),
    .Y(\reg_module/_02718_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09992_  (.A(\reg_module/gprf[770] ),
    .B(net570),
    .Y(\reg_module/_02719_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09993_  (.A(\reg_module/_02718_ ),
    .B(net474),
    .C(\reg_module/_02719_ ),
    .Y(\reg_module/_02720_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09994_  (.A(\reg_module/_02536_ ),
    .B(\reg_module/gprf[866] ),
    .Y(\reg_module/_02721_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_09995_  (.A(\reg_module/_02538_ ),
    .X(\reg_module/_02722_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09996_  (.A(\reg_module/gprf[834] ),
    .B(net572),
    .Y(\reg_module/_02723_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_09997_  (.A(\reg_module/_02721_ ),
    .B(\reg_module/_02722_ ),
    .C(\reg_module/_02723_ ),
    .Y(\reg_module/_02724_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09998_  (.A(\reg_module/_02720_ ),
    .B(\reg_module/_02724_ ),
    .Y(\reg_module/_02725_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_09999_  (.A(\reg_module/_02725_ ),
    .B(net423),
    .Y(\reg_module/_02726_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10000_  (.A(\reg_module/_02546_ ),
    .B(\reg_module/gprf[930] ),
    .Y(\reg_module/_02727_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10001_  (.A(\reg_module/gprf[898] ),
    .B(net562),
    .Y(\reg_module/_02728_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10002_  (.A(\reg_module/_02727_ ),
    .B(net470),
    .C(\reg_module/_02728_ ),
    .Y(\reg_module/_02729_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_10003_  (.A(\reg_module/_02550_ ),
    .X(\reg_module/_02730_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10004_  (.A(\reg_module/_02730_ ),
    .B(\reg_module/gprf[994] ),
    .Y(\reg_module/_02731_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10005_  (.A(\reg_module/gprf[962] ),
    .B(net562),
    .Y(\reg_module/_02732_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10006_  (.A(\reg_module/_02731_ ),
    .B(\reg_module/_02554_ ),
    .C(\reg_module/_02732_ ),
    .Y(\reg_module/_02733_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10007_  (.A(\reg_module/_02729_ ),
    .B(\reg_module/_02733_ ),
    .Y(\reg_module/_02734_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_10008_  (.A(\reg_module/_02521_ ),
    .X(\reg_module/_02735_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_10009_  (.A(\reg_module/_02735_ ),
    .X(\reg_module/_02736_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10010_  (.A(\reg_module/_02734_ ),
    .B(\reg_module/_02736_ ),
    .Y(\reg_module/_02737_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_10011_  (.A(\reg_module/_02526_ ),
    .X(\reg_module/_02738_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10012_  (.A(\reg_module/_02726_ ),
    .B(\reg_module/_02737_ ),
    .C(\reg_module/_02738_ ),
    .Y(\reg_module/_02739_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10013_  (.A(\reg_module/_02716_ ),
    .B(\reg_module/_02739_ ),
    .Y(\reg_module/_02740_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10014_  (.A(\reg_module/_02740_ ),
    .B(\reg_module/_02563_ ),
    .Y(\reg_module/_02741_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10015_  (.A(\reg_module/_02566_ ),
    .B(\reg_module/gprf[290] ),
    .Y(\reg_module/_02742_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10016_  (.A(\reg_module/gprf[258] ),
    .B(net570),
    .Y(\reg_module/_02743_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10017_  (.A(\reg_module/_02742_ ),
    .B(net474),
    .C(\reg_module/_02743_ ),
    .Y(\reg_module/_02744_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10018_  (.A(\reg_module/_02665_ ),
    .B(\reg_module/gprf[354] ),
    .Y(\reg_module/_02745_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10019_  (.A(\reg_module/gprf[322] ),
    .B(net571),
    .Y(\reg_module/_02746_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10020_  (.A(\reg_module/_02745_ ),
    .B(\reg_module/_02574_ ),
    .C(\reg_module/_02746_ ),
    .Y(\reg_module/_02747_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10021_  (.A(\reg_module/_02744_ ),
    .B(\reg_module/_02747_ ),
    .Y(\reg_module/_02748_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10022_  (.A(\reg_module/_02748_ ),
    .B(net423),
    .Y(\reg_module/_02749_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10023_  (.A(\reg_module/_02579_ ),
    .X(\reg_module/_02750_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10024_  (.A(\reg_module/_02750_ ),
    .B(\reg_module/gprf[418] ),
    .Y(\reg_module/_02751_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10025_  (.A(\reg_module/gprf[386] ),
    .B(net562),
    .Y(\reg_module/_02752_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10026_  (.A(\reg_module/_02751_ ),
    .B(net469),
    .C(\reg_module/_02752_ ),
    .Y(\reg_module/_02753_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10027_  (.A(\reg_module/_02585_ ),
    .B(\reg_module/gprf[482] ),
    .Y(\reg_module/_02754_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10028_  (.A(\reg_module/_02587_ ),
    .X(\reg_module/_02755_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10029_  (.A(\reg_module/gprf[450] ),
    .B(net562),
    .Y(\reg_module/_02756_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10030_  (.A(\reg_module/_02754_ ),
    .B(\reg_module/_02755_ ),
    .C(\reg_module/_02756_ ),
    .Y(\reg_module/_02757_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10031_  (.A(\reg_module/_02753_ ),
    .B(\reg_module/_02757_ ),
    .Y(\reg_module/_02758_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10032_  (.A(\reg_module/_02758_ ),
    .B(\reg_module/_02593_ ),
    .Y(\reg_module/_02759_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10033_  (.A(\reg_module/_02595_ ),
    .X(\reg_module/_02760_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10034_  (.A(\reg_module/_02749_ ),
    .B(\reg_module/_02759_ ),
    .C(\reg_module/_02760_ ),
    .Y(\reg_module/_02761_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10035_  (.A(\reg_module/_02665_ ),
    .B(\reg_module/gprf[34] ),
    .Y(\reg_module/_02762_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10036_  (.A(\reg_module/gprf[2] ),
    .B(net561),
    .Y(\reg_module/_02763_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10037_  (.A(\reg_module/_02762_ ),
    .B(net469),
    .C(\reg_module/_02763_ ),
    .Y(\reg_module/_02764_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_10038_  (.A(\reg_module/_02601_ ),
    .X(\reg_module/_02765_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10039_  (.A(\reg_module/_02765_ ),
    .B(\reg_module/gprf[98] ),
    .Y(\reg_module/_02766_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10040_  (.A(\reg_module/gprf[66] ),
    .B(net561),
    .Y(\reg_module/_02767_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10041_  (.A(\reg_module/_02766_ ),
    .B(\reg_module/_02605_ ),
    .C(\reg_module/_02767_ ),
    .Y(\reg_module/_02768_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10042_  (.A(\reg_module/_02764_ ),
    .B(\reg_module/_02768_ ),
    .Y(\reg_module/_02769_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10043_  (.A(\reg_module/_02769_ ),
    .B(net421),
    .Y(\reg_module/_02770_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10044_  (.A(\reg_module/_02610_ ),
    .B(\reg_module/gprf[162] ),
    .Y(\reg_module/_02771_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10045_  (.A(\reg_module/gprf[130] ),
    .B(net564),
    .Y(\reg_module/_02772_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10046_  (.A(\reg_module/_02771_ ),
    .B(net469),
    .C(\reg_module/_02772_ ),
    .Y(\reg_module/_02773_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10047_  (.A(\reg_module/_02615_ ),
    .B(\reg_module/gprf[226] ),
    .Y(\reg_module/_02774_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10048_  (.A(\reg_module/gprf[194] ),
    .B(net561),
    .Y(\reg_module/_02775_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10049_  (.A(\reg_module/_02774_ ),
    .B(\reg_module/_02617_ ),
    .C(\reg_module/_02775_ ),
    .Y(\reg_module/_02776_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10050_  (.A(\reg_module/_02773_ ),
    .B(\reg_module/_02776_ ),
    .Y(\reg_module/_02777_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10051_  (.A(\reg_module/_02777_ ),
    .B(\reg_module/_02621_ ),
    .Y(\reg_module/_02778_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10052_  (.A(\reg_module/_02770_ ),
    .B(\reg_module/_02778_ ),
    .C(net396),
    .Y(\reg_module/_02779_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10053_  (.A(\reg_module/_02761_ ),
    .B(\reg_module/_02779_ ),
    .Y(\reg_module/_02780_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10054_  (.A(\reg_module/_02780_ ),
    .B(net381),
    .Y(\reg_module/_02781_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_10055_  (.A(\reg_module/_02741_ ),
    .B(\reg_module/_02781_ ),
    .Y(\wRs2Data[2] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10056_  (.A(\reg_module/_02493_ ),
    .B(\reg_module/gprf[803] ),
    .Y(\reg_module/_02782_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10057_  (.A(\reg_module/gprf[771] ),
    .B(net572),
    .Y(\reg_module/_02783_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10058_  (.A(\reg_module/_02782_ ),
    .B(net475),
    .C(\reg_module/_02783_ ),
    .Y(\reg_module/_02784_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10059_  (.A(\reg_module/_02499_ ),
    .B(\reg_module/gprf[867] ),
    .Y(\reg_module/_02785_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10060_  (.A(\reg_module/gprf[835] ),
    .B(net567),
    .Y(\reg_module/_02786_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10061_  (.A(\reg_module/_02785_ ),
    .B(\reg_module/_02504_ ),
    .C(\reg_module/_02786_ ),
    .Y(\reg_module/_02787_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10062_  (.A(\reg_module/_02784_ ),
    .B(\reg_module/_02787_ ),
    .Y(\reg_module/_02788_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10063_  (.A(\reg_module/_02788_ ),
    .B(net422),
    .Y(\reg_module/_02789_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10064_  (.A(\reg_module/_02509_ ),
    .B(\reg_module/gprf[931] ),
    .Y(\reg_module/_02790_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10065_  (.A(\reg_module/gprf[899] ),
    .B(net567),
    .Y(\reg_module/_02791_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10066_  (.A(\reg_module/_02790_ ),
    .B(net472),
    .C(\reg_module/_02791_ ),
    .Y(\reg_module/_02792_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10067_  (.A(\reg_module/_02514_ ),
    .B(\reg_module/gprf[995] ),
    .Y(\reg_module/_02793_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10068_  (.A(\reg_module/gprf[963] ),
    .B(net567),
    .Y(\reg_module/_02794_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10069_  (.A(\reg_module/_02793_ ),
    .B(\reg_module/_02517_ ),
    .C(\reg_module/_02794_ ),
    .Y(\reg_module/_02795_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10070_  (.A(\reg_module/_02792_ ),
    .B(\reg_module/_02795_ ),
    .Y(\reg_module/_02796_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10071_  (.A(\reg_module/_02796_ ),
    .B(\reg_module/_02714_ ),
    .Y(\reg_module/_02797_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10072_  (.A(\reg_module/_02789_ ),
    .B(\reg_module/_02797_ ),
    .C(\reg_module/_02528_ ),
    .Y(\reg_module/_02798_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10073_  (.A(\reg_module/_02717_ ),
    .B(\reg_module/gprf[675] ),
    .Y(\reg_module/_02799_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10074_  (.A(\reg_module/gprf[643] ),
    .B(net566),
    .Y(\reg_module/_02800_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10075_  (.A(\reg_module/_02799_ ),
    .B(net471),
    .C(\reg_module/_02800_ ),
    .Y(\reg_module/_02801_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10076_  (.A(\reg_module/_02536_ ),
    .B(\reg_module/gprf[739] ),
    .Y(\reg_module/_02802_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10077_  (.A(\reg_module/gprf[707] ),
    .B(net566),
    .Y(\reg_module/_02803_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10078_  (.A(\reg_module/_02802_ ),
    .B(\reg_module/_02722_ ),
    .C(\reg_module/_02803_ ),
    .Y(\reg_module/_02804_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10079_  (.A(\reg_module/_02801_ ),
    .B(\reg_module/_02804_ ),
    .Y(\reg_module/_02805_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10080_  (.A(\reg_module/_02805_ ),
    .B(\reg_module/_02543_ ),
    .Y(\reg_module/_02806_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10081_  (.A(\reg_module/_02546_ ),
    .B(\reg_module/gprf[547] ),
    .Y(\reg_module/_02807_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10082_  (.A(\reg_module/gprf[515] ),
    .B(net579),
    .Y(\reg_module/_02808_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10083_  (.A(\reg_module/_02807_ ),
    .B(net478),
    .C(\reg_module/_02808_ ),
    .Y(\reg_module/_02809_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10084_  (.A(\reg_module/_02730_ ),
    .B(\reg_module/gprf[611] ),
    .Y(\reg_module/_02810_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10085_  (.A(\reg_module/gprf[579] ),
    .B(net580),
    .Y(\reg_module/_02811_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10086_  (.A(\reg_module/_02810_ ),
    .B(\reg_module/_02554_ ),
    .C(\reg_module/_02811_ ),
    .Y(\reg_module/_02812_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10087_  (.A(\reg_module/_02809_ ),
    .B(\reg_module/_02812_ ),
    .Y(\reg_module/_02813_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10088_  (.A(\reg_module/_02813_ ),
    .B(net421),
    .Y(\reg_module/_02814_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10089_  (.A(\reg_module/_02806_ ),
    .B(\reg_module/_02814_ ),
    .C(net396),
    .Y(\reg_module/_02815_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10090_  (.A(\reg_module/_02798_ ),
    .B(\reg_module/_02815_ ),
    .Y(\reg_module/_02816_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10091_  (.A(\reg_module/_02816_ ),
    .B(\reg_module/_02563_ ),
    .Y(\reg_module/_02817_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10092_  (.A(\reg_module/_02566_ ),
    .B(\reg_module/gprf[291] ),
    .Y(\reg_module/_02818_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10093_  (.A(\reg_module/gprf[259] ),
    .B(net570),
    .Y(\reg_module/_02819_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10094_  (.A(\reg_module/_02818_ ),
    .B(net474),
    .C(\reg_module/_02819_ ),
    .Y(\reg_module/_02820_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10095_  (.A(\reg_module/_02665_ ),
    .B(\reg_module/gprf[355] ),
    .Y(\reg_module/_02821_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10096_  (.A(\reg_module/gprf[323] ),
    .B(net572),
    .Y(\reg_module/_02822_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10097_  (.A(\reg_module/_02821_ ),
    .B(\reg_module/_02574_ ),
    .C(\reg_module/_02822_ ),
    .Y(\reg_module/_02823_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10098_  (.A(\reg_module/_02820_ ),
    .B(\reg_module/_02823_ ),
    .Y(\reg_module/_02824_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10099_  (.A(\reg_module/_02824_ ),
    .B(net421),
    .Y(\reg_module/_02825_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10100_  (.A(\reg_module/_02750_ ),
    .B(\reg_module/gprf[419] ),
    .Y(\reg_module/_02826_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10101_  (.A(\reg_module/gprf[387] ),
    .B(net562),
    .Y(\reg_module/_02827_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10102_  (.A(\reg_module/_02826_ ),
    .B(net470),
    .C(\reg_module/_02827_ ),
    .Y(\reg_module/_02828_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10103_  (.A(\reg_module/_02585_ ),
    .B(\reg_module/gprf[483] ),
    .Y(\reg_module/_02829_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10104_  (.A(\reg_module/gprf[451] ),
    .B(net562),
    .Y(\reg_module/_02830_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10105_  (.A(\reg_module/_02829_ ),
    .B(\reg_module/_02755_ ),
    .C(\reg_module/_02830_ ),
    .Y(\reg_module/_02831_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10106_  (.A(\reg_module/_02828_ ),
    .B(\reg_module/_02831_ ),
    .Y(\reg_module/_02832_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10107_  (.A(\reg_module/_02832_ ),
    .B(\reg_module/_02593_ ),
    .Y(\reg_module/_02833_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10108_  (.A(\reg_module/_02825_ ),
    .B(\reg_module/_02833_ ),
    .C(\reg_module/_02760_ ),
    .Y(\reg_module/_02834_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10109_  (.A(\reg_module/_02665_ ),
    .B(\reg_module/gprf[35] ),
    .Y(\reg_module/_02835_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10110_  (.A(\reg_module/gprf[3] ),
    .B(net561),
    .Y(\reg_module/_02836_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10111_  (.A(\reg_module/_02835_ ),
    .B(net469),
    .C(\reg_module/_02836_ ),
    .Y(\reg_module/_02837_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10112_  (.A(\reg_module/_02765_ ),
    .B(\reg_module/gprf[99] ),
    .Y(\reg_module/_02838_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10113_  (.A(\reg_module/gprf[67] ),
    .B(net564),
    .Y(\reg_module/_02839_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10114_  (.A(\reg_module/_02838_ ),
    .B(\reg_module/_02605_ ),
    .C(\reg_module/_02839_ ),
    .Y(\reg_module/_02840_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10115_  (.A(\reg_module/_02837_ ),
    .B(\reg_module/_02840_ ),
    .Y(\reg_module/_02841_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10116_  (.A(\reg_module/_02841_ ),
    .B(net421),
    .Y(\reg_module/_02842_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10117_  (.A(\reg_module/_02610_ ),
    .B(\reg_module/gprf[163] ),
    .Y(\reg_module/_02843_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10118_  (.A(\reg_module/gprf[131] ),
    .B(net565),
    .Y(\reg_module/_02844_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10119_  (.A(\reg_module/_02843_ ),
    .B(net471),
    .C(\reg_module/_02844_ ),
    .Y(\reg_module/_02845_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10120_  (.A(\reg_module/_02615_ ),
    .B(\reg_module/gprf[227] ),
    .Y(\reg_module/_02846_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10121_  (.A(\reg_module/gprf[195] ),
    .B(net565),
    .Y(\reg_module/_02847_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10122_  (.A(\reg_module/_02846_ ),
    .B(\reg_module/_02617_ ),
    .C(\reg_module/_02847_ ),
    .Y(\reg_module/_02848_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10123_  (.A(\reg_module/_02845_ ),
    .B(\reg_module/_02848_ ),
    .Y(\reg_module/_02849_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10124_  (.A(\reg_module/_02849_ ),
    .B(\reg_module/_02621_ ),
    .Y(\reg_module/_02850_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10125_  (.A(\reg_module/_02842_ ),
    .B(\reg_module/_02850_ ),
    .C(net396),
    .Y(\reg_module/_02851_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10126_  (.A(\reg_module/_02834_ ),
    .B(\reg_module/_02851_ ),
    .Y(\reg_module/_02852_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10127_  (.A(\reg_module/_02852_ ),
    .B(net380),
    .Y(\reg_module/_02853_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_10128_  (.A(\reg_module/_02817_ ),
    .B(\reg_module/_02853_ ),
    .Y(\wRs2Data[3] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10129_  (.A(\reg_module/_02493_ ),
    .B(\reg_module/gprf[804] ),
    .Y(\reg_module/_02854_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10130_  (.A(\reg_module/gprf[772] ),
    .B(net584),
    .Y(\reg_module/_02855_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10131_  (.A(\reg_module/_02854_ ),
    .B(net480),
    .C(\reg_module/_02855_ ),
    .Y(\reg_module/_02856_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10132_  (.A(\reg_module/_02499_ ),
    .B(\reg_module/gprf[868] ),
    .Y(\reg_module/_02857_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10133_  (.A(\reg_module/gprf[836] ),
    .B(net580),
    .Y(\reg_module/_02858_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10134_  (.A(\reg_module/_02857_ ),
    .B(\reg_module/_02504_ ),
    .C(\reg_module/_02858_ ),
    .Y(\reg_module/_02859_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10135_  (.A(\reg_module/_02856_ ),
    .B(\reg_module/_02859_ ),
    .Y(\reg_module/_02860_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10136_  (.A(\reg_module/_02860_ ),
    .B(net421),
    .Y(\reg_module/_02861_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10137_  (.A(\reg_module/_02570_ ),
    .X(\reg_module/_02862_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10138_  (.A(\reg_module/_02862_ ),
    .B(\reg_module/gprf[932] ),
    .Y(\reg_module/_02863_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10139_  (.A(\reg_module/gprf[900] ),
    .B(net568),
    .Y(\reg_module/_02864_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10140_  (.A(\reg_module/_02863_ ),
    .B(net472),
    .C(\reg_module/_02864_ ),
    .Y(\reg_module/_02865_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10141_  (.A(\reg_module/_02513_ ),
    .X(\reg_module/_02866_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10142_  (.A(\reg_module/_02866_ ),
    .B(\reg_module/gprf[996] ),
    .Y(\reg_module/_02867_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10143_  (.A(\reg_module/gprf[964] ),
    .B(net568),
    .Y(\reg_module/_02868_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10144_  (.A(\reg_module/_02867_ ),
    .B(\reg_module/_02517_ ),
    .C(\reg_module/_02868_ ),
    .Y(\reg_module/_02869_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10145_  (.A(\reg_module/_02865_ ),
    .B(\reg_module/_02869_ ),
    .Y(\reg_module/_02870_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10146_  (.A(\reg_module/_02870_ ),
    .B(\reg_module/_02714_ ),
    .Y(\reg_module/_02871_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10147_  (.A(\reg_module/_02861_ ),
    .B(\reg_module/_02871_ ),
    .C(\reg_module/_02528_ ),
    .Y(\reg_module/_02872_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10148_  (.A(\reg_module/_02717_ ),
    .B(\reg_module/gprf[676] ),
    .Y(\reg_module/_02873_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10149_  (.A(\reg_module/gprf[644] ),
    .B(net565),
    .Y(\reg_module/_02874_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10150_  (.A(\reg_module/_02873_ ),
    .B(net471),
    .C(\reg_module/_02874_ ),
    .Y(\reg_module/_02875_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10151_  (.A(\reg_module/_02535_ ),
    .X(\reg_module/_02876_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10152_  (.A(\reg_module/_02876_ ),
    .B(\reg_module/gprf[740] ),
    .Y(\reg_module/_02877_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10153_  (.A(\reg_module/gprf[708] ),
    .B(net566),
    .Y(\reg_module/_02878_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10154_  (.A(\reg_module/_02877_ ),
    .B(\reg_module/_02722_ ),
    .C(\reg_module/_02878_ ),
    .Y(\reg_module/_02879_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10155_  (.A(\reg_module/_02875_ ),
    .B(\reg_module/_02879_ ),
    .Y(\reg_module/_02880_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10156_  (.A(\reg_module/_02880_ ),
    .B(\reg_module/_02543_ ),
    .Y(\reg_module/_02881_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10157_  (.A(\reg_module/_02546_ ),
    .B(\reg_module/gprf[548] ),
    .Y(\reg_module/_02882_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10158_  (.A(\reg_module/gprf[516] ),
    .B(net579),
    .Y(\reg_module/_02883_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10159_  (.A(\reg_module/_02882_ ),
    .B(net478),
    .C(\reg_module/_02883_ ),
    .Y(\reg_module/_02884_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10160_  (.A(\reg_module/_02730_ ),
    .B(\reg_module/gprf[612] ),
    .Y(\reg_module/_02885_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10161_  (.A(\reg_module/gprf[580] ),
    .B(net580),
    .Y(\reg_module/_02886_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10162_  (.A(\reg_module/_02885_ ),
    .B(\reg_module/_02554_ ),
    .C(\reg_module/_02886_ ),
    .Y(\reg_module/_02887_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10163_  (.A(\reg_module/_02884_ ),
    .B(\reg_module/_02887_ ),
    .Y(\reg_module/_02888_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10164_  (.A(\reg_module/_02888_ ),
    .B(net426),
    .Y(\reg_module/_02889_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10165_  (.A(\reg_module/_02881_ ),
    .B(\reg_module/_02889_ ),
    .C(net396),
    .Y(\reg_module/_02890_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10166_  (.A(\reg_module/_02872_ ),
    .B(\reg_module/_02890_ ),
    .Y(\reg_module/_02891_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10167_  (.A(\reg_module/_02891_ ),
    .B(\reg_module/_02563_ ),
    .Y(\reg_module/_02892_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10168_  (.A(\reg_module/_02565_ ),
    .X(\reg_module/_02893_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10169_  (.A(\reg_module/_02893_ ),
    .B(\reg_module/gprf[292] ),
    .Y(\reg_module/_02894_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10170_  (.A(\reg_module/gprf[260] ),
    .B(net585),
    .Y(\reg_module/_02895_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10171_  (.A(\reg_module/_02894_ ),
    .B(net480),
    .C(\reg_module/_02895_ ),
    .Y(\reg_module/_02896_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_10172_  (.A(\reg_module/_02497_ ),
    .X(\reg_module/_02897_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10173_  (.A(\reg_module/_02897_ ),
    .X(\reg_module/_02898_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10174_  (.A(\reg_module/_02898_ ),
    .B(\reg_module/gprf[356] ),
    .Y(\reg_module/_02899_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10175_  (.A(\reg_module/_02573_ ),
    .X(\reg_module/_02900_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10176_  (.A(\reg_module/gprf[324] ),
    .B(net580),
    .Y(\reg_module/_02901_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10177_  (.A(\reg_module/_02899_ ),
    .B(\reg_module/_02900_ ),
    .C(\reg_module/_02901_ ),
    .Y(\reg_module/_02902_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10178_  (.A(\reg_module/_02896_ ),
    .B(\reg_module/_02902_ ),
    .Y(\reg_module/_02903_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10179_  (.A(\reg_module/_02903_ ),
    .B(net426),
    .Y(\reg_module/_02904_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10180_  (.A(\reg_module/_02750_ ),
    .B(\reg_module/gprf[420] ),
    .Y(\reg_module/_02905_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10181_  (.A(\reg_module/gprf[388] ),
    .B(net563),
    .Y(\reg_module/_02906_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10182_  (.A(\reg_module/_02905_ ),
    .B(net470),
    .C(\reg_module/_02906_ ),
    .Y(\reg_module/_02907_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10183_  (.A(\reg_module/_02550_ ),
    .X(\reg_module/_02908_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10184_  (.A(\reg_module/_02908_ ),
    .B(\reg_module/gprf[484] ),
    .Y(\reg_module/_02909_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10185_  (.A(\reg_module/gprf[452] ),
    .B(net563),
    .Y(\reg_module/_02910_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10186_  (.A(\reg_module/_02909_ ),
    .B(\reg_module/_02755_ ),
    .C(\reg_module/_02910_ ),
    .Y(\reg_module/_02911_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10187_  (.A(\reg_module/_02907_ ),
    .B(\reg_module/_02911_ ),
    .Y(\reg_module/_02912_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10188_  (.A(\reg_module/_02912_ ),
    .B(\reg_module/_02593_ ),
    .Y(\reg_module/_02913_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10189_  (.A(\reg_module/_02904_ ),
    .B(\reg_module/_02913_ ),
    .C(\reg_module/_02760_ ),
    .Y(\reg_module/_02914_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10190_  (.A(\reg_module/_02898_ ),
    .B(\reg_module/gprf[36] ),
    .Y(\reg_module/_02915_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10191_  (.A(\reg_module/gprf[4] ),
    .B(net581),
    .Y(\reg_module/_02916_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10192_  (.A(\reg_module/_02915_ ),
    .B(net479),
    .C(\reg_module/_02916_ ),
    .Y(\reg_module/_02917_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10193_  (.A(\reg_module/_02765_ ),
    .B(\reg_module/gprf[100] ),
    .Y(\reg_module/_02918_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10194_  (.A(\reg_module/_02604_ ),
    .X(\reg_module/_02919_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10195_  (.A(\reg_module/gprf[68] ),
    .B(net581),
    .Y(\reg_module/_02920_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10196_  (.A(\reg_module/_02918_ ),
    .B(\reg_module/_02919_ ),
    .C(\reg_module/_02920_ ),
    .Y(\reg_module/_02921_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10197_  (.A(\reg_module/_02917_ ),
    .B(\reg_module/_02921_ ),
    .Y(\reg_module/_02922_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10198_  (.A(\reg_module/_02922_ ),
    .B(net426),
    .Y(\reg_module/_02923_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10199_  (.A(\reg_module/_02610_ ),
    .B(\reg_module/gprf[164] ),
    .Y(\reg_module/_02924_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10200_  (.A(\reg_module/gprf[132] ),
    .B(net579),
    .Y(\reg_module/_02925_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10201_  (.A(\reg_module/_02924_ ),
    .B(net478),
    .C(\reg_module/_02925_ ),
    .Y(\reg_module/_02926_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10202_  (.A(\reg_module/_02615_ ),
    .B(\reg_module/gprf[228] ),
    .Y(\reg_module/_02927_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10203_  (.A(\reg_module/_02502_ ),
    .X(\reg_module/_02928_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10204_  (.A(\reg_module/gprf[196] ),
    .B(net579),
    .Y(\reg_module/_02929_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10205_  (.A(\reg_module/_02927_ ),
    .B(\reg_module/_02928_ ),
    .C(\reg_module/_02929_ ),
    .Y(\reg_module/_02930_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10206_  (.A(\reg_module/_02926_ ),
    .B(\reg_module/_02930_ ),
    .Y(\reg_module/_02931_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10207_  (.A(\reg_module/_02931_ ),
    .B(\reg_module/_02621_ ),
    .Y(\reg_module/_02932_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10208_  (.A(\reg_module/_02923_ ),
    .B(\reg_module/_02932_ ),
    .C(net404),
    .Y(\reg_module/_02933_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10209_  (.A(\reg_module/_02914_ ),
    .B(\reg_module/_02933_ ),
    .Y(\reg_module/_02934_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10210_  (.A(\reg_module/_02934_ ),
    .B(net380),
    .Y(\reg_module/_02935_ ));
 sky130_fd_sc_hd__nand2_4 \reg_module/_10211_  (.A(\reg_module/_02892_ ),
    .B(\reg_module/_02935_ ),
    .Y(\wRs2Data[4] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10212_  (.A(\reg_module/_02493_ ),
    .B(\reg_module/gprf[549] ),
    .Y(\reg_module/_02936_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10213_  (.A(\reg_module/gprf[517] ),
    .B(net579),
    .Y(\reg_module/_02937_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10214_  (.A(\reg_module/_02936_ ),
    .B(net478),
    .C(\reg_module/_02937_ ),
    .Y(\reg_module/_02938_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10215_  (.A(\reg_module/_02499_ ),
    .B(\reg_module/gprf[613] ),
    .Y(\reg_module/_02939_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10216_  (.A(\reg_module/gprf[581] ),
    .B(net580),
    .Y(\reg_module/_02940_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10217_  (.A(\reg_module/_02939_ ),
    .B(\reg_module/_02504_ ),
    .C(\reg_module/_02940_ ),
    .Y(\reg_module/_02941_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10218_  (.A(\reg_module/_02938_ ),
    .B(\reg_module/_02941_ ),
    .Y(\reg_module/_02942_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10219_  (.A(\reg_module/_02942_ ),
    .B(net422),
    .Y(\reg_module/_02943_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10220_  (.A(\reg_module/_02862_ ),
    .B(\reg_module/gprf[677] ),
    .Y(\reg_module/_02944_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10221_  (.A(\reg_module/gprf[645] ),
    .B(net566),
    .Y(\reg_module/_02945_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10222_  (.A(\reg_module/_02944_ ),
    .B(net471),
    .C(\reg_module/_02945_ ),
    .Y(\reg_module/_02946_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10223_  (.A(\reg_module/_02866_ ),
    .B(\reg_module/gprf[741] ),
    .Y(\reg_module/_02947_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10224_  (.A(\reg_module/gprf[709] ),
    .B(net568),
    .Y(\reg_module/_02948_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10225_  (.A(\reg_module/_02947_ ),
    .B(\reg_module/_02517_ ),
    .C(\reg_module/_02948_ ),
    .Y(\reg_module/_02949_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10226_  (.A(\reg_module/_02946_ ),
    .B(\reg_module/_02949_ ),
    .Y(\reg_module/_02950_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10227_  (.A(\reg_module/_02950_ ),
    .B(\reg_module/_02714_ ),
    .Y(\reg_module/_02951_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10228_  (.A(\reg_module/_02943_ ),
    .B(\reg_module/_02951_ ),
    .C(net396),
    .Y(\reg_module/_02952_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10229_  (.A(\reg_module/_02717_ ),
    .B(\reg_module/gprf[805] ),
    .Y(\reg_module/_02953_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10230_  (.A(\reg_module/gprf[773] ),
    .B(net573),
    .Y(\reg_module/_02954_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10231_  (.A(\reg_module/_02953_ ),
    .B(net475),
    .C(\reg_module/_02954_ ),
    .Y(\reg_module/_02955_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10232_  (.A(\reg_module/_02876_ ),
    .B(\reg_module/gprf[869] ),
    .Y(\reg_module/_02956_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10233_  (.A(\reg_module/gprf[837] ),
    .B(net567),
    .Y(\reg_module/_02957_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10234_  (.A(\reg_module/_02956_ ),
    .B(\reg_module/_02722_ ),
    .C(\reg_module/_02957_ ),
    .Y(\reg_module/_02958_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10235_  (.A(\reg_module/_02955_ ),
    .B(\reg_module/_02958_ ),
    .Y(\reg_module/_02959_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10236_  (.A(\reg_module/_02959_ ),
    .B(net422),
    .Y(\reg_module/_02960_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10237_  (.A(\reg_module/_02546_ ),
    .B(\reg_module/gprf[933] ),
    .Y(\reg_module/_02961_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10238_  (.A(\reg_module/gprf[901] ),
    .B(net568),
    .Y(\reg_module/_02962_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10239_  (.A(\reg_module/_02961_ ),
    .B(net472),
    .C(\reg_module/_02962_ ),
    .Y(\reg_module/_02963_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10240_  (.A(\reg_module/_02730_ ),
    .B(\reg_module/gprf[997] ),
    .Y(\reg_module/_02964_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10241_  (.A(\reg_module/gprf[965] ),
    .B(net567),
    .Y(\reg_module/_02965_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10242_  (.A(\reg_module/_02964_ ),
    .B(\reg_module/_02554_ ),
    .C(\reg_module/_02965_ ),
    .Y(\reg_module/_02966_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10243_  (.A(\reg_module/_02963_ ),
    .B(\reg_module/_02966_ ),
    .Y(\reg_module/_02967_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10244_  (.A(\reg_module/_02967_ ),
    .B(\reg_module/_02736_ ),
    .Y(\reg_module/_02968_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10245_  (.A(\reg_module/_02960_ ),
    .B(\reg_module/_02968_ ),
    .C(\reg_module/_02738_ ),
    .Y(\reg_module/_02969_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10246_  (.A(\reg_module/_02952_ ),
    .B(\reg_module/_02969_ ),
    .Y(\reg_module/_02970_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10247_  (.A(\reg_module/_02970_ ),
    .B(\reg_module/_02563_ ),
    .Y(\reg_module/_02971_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10248_  (.A(\reg_module/_02893_ ),
    .B(\reg_module/gprf[293] ),
    .Y(\reg_module/_02972_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10249_  (.A(\reg_module/gprf[261] ),
    .B(net581),
    .Y(\reg_module/_02973_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10250_  (.A(\reg_module/_02972_ ),
    .B(net478),
    .C(\reg_module/_02973_ ),
    .Y(\reg_module/_02974_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10251_  (.A(\reg_module/_02898_ ),
    .B(\reg_module/gprf[357] ),
    .Y(\reg_module/_02975_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10252_  (.A(\reg_module/gprf[325] ),
    .B(net580),
    .Y(\reg_module/_02976_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10253_  (.A(\reg_module/_02975_ ),
    .B(\reg_module/_02900_ ),
    .C(\reg_module/_02976_ ),
    .Y(\reg_module/_02977_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10254_  (.A(\reg_module/_02974_ ),
    .B(\reg_module/_02977_ ),
    .Y(\reg_module/_02978_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10255_  (.A(\reg_module/_02978_ ),
    .B(net426),
    .Y(\reg_module/_02979_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10256_  (.A(\reg_module/_02750_ ),
    .B(\reg_module/gprf[421] ),
    .Y(\reg_module/_02980_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10257_  (.A(\reg_module/gprf[389] ),
    .B(net563),
    .Y(\reg_module/_02981_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10258_  (.A(\reg_module/_02980_ ),
    .B(net470),
    .C(\reg_module/_02981_ ),
    .Y(\reg_module/_02982_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10259_  (.A(\reg_module/_02908_ ),
    .B(\reg_module/gprf[485] ),
    .Y(\reg_module/_02983_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10260_  (.A(\reg_module/gprf[453] ),
    .B(net563),
    .Y(\reg_module/_02984_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10261_  (.A(\reg_module/_02983_ ),
    .B(\reg_module/_02755_ ),
    .C(\reg_module/_02984_ ),
    .Y(\reg_module/_02985_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10262_  (.A(\reg_module/_02982_ ),
    .B(\reg_module/_02985_ ),
    .Y(\reg_module/_02986_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10263_  (.A(\reg_module/_02986_ ),
    .B(\reg_module/_02593_ ),
    .Y(\reg_module/_02987_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10264_  (.A(\reg_module/_02979_ ),
    .B(\reg_module/_02987_ ),
    .C(\reg_module/_02760_ ),
    .Y(\reg_module/_02988_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10265_  (.A(\reg_module/_02898_ ),
    .B(\reg_module/gprf[37] ),
    .Y(\reg_module/_02989_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10266_  (.A(\reg_module/gprf[5] ),
    .B(net583),
    .Y(\reg_module/_02990_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10267_  (.A(\reg_module/_02989_ ),
    .B(net479),
    .C(\reg_module/_02990_ ),
    .Y(\reg_module/_02991_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10268_  (.A(\reg_module/_02765_ ),
    .B(\reg_module/gprf[101] ),
    .Y(\reg_module/_02992_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10269_  (.A(\reg_module/gprf[69] ),
    .B(net583),
    .Y(\reg_module/_02993_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10270_  (.A(\reg_module/_02992_ ),
    .B(\reg_module/_02919_ ),
    .C(\reg_module/_02993_ ),
    .Y(\reg_module/_02994_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10271_  (.A(\reg_module/_02991_ ),
    .B(\reg_module/_02994_ ),
    .Y(\reg_module/_02995_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10272_  (.A(\reg_module/_02995_ ),
    .B(net426),
    .Y(\reg_module/_02996_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10273_  (.A(\reg_module/_02610_ ),
    .B(\reg_module/gprf[165] ),
    .Y(\reg_module/_02997_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10274_  (.A(\reg_module/gprf[133] ),
    .B(net579),
    .Y(\reg_module/_02998_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10275_  (.A(\reg_module/_02997_ ),
    .B(net478),
    .C(\reg_module/_02998_ ),
    .Y(\reg_module/_02999_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10276_  (.A(\reg_module/_02615_ ),
    .B(\reg_module/gprf[229] ),
    .Y(\reg_module/_03000_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10277_  (.A(\reg_module/gprf[197] ),
    .B(net582),
    .Y(\reg_module/_03001_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10278_  (.A(\reg_module/_03000_ ),
    .B(\reg_module/_02928_ ),
    .C(\reg_module/_03001_ ),
    .Y(\reg_module/_03002_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10279_  (.A(\reg_module/_02999_ ),
    .B(\reg_module/_03002_ ),
    .Y(\reg_module/_03003_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10280_  (.A(\reg_module/_03003_ ),
    .B(\reg_module/_02621_ ),
    .Y(\reg_module/_03004_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10281_  (.A(\reg_module/_02996_ ),
    .B(\reg_module/_03004_ ),
    .C(net404),
    .Y(\reg_module/_03005_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10282_  (.A(\reg_module/_02988_ ),
    .B(\reg_module/_03005_ ),
    .Y(\reg_module/_03006_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10283_  (.A(\reg_module/_03006_ ),
    .B(net380),
    .Y(\reg_module/_03007_ ));
 sky130_fd_sc_hd__nand2_4 \reg_module/_10284_  (.A(\reg_module/_02971_ ),
    .B(\reg_module/_03007_ ),
    .Y(\wRs2Data[5] ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10285_  (.A(\reg_module/_02492_ ),
    .X(\reg_module/_03008_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10286_  (.A(\reg_module/_03008_ ),
    .B(\reg_module/gprf[806] ),
    .Y(\reg_module/_03009_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10287_  (.A(\reg_module/gprf[774] ),
    .B(net584),
    .Y(\reg_module/_03010_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10288_  (.A(\reg_module/_03009_ ),
    .B(net480),
    .C(\reg_module/_03010_ ),
    .Y(\reg_module/_03011_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10289_  (.A(\reg_module/_02498_ ),
    .X(\reg_module/_03012_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10290_  (.A(\reg_module/_03012_ ),
    .B(\reg_module/gprf[870] ),
    .Y(\reg_module/_03013_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10291_  (.A(\reg_module/_02503_ ),
    .X(\reg_module/_03014_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10292_  (.A(\reg_module/gprf[838] ),
    .B(net584),
    .Y(\reg_module/_03015_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10293_  (.A(\reg_module/_03013_ ),
    .B(\reg_module/_03014_ ),
    .C(\reg_module/_03015_ ),
    .Y(\reg_module/_03016_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10294_  (.A(\reg_module/_03011_ ),
    .B(\reg_module/_03016_ ),
    .Y(\reg_module/_03017_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10295_  (.A(\reg_module/_03017_ ),
    .B(net424),
    .Y(\reg_module/_03018_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10296_  (.A(\reg_module/_02862_ ),
    .B(\reg_module/gprf[934] ),
    .Y(\reg_module/_03019_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10297_  (.A(\reg_module/gprf[902] ),
    .B(net575),
    .Y(\reg_module/_03020_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10298_  (.A(\reg_module/_03019_ ),
    .B(net476),
    .C(\reg_module/_03020_ ),
    .Y(\reg_module/_03021_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10299_  (.A(\reg_module/_02866_ ),
    .B(\reg_module/gprf[998] ),
    .Y(\reg_module/_03022_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10300_  (.A(\reg_module/_02516_ ),
    .X(\reg_module/_03023_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10301_  (.A(\reg_module/gprf[966] ),
    .B(net572),
    .Y(\reg_module/_03024_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10302_  (.A(\reg_module/_03022_ ),
    .B(\reg_module/_03023_ ),
    .C(\reg_module/_03024_ ),
    .Y(\reg_module/_03025_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10303_  (.A(\reg_module/_03021_ ),
    .B(\reg_module/_03025_ ),
    .Y(\reg_module/_03026_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10304_  (.A(\reg_module/_03026_ ),
    .B(\reg_module/_02714_ ),
    .Y(\reg_module/_03027_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10305_  (.A(\reg_module/_03018_ ),
    .B(\reg_module/_03027_ ),
    .C(\reg_module/_02528_ ),
    .Y(\reg_module/_03028_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10306_  (.A(\reg_module/_02717_ ),
    .B(\reg_module/gprf[678] ),
    .Y(\reg_module/_03029_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10307_  (.A(\reg_module/gprf[646] ),
    .B(net573),
    .Y(\reg_module/_03030_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10308_  (.A(\reg_module/_03029_ ),
    .B(net475),
    .C(\reg_module/_03030_ ),
    .Y(\reg_module/_03031_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10309_  (.A(\reg_module/_02876_ ),
    .B(\reg_module/gprf[742] ),
    .Y(\reg_module/_03032_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10310_  (.A(\reg_module/gprf[710] ),
    .B(net573),
    .Y(\reg_module/_03033_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10311_  (.A(\reg_module/_03032_ ),
    .B(\reg_module/_02722_ ),
    .C(\reg_module/_03033_ ),
    .Y(\reg_module/_03034_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10312_  (.A(\reg_module/_03031_ ),
    .B(\reg_module/_03034_ ),
    .Y(\reg_module/_03035_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10313_  (.A(\reg_module/_03035_ ),
    .B(\reg_module/_02543_ ),
    .Y(\reg_module/_03036_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10314_  (.A(\reg_module/_02545_ ),
    .X(\reg_module/_03037_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10315_  (.A(\reg_module/_03037_ ),
    .B(\reg_module/gprf[550] ),
    .Y(\reg_module/_03038_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10316_  (.A(\reg_module/gprf[518] ),
    .B(net589),
    .Y(\reg_module/_03039_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10317_  (.A(\reg_module/_03038_ ),
    .B(net481),
    .C(\reg_module/_03039_ ),
    .Y(\reg_module/_03040_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10318_  (.A(\reg_module/_02730_ ),
    .B(\reg_module/gprf[614] ),
    .Y(\reg_module/_03041_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10319_  (.A(\reg_module/_02553_ ),
    .X(\reg_module/_03042_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10320_  (.A(\reg_module/gprf[582] ),
    .B(net590),
    .Y(\reg_module/_03043_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10321_  (.A(\reg_module/_03041_ ),
    .B(\reg_module/_03042_ ),
    .C(\reg_module/_03043_ ),
    .Y(\reg_module/_03044_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10322_  (.A(\reg_module/_03040_ ),
    .B(\reg_module/_03044_ ),
    .Y(\reg_module/_03045_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10323_  (.A(\reg_module/_03045_ ),
    .B(net425),
    .Y(\reg_module/_03046_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10324_  (.A(\reg_module/_03036_ ),
    .B(\reg_module/_03046_ ),
    .C(net397),
    .Y(\reg_module/_03047_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10325_  (.A(\reg_module/_03028_ ),
    .B(\reg_module/_03047_ ),
    .Y(\reg_module/_03048_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10326_  (.A(\reg_module/_02562_ ),
    .X(\reg_module/_03049_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10327_  (.A(\reg_module/_03048_ ),
    .B(\reg_module/_03049_ ),
    .Y(\reg_module/_03050_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10328_  (.A(\reg_module/_02893_ ),
    .B(\reg_module/gprf[294] ),
    .Y(\reg_module/_03051_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10329_  (.A(\reg_module/gprf[262] ),
    .B(net585),
    .Y(\reg_module/_03052_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10330_  (.A(\reg_module/_03051_ ),
    .B(net480),
    .C(\reg_module/_03052_ ),
    .Y(\reg_module/_03053_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10331_  (.A(\reg_module/_02898_ ),
    .B(\reg_module/gprf[358] ),
    .Y(\reg_module/_03054_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10332_  (.A(\reg_module/gprf[326] ),
    .B(net584),
    .Y(\reg_module/_03055_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10333_  (.A(\reg_module/_03054_ ),
    .B(\reg_module/_02900_ ),
    .C(\reg_module/_03055_ ),
    .Y(\reg_module/_03056_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10334_  (.A(\reg_module/_03053_ ),
    .B(\reg_module/_03056_ ),
    .Y(\reg_module/_03057_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10335_  (.A(\reg_module/_03057_ ),
    .B(net424),
    .Y(\reg_module/_03058_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10336_  (.A(\reg_module/_02750_ ),
    .B(\reg_module/gprf[422] ),
    .Y(\reg_module/_03059_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10337_  (.A(\reg_module/gprf[390] ),
    .B(net570),
    .Y(\reg_module/_03060_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10338_  (.A(\reg_module/_03059_ ),
    .B(net474),
    .C(\reg_module/_03060_ ),
    .Y(\reg_module/_03061_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10339_  (.A(\reg_module/_02908_ ),
    .B(\reg_module/gprf[486] ),
    .Y(\reg_module/_03062_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10340_  (.A(\reg_module/gprf[454] ),
    .B(net570),
    .Y(\reg_module/_03063_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10341_  (.A(\reg_module/_03062_ ),
    .B(\reg_module/_02755_ ),
    .C(\reg_module/_03063_ ),
    .Y(\reg_module/_03064_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10342_  (.A(\reg_module/_03061_ ),
    .B(\reg_module/_03064_ ),
    .Y(\reg_module/_03065_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10343_  (.A(\reg_module/_02735_ ),
    .X(\reg_module/_03066_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10344_  (.A(\reg_module/_03065_ ),
    .B(\reg_module/_03066_ ),
    .Y(\reg_module/_03067_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10345_  (.A(\reg_module/_03058_ ),
    .B(\reg_module/_03067_ ),
    .C(\reg_module/_02760_ ),
    .Y(\reg_module/_03068_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10346_  (.A(\reg_module/_02898_ ),
    .B(\reg_module/gprf[38] ),
    .Y(\reg_module/_03069_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10347_  (.A(\reg_module/gprf[6] ),
    .B(net587),
    .Y(\reg_module/_03070_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10348_  (.A(\reg_module/_03069_ ),
    .B(net482),
    .C(\reg_module/_03070_ ),
    .Y(\reg_module/_03071_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10349_  (.A(\reg_module/_02765_ ),
    .B(\reg_module/gprf[102] ),
    .Y(\reg_module/_03072_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10350_  (.A(\reg_module/gprf[70] ),
    .B(net588),
    .Y(\reg_module/_03073_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10351_  (.A(\reg_module/_03072_ ),
    .B(\reg_module/_02919_ ),
    .C(\reg_module/_03073_ ),
    .Y(\reg_module/_03074_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10352_  (.A(\reg_module/_03071_ ),
    .B(\reg_module/_03074_ ),
    .Y(\reg_module/_03075_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10353_  (.A(\reg_module/_03075_ ),
    .B(net425),
    .Y(\reg_module/_03076_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10354_  (.A(\reg_module/_02584_ ),
    .X(\reg_module/_03077_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10355_  (.A(\reg_module/_03077_ ),
    .B(\reg_module/gprf[166] ),
    .Y(\reg_module/_03078_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10356_  (.A(\reg_module/gprf[134] ),
    .B(net592),
    .Y(\reg_module/_03079_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10357_  (.A(\reg_module/_03078_ ),
    .B(net479),
    .C(\reg_module/_03079_ ),
    .Y(\reg_module/_03080_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10358_  (.A(\reg_module/_02614_ ),
    .X(\reg_module/_03081_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10359_  (.A(\reg_module/_03081_ ),
    .B(\reg_module/gprf[230] ),
    .Y(\reg_module/_03082_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10360_  (.A(\reg_module/gprf[198] ),
    .B(net583),
    .Y(\reg_module/_03083_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10361_  (.A(\reg_module/_03082_ ),
    .B(\reg_module/_02928_ ),
    .C(\reg_module/_03083_ ),
    .Y(\reg_module/_03084_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10362_  (.A(\reg_module/_03080_ ),
    .B(\reg_module/_03084_ ),
    .Y(\reg_module/_03085_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_10363_  (.A(\reg_module/_02522_ ),
    .X(\reg_module/_03086_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10364_  (.A(\reg_module/_03085_ ),
    .B(\reg_module/_03086_ ),
    .Y(\reg_module/_03087_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10365_  (.A(\reg_module/_03076_ ),
    .B(\reg_module/_03087_ ),
    .C(net398),
    .Y(\reg_module/_03088_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10366_  (.A(\reg_module/_03068_ ),
    .B(\reg_module/_03088_ ),
    .Y(\reg_module/_03089_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10367_  (.A(\reg_module/_03089_ ),
    .B(net380),
    .Y(\reg_module/_03090_ ));
 sky130_fd_sc_hd__nand2_4 \reg_module/_10368_  (.A(\reg_module/_03050_ ),
    .B(\reg_module/_03090_ ),
    .Y(\wRs2Data[6] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10369_  (.A(\reg_module/_03008_ ),
    .B(\reg_module/gprf[807] ),
    .Y(\reg_module/_03091_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10370_  (.A(\reg_module/gprf[775] ),
    .B(net591),
    .Y(\reg_module/_03092_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10371_  (.A(\reg_module/_03091_ ),
    .B(net483),
    .C(\reg_module/_03092_ ),
    .Y(\reg_module/_03093_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10372_  (.A(\reg_module/_03012_ ),
    .B(\reg_module/gprf[871] ),
    .Y(\reg_module/_03094_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10373_  (.A(\reg_module/gprf[839] ),
    .B(net585),
    .Y(\reg_module/_03095_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10374_  (.A(\reg_module/_03094_ ),
    .B(\reg_module/_03014_ ),
    .C(\reg_module/_03095_ ),
    .Y(\reg_module/_03096_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10375_  (.A(\reg_module/_03093_ ),
    .B(\reg_module/_03096_ ),
    .Y(\reg_module/_03097_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10376_  (.A(\reg_module/_03097_ ),
    .B(net424),
    .Y(\reg_module/_03098_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10377_  (.A(\reg_module/_02862_ ),
    .B(\reg_module/gprf[935] ),
    .Y(\reg_module/_03099_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10378_  (.A(\reg_module/gprf[903] ),
    .B(net574),
    .Y(\reg_module/_03100_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10379_  (.A(\reg_module/_03099_ ),
    .B(net475),
    .C(\reg_module/_03100_ ),
    .Y(\reg_module/_03101_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10380_  (.A(\reg_module/_02866_ ),
    .B(\reg_module/gprf[999] ),
    .Y(\reg_module/_03102_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10381_  (.A(\reg_module/gprf[967] ),
    .B(net574),
    .Y(\reg_module/_03103_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10382_  (.A(\reg_module/_03102_ ),
    .B(\reg_module/_03023_ ),
    .C(\reg_module/_03103_ ),
    .Y(\reg_module/_03104_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10383_  (.A(\reg_module/_03101_ ),
    .B(\reg_module/_03104_ ),
    .Y(\reg_module/_03105_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10384_  (.A(\reg_module/_03105_ ),
    .B(\reg_module/_02714_ ),
    .Y(\reg_module/_03106_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10385_  (.A(\reg_module/_03098_ ),
    .B(\reg_module/_03106_ ),
    .C(\reg_module/_02528_ ),
    .Y(\reg_module/_03107_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10386_  (.A(\reg_module/_02717_ ),
    .B(\reg_module/gprf[679] ),
    .Y(\reg_module/_03108_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10387_  (.A(\reg_module/gprf[647] ),
    .B(net572),
    .Y(\reg_module/_03109_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10388_  (.A(\reg_module/_03108_ ),
    .B(net475),
    .C(\reg_module/_03109_ ),
    .Y(\reg_module/_03110_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10389_  (.A(\reg_module/_02876_ ),
    .B(\reg_module/gprf[743] ),
    .Y(\reg_module/_03111_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10390_  (.A(\reg_module/gprf[711] ),
    .B(net572),
    .Y(\reg_module/_03112_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10391_  (.A(\reg_module/_03111_ ),
    .B(\reg_module/_02722_ ),
    .C(\reg_module/_03112_ ),
    .Y(\reg_module/_03113_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10392_  (.A(\reg_module/_03110_ ),
    .B(\reg_module/_03113_ ),
    .Y(\reg_module/_03114_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10393_  (.A(\reg_module/_03114_ ),
    .B(\reg_module/_02543_ ),
    .Y(\reg_module/_03115_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10394_  (.A(\reg_module/_03037_ ),
    .B(\reg_module/gprf[551] ),
    .Y(\reg_module/_03116_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10395_  (.A(\reg_module/gprf[519] ),
    .B(net590),
    .Y(\reg_module/_03117_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10396_  (.A(\reg_module/_03116_ ),
    .B(net483),
    .C(\reg_module/_03117_ ),
    .Y(\reg_module/_03118_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10397_  (.A(\reg_module/_02730_ ),
    .B(\reg_module/gprf[615] ),
    .Y(\reg_module/_03119_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10398_  (.A(\reg_module/gprf[583] ),
    .B(net589),
    .Y(\reg_module/_03120_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10399_  (.A(\reg_module/_03119_ ),
    .B(\reg_module/_03042_ ),
    .C(\reg_module/_03120_ ),
    .Y(\reg_module/_03121_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10400_  (.A(\reg_module/_03118_ ),
    .B(\reg_module/_03121_ ),
    .Y(\reg_module/_03122_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10401_  (.A(\reg_module/_03122_ ),
    .B(net425),
    .Y(\reg_module/_03123_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10402_  (.A(\reg_module/_03115_ ),
    .B(\reg_module/_03123_ ),
    .C(net397),
    .Y(\reg_module/_03124_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10403_  (.A(\reg_module/_03107_ ),
    .B(\reg_module/_03124_ ),
    .Y(\reg_module/_03125_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10404_  (.A(\reg_module/_03125_ ),
    .B(\reg_module/_03049_ ),
    .Y(\reg_module/_03126_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10405_  (.A(\reg_module/_02893_ ),
    .B(\reg_module/gprf[295] ),
    .Y(\reg_module/_03127_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10406_  (.A(\reg_module/gprf[263] ),
    .B(net584),
    .Y(\reg_module/_03128_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10407_  (.A(\reg_module/_03127_ ),
    .B(net480),
    .C(\reg_module/_03128_ ),
    .Y(\reg_module/_03129_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10408_  (.A(\reg_module/_02897_ ),
    .X(\reg_module/_03130_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10409_  (.A(\reg_module/_03130_ ),
    .B(\reg_module/gprf[359] ),
    .Y(\reg_module/_03131_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10410_  (.A(\reg_module/gprf[327] ),
    .B(net584),
    .Y(\reg_module/_03132_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10411_  (.A(\reg_module/_03131_ ),
    .B(\reg_module/_02900_ ),
    .C(\reg_module/_03132_ ),
    .Y(\reg_module/_03133_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10412_  (.A(\reg_module/_03129_ ),
    .B(\reg_module/_03133_ ),
    .Y(\reg_module/_03134_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10413_  (.A(\reg_module/_03134_ ),
    .B(net424),
    .Y(\reg_module/_03135_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10414_  (.A(\reg_module/_02750_ ),
    .B(\reg_module/gprf[423] ),
    .Y(\reg_module/_03136_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10415_  (.A(\reg_module/gprf[391] ),
    .B(net571),
    .Y(\reg_module/_03137_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10416_  (.A(\reg_module/_03136_ ),
    .B(net474),
    .C(\reg_module/_03137_ ),
    .Y(\reg_module/_03138_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10417_  (.A(\reg_module/_02908_ ),
    .B(\reg_module/gprf[487] ),
    .Y(\reg_module/_03139_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10418_  (.A(\reg_module/gprf[455] ),
    .B(net577),
    .Y(\reg_module/_03140_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10419_  (.A(\reg_module/_03139_ ),
    .B(\reg_module/_02755_ ),
    .C(\reg_module/_03140_ ),
    .Y(\reg_module/_03141_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10420_  (.A(\reg_module/_03138_ ),
    .B(\reg_module/_03141_ ),
    .Y(\reg_module/_03142_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10421_  (.A(\reg_module/_03142_ ),
    .B(\reg_module/_03066_ ),
    .Y(\reg_module/_03143_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10422_  (.A(\reg_module/_03135_ ),
    .B(\reg_module/_03143_ ),
    .C(\reg_module/_02760_ ),
    .Y(\reg_module/_03144_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10423_  (.A(\reg_module/_03130_ ),
    .B(\reg_module/gprf[39] ),
    .Y(\reg_module/_03145_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10424_  (.A(\reg_module/gprf[7] ),
    .B(net589),
    .Y(\reg_module/_03146_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10425_  (.A(\reg_module/_03145_ ),
    .B(net481),
    .C(\reg_module/_03146_ ),
    .Y(\reg_module/_03147_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10426_  (.A(\reg_module/_02765_ ),
    .B(\reg_module/gprf[103] ),
    .Y(\reg_module/_03148_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10427_  (.A(\reg_module/gprf[71] ),
    .B(net589),
    .Y(\reg_module/_03149_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10428_  (.A(\reg_module/_03148_ ),
    .B(\reg_module/_02919_ ),
    .C(\reg_module/_03149_ ),
    .Y(\reg_module/_03150_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10429_  (.A(\reg_module/_03147_ ),
    .B(\reg_module/_03150_ ),
    .Y(\reg_module/_03151_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10430_  (.A(\reg_module/_03151_ ),
    .B(net425),
    .Y(\reg_module/_03152_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10431_  (.A(\reg_module/_03077_ ),
    .B(\reg_module/gprf[167] ),
    .Y(\reg_module/_03153_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10432_  (.A(\reg_module/gprf[135] ),
    .B(net583),
    .Y(\reg_module/_03154_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10433_  (.A(\reg_module/_03153_ ),
    .B(net479),
    .C(\reg_module/_03154_ ),
    .Y(\reg_module/_03155_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10434_  (.A(\reg_module/_03081_ ),
    .B(\reg_module/gprf[231] ),
    .Y(\reg_module/_03156_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10435_  (.A(\reg_module/gprf[199] ),
    .B(net583),
    .Y(\reg_module/_03157_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10436_  (.A(\reg_module/_03156_ ),
    .B(\reg_module/_02928_ ),
    .C(\reg_module/_03157_ ),
    .Y(\reg_module/_03158_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10437_  (.A(\reg_module/_03155_ ),
    .B(\reg_module/_03158_ ),
    .Y(\reg_module/_03159_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10438_  (.A(\reg_module/_03159_ ),
    .B(\reg_module/_03086_ ),
    .Y(\reg_module/_03160_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10439_  (.A(\reg_module/_03152_ ),
    .B(\reg_module/_03160_ ),
    .C(net398),
    .Y(\reg_module/_03161_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10440_  (.A(\reg_module/_03144_ ),
    .B(\reg_module/_03161_ ),
    .Y(\reg_module/_03162_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10441_  (.A(\reg_module/_03162_ ),
    .B(net381),
    .Y(\reg_module/_03163_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_10442_  (.A(\reg_module/_03126_ ),
    .B(\reg_module/_03163_ ),
    .Y(\wRs2Data[7] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10443_  (.A(\reg_module/_03008_ ),
    .B(\reg_module/gprf[552] ),
    .Y(\reg_module/_03164_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10444_  (.A(\reg_module/gprf[520] ),
    .B(net586),
    .Y(\reg_module/_03165_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10445_  (.A(\reg_module/_03164_ ),
    .B(net483),
    .C(\reg_module/_03165_ ),
    .Y(\reg_module/_03166_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10446_  (.A(\reg_module/_03012_ ),
    .B(\reg_module/gprf[616] ),
    .Y(\reg_module/_03167_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10447_  (.A(\reg_module/gprf[584] ),
    .B(net586),
    .Y(\reg_module/_03168_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10448_  (.A(\reg_module/_03167_ ),
    .B(\reg_module/_03014_ ),
    .C(\reg_module/_03168_ ),
    .Y(\reg_module/_03169_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10449_  (.A(\reg_module/_03166_ ),
    .B(\reg_module/_03169_ ),
    .Y(\reg_module/_03170_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10450_  (.A(\reg_module/_03170_ ),
    .B(net423),
    .Y(\reg_module/_03171_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10451_  (.A(\reg_module/_02862_ ),
    .B(\reg_module/gprf[680] ),
    .Y(\reg_module/_03172_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10452_  (.A(\reg_module/gprf[648] ),
    .B(net574),
    .Y(\reg_module/_03173_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10453_  (.A(\reg_module/_03172_ ),
    .B(net476),
    .C(\reg_module/_03173_ ),
    .Y(\reg_module/_03174_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10454_  (.A(\reg_module/_02866_ ),
    .B(\reg_module/gprf[744] ),
    .Y(\reg_module/_03175_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10455_  (.A(\reg_module/gprf[712] ),
    .B(net574),
    .Y(\reg_module/_03176_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10456_  (.A(\reg_module/_03175_ ),
    .B(\reg_module/_03023_ ),
    .C(\reg_module/_03176_ ),
    .Y(\reg_module/_03177_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10457_  (.A(\reg_module/_03174_ ),
    .B(\reg_module/_03177_ ),
    .Y(\reg_module/_03178_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10458_  (.A(\reg_module/_02592_ ),
    .X(\reg_module/_03179_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10459_  (.A(\reg_module/_03178_ ),
    .B(\reg_module/_03179_ ),
    .Y(\reg_module/_03180_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10460_  (.A(\reg_module/_03171_ ),
    .B(\reg_module/_03180_ ),
    .C(net397),
    .Y(\reg_module/_03181_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10461_  (.A(\reg_module/_02530_ ),
    .X(\reg_module/_03182_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10462_  (.A(\reg_module/_03182_ ),
    .B(\reg_module/gprf[808] ),
    .Y(\reg_module/_03183_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10463_  (.A(\reg_module/gprf[776] ),
    .B(net591),
    .Y(\reg_module/_03184_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10464_  (.A(\reg_module/_03183_ ),
    .B(net480),
    .C(\reg_module/_03184_ ),
    .Y(\reg_module/_03185_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10465_  (.A(\reg_module/_02876_ ),
    .B(\reg_module/gprf[872] ),
    .Y(\reg_module/_03186_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10466_  (.A(\reg_module/_02538_ ),
    .X(\reg_module/_03187_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10467_  (.A(\reg_module/gprf[840] ),
    .B(net597),
    .Y(\reg_module/_03188_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10468_  (.A(\reg_module/_03186_ ),
    .B(\reg_module/_03187_ ),
    .C(\reg_module/_03188_ ),
    .Y(\reg_module/_03189_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10469_  (.A(\reg_module/_03185_ ),
    .B(\reg_module/_03189_ ),
    .Y(\reg_module/_03190_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10470_  (.A(\reg_module/_03190_ ),
    .B(net423),
    .Y(\reg_module/_03191_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10471_  (.A(\reg_module/_03037_ ),
    .B(\reg_module/gprf[936] ),
    .Y(\reg_module/_03192_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10472_  (.A(\reg_module/gprf[904] ),
    .B(net574),
    .Y(\reg_module/_03193_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10473_  (.A(\reg_module/_03192_ ),
    .B(net475),
    .C(\reg_module/_03193_ ),
    .Y(\reg_module/_03194_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10474_  (.A(\reg_module/_02614_ ),
    .X(\reg_module/_03195_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10475_  (.A(\reg_module/_03195_ ),
    .B(\reg_module/gprf[1000] ),
    .Y(\reg_module/_03196_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10476_  (.A(\reg_module/gprf[968] ),
    .B(net575),
    .Y(\reg_module/_03197_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10477_  (.A(\reg_module/_03196_ ),
    .B(\reg_module/_03042_ ),
    .C(\reg_module/_03197_ ),
    .Y(\reg_module/_03198_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10478_  (.A(\reg_module/_03194_ ),
    .B(\reg_module/_03198_ ),
    .Y(\reg_module/_03199_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10479_  (.A(\reg_module/_03199_ ),
    .B(\reg_module/_02736_ ),
    .Y(\reg_module/_03200_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10480_  (.A(\reg_module/_03191_ ),
    .B(\reg_module/_03200_ ),
    .C(\reg_module/_02738_ ),
    .Y(\reg_module/_03201_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10481_  (.A(\reg_module/_03181_ ),
    .B(\reg_module/_03201_ ),
    .Y(\reg_module/_03202_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10482_  (.A(\reg_module/_03202_ ),
    .B(\reg_module/_03049_ ),
    .Y(\reg_module/_03203_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10483_  (.A(\reg_module/_02893_ ),
    .B(\reg_module/gprf[296] ),
    .Y(\reg_module/_03204_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10484_  (.A(\reg_module/gprf[264] ),
    .B(net590),
    .Y(\reg_module/_03205_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10485_  (.A(\reg_module/_03204_ ),
    .B(net481),
    .C(\reg_module/_03205_ ),
    .Y(\reg_module/_03206_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10486_  (.A(\reg_module/_03130_ ),
    .B(\reg_module/gprf[360] ),
    .Y(\reg_module/_03207_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10487_  (.A(\reg_module/gprf[328] ),
    .B(net586),
    .Y(\reg_module/_03208_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10488_  (.A(\reg_module/_03207_ ),
    .B(\reg_module/_02900_ ),
    .C(\reg_module/_03208_ ),
    .Y(\reg_module/_03209_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10489_  (.A(\reg_module/_03206_ ),
    .B(\reg_module/_03209_ ),
    .Y(\reg_module/_03210_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10490_  (.A(\reg_module/_03210_ ),
    .B(net424),
    .Y(\reg_module/_03211_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10491_  (.A(\reg_module/_02579_ ),
    .X(\reg_module/_03212_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10492_  (.A(\reg_module/_03212_ ),
    .B(\reg_module/gprf[424] ),
    .Y(\reg_module/_03213_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10493_  (.A(\reg_module/gprf[392] ),
    .B(net571),
    .Y(\reg_module/_03214_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10494_  (.A(\reg_module/_03213_ ),
    .B(net477),
    .C(\reg_module/_03214_ ),
    .Y(\reg_module/_03215_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10495_  (.A(\reg_module/_02908_ ),
    .B(\reg_module/gprf[488] ),
    .Y(\reg_module/_03216_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10496_  (.A(\reg_module/_02587_ ),
    .X(\reg_module/_03217_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10497_  (.A(\reg_module/gprf[456] ),
    .B(net571),
    .Y(\reg_module/_03218_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10498_  (.A(\reg_module/_03216_ ),
    .B(\reg_module/_03217_ ),
    .C(\reg_module/_03218_ ),
    .Y(\reg_module/_03219_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10499_  (.A(\reg_module/_03215_ ),
    .B(\reg_module/_03219_ ),
    .Y(\reg_module/_03220_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10500_  (.A(\reg_module/_03220_ ),
    .B(\reg_module/_03066_ ),
    .Y(\reg_module/_03221_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10501_  (.A(\reg_module/_02595_ ),
    .X(\reg_module/_03222_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10502_  (.A(\reg_module/_03211_ ),
    .B(\reg_module/_03221_ ),
    .C(\reg_module/_03222_ ),
    .Y(\reg_module/_03223_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10503_  (.A(\reg_module/_03130_ ),
    .B(\reg_module/gprf[40] ),
    .Y(\reg_module/_03224_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10504_  (.A(\reg_module/gprf[8] ),
    .B(net590),
    .Y(\reg_module/_03225_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10505_  (.A(\reg_module/_03224_ ),
    .B(net481),
    .C(\reg_module/_03225_ ),
    .Y(\reg_module/_03226_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10506_  (.A(\reg_module/_02601_ ),
    .X(\reg_module/_03227_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10507_  (.A(\reg_module/_03227_ ),
    .B(\reg_module/gprf[104] ),
    .Y(\reg_module/_03228_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10508_  (.A(\reg_module/gprf[72] ),
    .B(net589),
    .Y(\reg_module/_03229_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10509_  (.A(\reg_module/_03228_ ),
    .B(\reg_module/_02919_ ),
    .C(\reg_module/_03229_ ),
    .Y(\reg_module/_03230_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10510_  (.A(\reg_module/_03226_ ),
    .B(\reg_module/_03230_ ),
    .Y(\reg_module/_03231_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10511_  (.A(\reg_module/_03231_ ),
    .B(net425),
    .Y(\reg_module/_03232_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10512_  (.A(\reg_module/_03077_ ),
    .B(\reg_module/gprf[168] ),
    .Y(\reg_module/_03233_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10513_  (.A(\reg_module/gprf[136] ),
    .B(net587),
    .Y(\reg_module/_03234_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10514_  (.A(\reg_module/_03233_ ),
    .B(net482),
    .C(\reg_module/_03234_ ),
    .Y(\reg_module/_03235_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10515_  (.A(\reg_module/_03081_ ),
    .B(\reg_module/gprf[232] ),
    .Y(\reg_module/_03236_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10516_  (.A(\reg_module/gprf[200] ),
    .B(net588),
    .Y(\reg_module/_03237_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10517_  (.A(\reg_module/_03236_ ),
    .B(\reg_module/_02928_ ),
    .C(\reg_module/_03237_ ),
    .Y(\reg_module/_03238_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10518_  (.A(\reg_module/_03235_ ),
    .B(\reg_module/_03238_ ),
    .Y(\reg_module/_03239_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10519_  (.A(\reg_module/_03239_ ),
    .B(\reg_module/_03086_ ),
    .Y(\reg_module/_03240_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10520_  (.A(\reg_module/_03232_ ),
    .B(\reg_module/_03240_ ),
    .C(net398),
    .Y(\reg_module/_03241_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10521_  (.A(\reg_module/_03223_ ),
    .B(\reg_module/_03241_ ),
    .Y(\reg_module/_03242_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10522_  (.A(\reg_module/_03242_ ),
    .B(net381),
    .Y(\reg_module/_03243_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_10523_  (.A(\reg_module/_03203_ ),
    .B(\reg_module/_03243_ ),
    .Y(\wRs2Data[8] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10524_  (.A(\reg_module/_03008_ ),
    .B(\reg_module/gprf[809] ),
    .Y(\reg_module/_03244_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10525_  (.A(\reg_module/gprf[777] ),
    .B(net612),
    .Y(\reg_module/_03245_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10526_  (.A(\reg_module/_03244_ ),
    .B(net494),
    .C(\reg_module/_03245_ ),
    .Y(\reg_module/_03246_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10527_  (.A(\reg_module/_03012_ ),
    .B(\reg_module/gprf[873] ),
    .Y(\reg_module/_03247_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10528_  (.A(\reg_module/gprf[841] ),
    .B(net612),
    .Y(\reg_module/_03248_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10529_  (.A(\reg_module/_03247_ ),
    .B(\reg_module/_03014_ ),
    .C(\reg_module/_03248_ ),
    .Y(\reg_module/_03249_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10530_  (.A(\reg_module/_03246_ ),
    .B(\reg_module/_03249_ ),
    .Y(\reg_module/_03250_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10531_  (.A(\reg_module/_03250_ ),
    .B(net431),
    .Y(\reg_module/_03251_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10532_  (.A(\reg_module/_02862_ ),
    .B(\reg_module/gprf[937] ),
    .Y(\reg_module/_03252_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10533_  (.A(\reg_module/gprf[905] ),
    .B(net596),
    .Y(\reg_module/_03253_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10534_  (.A(\reg_module/_03252_ ),
    .B(net476),
    .C(\reg_module/_03253_ ),
    .Y(\reg_module/_03254_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10535_  (.A(\reg_module/_02866_ ),
    .B(\reg_module/gprf[1001] ),
    .Y(\reg_module/_03255_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10536_  (.A(\reg_module/gprf[969] ),
    .B(net574),
    .Y(\reg_module/_03256_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10537_  (.A(\reg_module/_03255_ ),
    .B(\reg_module/_03023_ ),
    .C(\reg_module/_03256_ ),
    .Y(\reg_module/_03257_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10538_  (.A(\reg_module/_03254_ ),
    .B(\reg_module/_03257_ ),
    .Y(\reg_module/_03258_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10539_  (.A(\reg_module/_03258_ ),
    .B(\reg_module/_03179_ ),
    .Y(\reg_module/_03259_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10540_  (.A(\reg_module/_02527_ ),
    .X(\reg_module/_03260_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10541_  (.A(\reg_module/_03251_ ),
    .B(\reg_module/_03259_ ),
    .C(\reg_module/_03260_ ),
    .Y(\reg_module/_03261_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10542_  (.A(\reg_module/_03182_ ),
    .B(\reg_module/gprf[681] ),
    .Y(\reg_module/_03262_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10543_  (.A(\reg_module/gprf[649] ),
    .B(net575),
    .Y(\reg_module/_03263_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10544_  (.A(\reg_module/_03262_ ),
    .B(net476),
    .C(\reg_module/_03263_ ),
    .Y(\reg_module/_03264_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10545_  (.A(\reg_module/_02876_ ),
    .B(\reg_module/gprf[745] ),
    .Y(\reg_module/_03265_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10546_  (.A(\reg_module/gprf[713] ),
    .B(net597),
    .Y(\reg_module/_03266_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10547_  (.A(\reg_module/_03265_ ),
    .B(\reg_module/_03187_ ),
    .C(\reg_module/_03266_ ),
    .Y(\reg_module/_03267_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10548_  (.A(\reg_module/_03264_ ),
    .B(\reg_module/_03267_ ),
    .Y(\reg_module/_03268_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10549_  (.A(\reg_module/_02523_ ),
    .X(\reg_module/_03269_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10550_  (.A(\reg_module/_03268_ ),
    .B(\reg_module/_03269_ ),
    .Y(\reg_module/_03270_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10551_  (.A(\reg_module/_03037_ ),
    .B(\reg_module/gprf[553] ),
    .Y(\reg_module/_03271_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10552_  (.A(\reg_module/gprf[521] ),
    .B(net615),
    .Y(\reg_module/_03272_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10553_  (.A(\reg_module/_03271_ ),
    .B(net495),
    .C(\reg_module/_03272_ ),
    .Y(\reg_module/_03273_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10554_  (.A(\reg_module/_03195_ ),
    .B(\reg_module/gprf[617] ),
    .Y(\reg_module/_03274_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10555_  (.A(\reg_module/gprf[585] ),
    .B(net616),
    .Y(\reg_module/_03275_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10556_  (.A(\reg_module/_03274_ ),
    .B(\reg_module/_03042_ ),
    .C(\reg_module/_03275_ ),
    .Y(\reg_module/_03276_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10557_  (.A(\reg_module/_03273_ ),
    .B(\reg_module/_03276_ ),
    .Y(\reg_module/_03277_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10558_  (.A(\reg_module/_03277_ ),
    .B(net432),
    .Y(\reg_module/_03278_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10559_  (.A(\reg_module/_03270_ ),
    .B(\reg_module/_03278_ ),
    .C(net399),
    .Y(\reg_module/_03279_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10560_  (.A(\reg_module/_03261_ ),
    .B(\reg_module/_03279_ ),
    .Y(\reg_module/_03280_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10561_  (.A(\reg_module/_03280_ ),
    .B(\reg_module/_03049_ ),
    .Y(\reg_module/_03281_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10562_  (.A(\reg_module/_02893_ ),
    .B(\reg_module/gprf[297] ),
    .Y(\reg_module/_03282_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10563_  (.A(\reg_module/gprf[265] ),
    .B(net590),
    .Y(\reg_module/_03283_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10564_  (.A(\reg_module/_03282_ ),
    .B(net481),
    .C(\reg_module/_03283_ ),
    .Y(\reg_module/_03284_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10565_  (.A(\reg_module/_03130_ ),
    .B(\reg_module/gprf[361] ),
    .Y(\reg_module/_03285_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10566_  (.A(\reg_module/gprf[329] ),
    .B(net586),
    .Y(\reg_module/_03286_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10567_  (.A(\reg_module/_03285_ ),
    .B(\reg_module/_02900_ ),
    .C(\reg_module/_03286_ ),
    .Y(\reg_module/_03287_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10568_  (.A(\reg_module/_03284_ ),
    .B(\reg_module/_03287_ ),
    .Y(\reg_module/_03288_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10569_  (.A(\reg_module/_03288_ ),
    .B(net424),
    .Y(\reg_module/_03289_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10570_  (.A(\reg_module/_03212_ ),
    .B(\reg_module/gprf[425] ),
    .Y(\reg_module/_03290_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10571_  (.A(\reg_module/gprf[393] ),
    .B(net577),
    .Y(\reg_module/_03291_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10572_  (.A(\reg_module/_03290_ ),
    .B(net477),
    .C(\reg_module/_03291_ ),
    .Y(\reg_module/_03292_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10573_  (.A(\reg_module/_02908_ ),
    .B(\reg_module/gprf[489] ),
    .Y(\reg_module/_03293_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10574_  (.A(\reg_module/gprf[457] ),
    .B(net571),
    .Y(\reg_module/_03294_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10575_  (.A(\reg_module/_03293_ ),
    .B(\reg_module/_03217_ ),
    .C(\reg_module/_03294_ ),
    .Y(\reg_module/_03295_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10576_  (.A(\reg_module/_03292_ ),
    .B(\reg_module/_03295_ ),
    .Y(\reg_module/_03296_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10577_  (.A(\reg_module/_03296_ ),
    .B(\reg_module/_03066_ ),
    .Y(\reg_module/_03297_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10578_  (.A(\reg_module/_03289_ ),
    .B(\reg_module/_03297_ ),
    .C(\reg_module/_03222_ ),
    .Y(\reg_module/_03298_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10579_  (.A(\reg_module/_03130_ ),
    .B(\reg_module/gprf[41] ),
    .Y(\reg_module/_03299_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10580_  (.A(\reg_module/gprf[9] ),
    .B(net589),
    .Y(\reg_module/_03300_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10581_  (.A(\reg_module/_03299_ ),
    .B(net481),
    .C(\reg_module/_03300_ ),
    .Y(\reg_module/_03301_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10582_  (.A(\reg_module/_03227_ ),
    .B(\reg_module/gprf[105] ),
    .Y(\reg_module/_03302_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10583_  (.A(\reg_module/gprf[73] ),
    .B(net616),
    .Y(\reg_module/_03303_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10584_  (.A(\reg_module/_03302_ ),
    .B(\reg_module/_02919_ ),
    .C(\reg_module/_03303_ ),
    .Y(\reg_module/_03304_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10585_  (.A(\reg_module/_03301_ ),
    .B(\reg_module/_03304_ ),
    .Y(\reg_module/_03305_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10586_  (.A(\reg_module/_03305_ ),
    .B(net425),
    .Y(\reg_module/_03306_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10587_  (.A(\reg_module/_03077_ ),
    .B(\reg_module/gprf[169] ),
    .Y(\reg_module/_03307_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10588_  (.A(\reg_module/gprf[137] ),
    .B(net587),
    .Y(\reg_module/_03308_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10589_  (.A(\reg_module/_03307_ ),
    .B(net482),
    .C(\reg_module/_03308_ ),
    .Y(\reg_module/_03309_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10590_  (.A(\reg_module/_03081_ ),
    .B(\reg_module/gprf[233] ),
    .Y(\reg_module/_03310_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10591_  (.A(\reg_module/gprf[201] ),
    .B(net587),
    .Y(\reg_module/_03311_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10592_  (.A(\reg_module/_03310_ ),
    .B(\reg_module/_02928_ ),
    .C(\reg_module/_03311_ ),
    .Y(\reg_module/_03312_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10593_  (.A(\reg_module/_03309_ ),
    .B(\reg_module/_03312_ ),
    .Y(\reg_module/_03313_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10594_  (.A(\reg_module/_03313_ ),
    .B(\reg_module/_03086_ ),
    .Y(\reg_module/_03314_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10595_  (.A(\reg_module/_03306_ ),
    .B(\reg_module/_03314_ ),
    .C(net398),
    .Y(\reg_module/_03315_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10596_  (.A(\reg_module/_03298_ ),
    .B(\reg_module/_03315_ ),
    .Y(\reg_module/_03316_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10597_  (.A(\reg_module/_03316_ ),
    .B(net381),
    .Y(\reg_module/_03317_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_10598_  (.A(\reg_module/_03281_ ),
    .B(\reg_module/_03317_ ),
    .Y(\wRs2Data[9] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10599_  (.A(\reg_module/_03008_ ),
    .B(\reg_module/gprf[810] ),
    .Y(\reg_module/_03318_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10600_  (.A(\reg_module/gprf[778] ),
    .B(net612),
    .Y(\reg_module/_03319_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10601_  (.A(\reg_module/_03318_ ),
    .B(net494),
    .C(\reg_module/_03319_ ),
    .Y(\reg_module/_03320_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10602_  (.A(\reg_module/_03012_ ),
    .B(\reg_module/gprf[874] ),
    .Y(\reg_module/_03321_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10603_  (.A(\reg_module/gprf[842] ),
    .B(net612),
    .Y(\reg_module/_03322_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10604_  (.A(\reg_module/_03321_ ),
    .B(\reg_module/_03014_ ),
    .C(\reg_module/_03322_ ),
    .Y(\reg_module/_03323_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10605_  (.A(\reg_module/_03320_ ),
    .B(\reg_module/_03323_ ),
    .Y(\reg_module/_03324_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10606_  (.A(\reg_module/_03324_ ),
    .B(net431),
    .Y(\reg_module/_03325_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10607_  (.A(\reg_module/_02570_ ),
    .X(\reg_module/_03326_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10608_  (.A(\reg_module/_03326_ ),
    .B(\reg_module/gprf[938] ),
    .Y(\reg_module/_03327_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10609_  (.A(\reg_module/gprf[906] ),
    .B(net596),
    .Y(\reg_module/_03328_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10610_  (.A(\reg_module/_03327_ ),
    .B(net486),
    .C(\reg_module/_03328_ ),
    .Y(\reg_module/_03329_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10611_  (.A(\reg_module/_02513_ ),
    .X(\reg_module/_03330_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10612_  (.A(\reg_module/_03330_ ),
    .B(\reg_module/gprf[1002] ),
    .Y(\reg_module/_03331_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10613_  (.A(\reg_module/gprf[970] ),
    .B(net596),
    .Y(\reg_module/_03332_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10614_  (.A(\reg_module/_03331_ ),
    .B(\reg_module/_03023_ ),
    .C(\reg_module/_03332_ ),
    .Y(\reg_module/_03333_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10615_  (.A(\reg_module/_03329_ ),
    .B(\reg_module/_03333_ ),
    .Y(\reg_module/_03334_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10616_  (.A(\reg_module/_03334_ ),
    .B(\reg_module/_03179_ ),
    .Y(\reg_module/_03335_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10617_  (.A(\reg_module/_03325_ ),
    .B(\reg_module/_03335_ ),
    .C(\reg_module/_03260_ ),
    .Y(\reg_module/_03336_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10618_  (.A(\reg_module/_03182_ ),
    .B(\reg_module/gprf[682] ),
    .Y(\reg_module/_03337_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10619_  (.A(\reg_module/gprf[650] ),
    .B(net612),
    .Y(\reg_module/_03338_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10620_  (.A(\reg_module/_03337_ ),
    .B(net486),
    .C(\reg_module/_03338_ ),
    .Y(\reg_module/_03339_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10621_  (.A(\reg_module/_02535_ ),
    .X(\reg_module/_03340_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10622_  (.A(\reg_module/_03340_ ),
    .B(\reg_module/gprf[746] ),
    .Y(\reg_module/_03341_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10623_  (.A(\reg_module/gprf[714] ),
    .B(net597),
    .Y(\reg_module/_03342_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10624_  (.A(\reg_module/_03341_ ),
    .B(\reg_module/_03187_ ),
    .C(\reg_module/_03342_ ),
    .Y(\reg_module/_03343_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10625_  (.A(\reg_module/_03339_ ),
    .B(\reg_module/_03343_ ),
    .Y(\reg_module/_03344_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10626_  (.A(\reg_module/_03344_ ),
    .B(\reg_module/_03269_ ),
    .Y(\reg_module/_03345_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10627_  (.A(\reg_module/_03037_ ),
    .B(\reg_module/gprf[554] ),
    .Y(\reg_module/_03346_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10628_  (.A(\reg_module/gprf[522] ),
    .B(net615),
    .Y(\reg_module/_03347_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10629_  (.A(\reg_module/_03346_ ),
    .B(net495),
    .C(\reg_module/_03347_ ),
    .Y(\reg_module/_03348_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10630_  (.A(\reg_module/_03195_ ),
    .B(\reg_module/gprf[618] ),
    .Y(\reg_module/_03349_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10631_  (.A(\reg_module/gprf[586] ),
    .B(net615),
    .Y(\reg_module/_03350_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10632_  (.A(\reg_module/_03349_ ),
    .B(\reg_module/_03042_ ),
    .C(\reg_module/_03350_ ),
    .Y(\reg_module/_03351_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10633_  (.A(\reg_module/_03348_ ),
    .B(\reg_module/_03351_ ),
    .Y(\reg_module/_03352_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10634_  (.A(\reg_module/_03352_ ),
    .B(net431),
    .Y(\reg_module/_03353_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10635_  (.A(\reg_module/_03345_ ),
    .B(\reg_module/_03353_ ),
    .C(net399),
    .Y(\reg_module/_03354_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10636_  (.A(\reg_module/_03336_ ),
    .B(\reg_module/_03354_ ),
    .Y(\reg_module/_03355_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10637_  (.A(\reg_module/_03355_ ),
    .B(\reg_module/_03049_ ),
    .Y(\reg_module/_03356_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10638_  (.A(\reg_module/_02565_ ),
    .X(\reg_module/_03357_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10639_  (.A(\reg_module/_03357_ ),
    .B(\reg_module/gprf[298] ),
    .Y(\reg_module/_03358_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10640_  (.A(\reg_module/gprf[266] ),
    .B(net614),
    .Y(\reg_module/_03359_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10641_  (.A(\reg_module/_03358_ ),
    .B(net494),
    .C(\reg_module/_03359_ ),
    .Y(\reg_module/_03360_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10642_  (.A(\reg_module/_02897_ ),
    .X(\reg_module/_03361_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10643_  (.A(\reg_module/_03361_ ),
    .B(\reg_module/gprf[362] ),
    .Y(\reg_module/_03362_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10644_  (.A(\reg_module/_02573_ ),
    .X(\reg_module/_03363_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10645_  (.A(\reg_module/gprf[330] ),
    .B(net614),
    .Y(\reg_module/_03364_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10646_  (.A(\reg_module/_03362_ ),
    .B(\reg_module/_03363_ ),
    .C(\reg_module/_03364_ ),
    .Y(\reg_module/_03365_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10647_  (.A(\reg_module/_03360_ ),
    .B(\reg_module/_03365_ ),
    .Y(\reg_module/_03366_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10648_  (.A(\reg_module/_03366_ ),
    .B(net431),
    .Y(\reg_module/_03367_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10649_  (.A(\reg_module/_03212_ ),
    .B(\reg_module/gprf[426] ),
    .Y(\reg_module/_03368_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10650_  (.A(\reg_module/gprf[394] ),
    .B(net594),
    .Y(\reg_module/_03369_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10651_  (.A(\reg_module/_03368_ ),
    .B(net485),
    .C(\reg_module/_03369_ ),
    .Y(\reg_module/_03370_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10652_  (.A(\reg_module/_02550_ ),
    .X(\reg_module/_03371_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10653_  (.A(\reg_module/_03371_ ),
    .B(\reg_module/gprf[490] ),
    .Y(\reg_module/_03372_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10654_  (.A(\reg_module/gprf[458] ),
    .B(net593),
    .Y(\reg_module/_03373_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10655_  (.A(\reg_module/_03372_ ),
    .B(\reg_module/_03217_ ),
    .C(\reg_module/_03373_ ),
    .Y(\reg_module/_03374_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10656_  (.A(\reg_module/_03370_ ),
    .B(\reg_module/_03374_ ),
    .Y(\reg_module/_03375_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10657_  (.A(\reg_module/_03375_ ),
    .B(\reg_module/_03066_ ),
    .Y(\reg_module/_03376_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10658_  (.A(\reg_module/_03367_ ),
    .B(\reg_module/_03376_ ),
    .C(\reg_module/_03222_ ),
    .Y(\reg_module/_03377_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10659_  (.A(\reg_module/_03361_ ),
    .B(\reg_module/gprf[42] ),
    .Y(\reg_module/_03378_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10660_  (.A(\reg_module/gprf[10] ),
    .B(net615),
    .Y(\reg_module/_03379_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10661_  (.A(\reg_module/_03378_ ),
    .B(net495),
    .C(\reg_module/_03379_ ),
    .Y(\reg_module/_03380_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10662_  (.A(\reg_module/_03227_ ),
    .B(\reg_module/gprf[106] ),
    .Y(\reg_module/_03381_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10663_  (.A(\reg_module/_02604_ ),
    .X(\reg_module/_03382_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10664_  (.A(\reg_module/gprf[74] ),
    .B(net615),
    .Y(\reg_module/_03383_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10665_  (.A(\reg_module/_03381_ ),
    .B(\reg_module/_03382_ ),
    .C(\reg_module/_03383_ ),
    .Y(\reg_module/_03384_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10666_  (.A(\reg_module/_03380_ ),
    .B(\reg_module/_03384_ ),
    .Y(\reg_module/_03385_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10667_  (.A(\reg_module/_03385_ ),
    .B(net432),
    .Y(\reg_module/_03386_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10668_  (.A(\reg_module/_03077_ ),
    .B(\reg_module/gprf[170] ),
    .Y(\reg_module/_03387_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10669_  (.A(\reg_module/gprf[138] ),
    .B(net587),
    .Y(\reg_module/_03388_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10670_  (.A(\reg_module/_03387_ ),
    .B(net482),
    .C(\reg_module/_03388_ ),
    .Y(\reg_module/_03389_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10671_  (.A(\reg_module/_03081_ ),
    .B(\reg_module/gprf[234] ),
    .Y(\reg_module/_03390_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10672_  (.A(\reg_module/_02502_ ),
    .X(\reg_module/_03391_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10673_  (.A(\reg_module/gprf[202] ),
    .B(net588),
    .Y(\reg_module/_03392_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10674_  (.A(\reg_module/_03390_ ),
    .B(\reg_module/_03391_ ),
    .C(\reg_module/_03392_ ),
    .Y(\reg_module/_03393_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10675_  (.A(\reg_module/_03389_ ),
    .B(\reg_module/_03393_ ),
    .Y(\reg_module/_03394_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10676_  (.A(\reg_module/_03394_ ),
    .B(\reg_module/_03086_ ),
    .Y(\reg_module/_03395_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10677_  (.A(\reg_module/_03386_ ),
    .B(\reg_module/_03395_ ),
    .C(net402),
    .Y(\reg_module/_03396_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10678_  (.A(\reg_module/_03377_ ),
    .B(\reg_module/_03396_ ),
    .Y(\reg_module/_03397_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10679_  (.A(\reg_module/_03397_ ),
    .B(net385),
    .Y(\reg_module/_03398_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_10680_  (.A(\reg_module/_03356_ ),
    .B(\reg_module/_03398_ ),
    .Y(\wRs2Data[10] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10681_  (.A(\reg_module/_03008_ ),
    .B(\reg_module/gprf[555] ),
    .Y(\reg_module/_03399_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10682_  (.A(\reg_module/gprf[523] ),
    .B(net613),
    .Y(\reg_module/_03400_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10683_  (.A(\reg_module/_03399_ ),
    .B(net494),
    .C(\reg_module/_03400_ ),
    .Y(\reg_module/_03401_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10684_  (.A(\reg_module/_03012_ ),
    .B(\reg_module/gprf[619] ),
    .Y(\reg_module/_03402_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10685_  (.A(\reg_module/gprf[587] ),
    .B(net613),
    .Y(\reg_module/_03403_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10686_  (.A(\reg_module/_03402_ ),
    .B(\reg_module/_03014_ ),
    .C(\reg_module/_03403_ ),
    .Y(\reg_module/_03404_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10687_  (.A(\reg_module/_03401_ ),
    .B(\reg_module/_03404_ ),
    .Y(\reg_module/_03405_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10688_  (.A(\reg_module/_03405_ ),
    .B(net431),
    .Y(\reg_module/_03406_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10689_  (.A(\reg_module/_03326_ ),
    .B(\reg_module/gprf[683] ),
    .Y(\reg_module/_03407_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10690_  (.A(\reg_module/gprf[651] ),
    .B(net596),
    .Y(\reg_module/_03408_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10691_  (.A(\reg_module/_03407_ ),
    .B(net486),
    .C(\reg_module/_03408_ ),
    .Y(\reg_module/_03409_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10692_  (.A(\reg_module/_03330_ ),
    .B(\reg_module/gprf[747] ),
    .Y(\reg_module/_03410_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10693_  (.A(\reg_module/gprf[715] ),
    .B(net596),
    .Y(\reg_module/_03411_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10694_  (.A(\reg_module/_03410_ ),
    .B(\reg_module/_03023_ ),
    .C(\reg_module/_03411_ ),
    .Y(\reg_module/_03412_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10695_  (.A(\reg_module/_03409_ ),
    .B(\reg_module/_03412_ ),
    .Y(\reg_module/_03413_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10696_  (.A(\reg_module/_03413_ ),
    .B(\reg_module/_03179_ ),
    .Y(\reg_module/_03414_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10697_  (.A(\reg_module/_03406_ ),
    .B(\reg_module/_03414_ ),
    .C(net399),
    .Y(\reg_module/_03415_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10698_  (.A(\reg_module/_03182_ ),
    .B(\reg_module/gprf[811] ),
    .Y(\reg_module/_03416_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10699_  (.A(\reg_module/gprf[779] ),
    .B(net612),
    .Y(\reg_module/_03417_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10700_  (.A(\reg_module/_03416_ ),
    .B(net494),
    .C(\reg_module/_03417_ ),
    .Y(\reg_module/_03418_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10701_  (.A(\reg_module/_03340_ ),
    .B(\reg_module/gprf[875] ),
    .Y(\reg_module/_03419_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10702_  (.A(\reg_module/gprf[843] ),
    .B(net613),
    .Y(\reg_module/_03420_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10703_  (.A(\reg_module/_03419_ ),
    .B(\reg_module/_03187_ ),
    .C(\reg_module/_03420_ ),
    .Y(\reg_module/_03421_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10704_  (.A(\reg_module/_03418_ ),
    .B(\reg_module/_03421_ ),
    .Y(\reg_module/_03422_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10705_  (.A(\reg_module/_03422_ ),
    .B(net430),
    .Y(\reg_module/_03423_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10706_  (.A(\reg_module/_03037_ ),
    .B(\reg_module/gprf[939] ),
    .Y(\reg_module/_03424_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10707_  (.A(\reg_module/gprf[907] ),
    .B(net596),
    .Y(\reg_module/_03425_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10708_  (.A(\reg_module/_03424_ ),
    .B(net486),
    .C(\reg_module/_03425_ ),
    .Y(\reg_module/_03426_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10709_  (.A(\reg_module/_03195_ ),
    .B(\reg_module/gprf[1003] ),
    .Y(\reg_module/_03427_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10710_  (.A(\reg_module/gprf[971] ),
    .B(net597),
    .Y(\reg_module/_03428_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10711_  (.A(\reg_module/_03427_ ),
    .B(\reg_module/_03042_ ),
    .C(\reg_module/_03428_ ),
    .Y(\reg_module/_03429_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10712_  (.A(\reg_module/_03426_ ),
    .B(\reg_module/_03429_ ),
    .Y(\reg_module/_03430_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10713_  (.A(\reg_module/_03430_ ),
    .B(\reg_module/_02736_ ),
    .Y(\reg_module/_03431_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10714_  (.A(\reg_module/_03423_ ),
    .B(\reg_module/_03431_ ),
    .C(\reg_module/_02738_ ),
    .Y(\reg_module/_03432_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10715_  (.A(\reg_module/_03415_ ),
    .B(\reg_module/_03432_ ),
    .Y(\reg_module/_03433_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10716_  (.A(\reg_module/_03433_ ),
    .B(\reg_module/_03049_ ),
    .Y(\reg_module/_03434_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10717_  (.A(\reg_module/_03357_ ),
    .B(\reg_module/gprf[299] ),
    .Y(\reg_module/_03435_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10718_  (.A(\reg_module/gprf[267] ),
    .B(net614),
    .Y(\reg_module/_03436_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10719_  (.A(\reg_module/_03435_ ),
    .B(net497),
    .C(\reg_module/_03436_ ),
    .Y(\reg_module/_03437_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10720_  (.A(\reg_module/_03361_ ),
    .B(\reg_module/gprf[363] ),
    .Y(\reg_module/_03438_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10721_  (.A(\reg_module/gprf[331] ),
    .B(net614),
    .Y(\reg_module/_03439_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10722_  (.A(\reg_module/_03438_ ),
    .B(\reg_module/_03363_ ),
    .C(\reg_module/_03439_ ),
    .Y(\reg_module/_03440_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10723_  (.A(\reg_module/_03437_ ),
    .B(\reg_module/_03440_ ),
    .Y(\reg_module/_03441_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10724_  (.A(\reg_module/_03441_ ),
    .B(net431),
    .Y(\reg_module/_03442_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10725_  (.A(\reg_module/_03212_ ),
    .B(\reg_module/gprf[427] ),
    .Y(\reg_module/_03443_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10726_  (.A(\reg_module/gprf[395] ),
    .B(net594),
    .Y(\reg_module/_03444_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10727_  (.A(\reg_module/_03443_ ),
    .B(net485),
    .C(\reg_module/_03444_ ),
    .Y(\reg_module/_03445_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10728_  (.A(\reg_module/_03371_ ),
    .B(\reg_module/gprf[491] ),
    .Y(\reg_module/_03446_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10729_  (.A(\reg_module/gprf[459] ),
    .B(net593),
    .Y(\reg_module/_03447_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10730_  (.A(\reg_module/_03446_ ),
    .B(\reg_module/_03217_ ),
    .C(\reg_module/_03447_ ),
    .Y(\reg_module/_03448_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10731_  (.A(\reg_module/_03445_ ),
    .B(\reg_module/_03448_ ),
    .Y(\reg_module/_03449_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10732_  (.A(\reg_module/_03449_ ),
    .B(\reg_module/_03066_ ),
    .Y(\reg_module/_03450_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10733_  (.A(\reg_module/_03442_ ),
    .B(\reg_module/_03450_ ),
    .C(\reg_module/_03222_ ),
    .Y(\reg_module/_03451_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10734_  (.A(\reg_module/_03361_ ),
    .B(\reg_module/gprf[43] ),
    .Y(\reg_module/_03452_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10735_  (.A(\reg_module/gprf[11] ),
    .B(net616),
    .Y(\reg_module/_03453_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10736_  (.A(\reg_module/_03452_ ),
    .B(net495),
    .C(\reg_module/_03453_ ),
    .Y(\reg_module/_03454_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10737_  (.A(\reg_module/_03227_ ),
    .B(\reg_module/gprf[107] ),
    .Y(\reg_module/_03455_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10738_  (.A(\reg_module/gprf[75] ),
    .B(net616),
    .Y(\reg_module/_03456_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10739_  (.A(\reg_module/_03455_ ),
    .B(\reg_module/_03382_ ),
    .C(\reg_module/_03456_ ),
    .Y(\reg_module/_03457_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10740_  (.A(\reg_module/_03454_ ),
    .B(\reg_module/_03457_ ),
    .Y(\reg_module/_03458_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10741_  (.A(\reg_module/_03458_ ),
    .B(net432),
    .Y(\reg_module/_03459_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10742_  (.A(\reg_module/_03077_ ),
    .B(\reg_module/gprf[171] ),
    .Y(\reg_module/_03460_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10743_  (.A(\reg_module/gprf[139] ),
    .B(net587),
    .Y(\reg_module/_03461_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10744_  (.A(\reg_module/_03460_ ),
    .B(net482),
    .C(\reg_module/_03461_ ),
    .Y(\reg_module/_03462_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10745_  (.A(\reg_module/_03081_ ),
    .B(\reg_module/gprf[235] ),
    .Y(\reg_module/_03463_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10746_  (.A(\reg_module/gprf[203] ),
    .B(net588),
    .Y(\reg_module/_03464_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10747_  (.A(\reg_module/_03463_ ),
    .B(\reg_module/_03391_ ),
    .C(\reg_module/_03464_ ),
    .Y(\reg_module/_03465_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10748_  (.A(\reg_module/_03462_ ),
    .B(\reg_module/_03465_ ),
    .Y(\reg_module/_03466_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10749_  (.A(\reg_module/_03466_ ),
    .B(\reg_module/_03086_ ),
    .Y(\reg_module/_03467_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10750_  (.A(\reg_module/_03459_ ),
    .B(\reg_module/_03467_ ),
    .C(net402),
    .Y(\reg_module/_03468_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10751_  (.A(\reg_module/_03451_ ),
    .B(\reg_module/_03468_ ),
    .Y(\reg_module/_03469_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10752_  (.A(\reg_module/_03469_ ),
    .B(net385),
    .Y(\reg_module/_03470_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_10753_  (.A(\reg_module/_03434_ ),
    .B(\reg_module/_03470_ ),
    .Y(\wRs2Data[11] ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10754_  (.A(\reg_module/_02492_ ),
    .X(\reg_module/_03471_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10755_  (.A(\reg_module/_03471_ ),
    .B(\reg_module/gprf[812] ),
    .Y(\reg_module/_03472_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10756_  (.A(\reg_module/gprf[780] ),
    .B(net622),
    .Y(\reg_module/_03473_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10757_  (.A(\reg_module/_03472_ ),
    .B(net498),
    .C(\reg_module/_03473_ ),
    .Y(\reg_module/_03474_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10758_  (.A(\reg_module/_02498_ ),
    .X(\reg_module/_03475_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10759_  (.A(\reg_module/_03475_ ),
    .B(\reg_module/gprf[876] ),
    .Y(\reg_module/_03476_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10760_  (.A(\reg_module/_02573_ ),
    .X(\reg_module/_03477_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10761_  (.A(\reg_module/gprf[844] ),
    .B(net622),
    .Y(\reg_module/_03478_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10762_  (.A(\reg_module/_03476_ ),
    .B(\reg_module/_03477_ ),
    .C(\reg_module/_03478_ ),
    .Y(\reg_module/_03479_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10763_  (.A(\reg_module/_03474_ ),
    .B(\reg_module/_03479_ ),
    .Y(\reg_module/_03480_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10764_  (.A(\reg_module/_03480_ ),
    .B(net433),
    .Y(\reg_module/_03481_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10765_  (.A(\reg_module/_03326_ ),
    .B(\reg_module/gprf[940] ),
    .Y(\reg_module/_03482_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10766_  (.A(\reg_module/gprf[908] ),
    .B(net598),
    .Y(\reg_module/_03483_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10767_  (.A(\reg_module/_03482_ ),
    .B(net487),
    .C(\reg_module/_03483_ ),
    .Y(\reg_module/_03484_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10768_  (.A(\reg_module/_03330_ ),
    .B(\reg_module/gprf[1004] ),
    .Y(\reg_module/_03485_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10769_  (.A(\reg_module/_02516_ ),
    .X(\reg_module/_03486_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10770_  (.A(\reg_module/gprf[972] ),
    .B(net598),
    .Y(\reg_module/_03487_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10771_  (.A(\reg_module/_03485_ ),
    .B(\reg_module/_03486_ ),
    .C(\reg_module/_03487_ ),
    .Y(\reg_module/_03488_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10772_  (.A(\reg_module/_03484_ ),
    .B(\reg_module/_03488_ ),
    .Y(\reg_module/_03489_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10773_  (.A(\reg_module/_03489_ ),
    .B(\reg_module/_03179_ ),
    .Y(\reg_module/_03490_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10774_  (.A(\reg_module/_03481_ ),
    .B(\reg_module/_03490_ ),
    .C(\reg_module/_03260_ ),
    .Y(\reg_module/_03491_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10775_  (.A(\reg_module/_03182_ ),
    .B(\reg_module/gprf[684] ),
    .Y(\reg_module/_03492_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10776_  (.A(\reg_module/gprf[652] ),
    .B(net600),
    .Y(\reg_module/_03493_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10777_  (.A(\reg_module/_03492_ ),
    .B(net486),
    .C(\reg_module/_03493_ ),
    .Y(\reg_module/_03494_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10778_  (.A(\reg_module/_03340_ ),
    .B(\reg_module/gprf[748] ),
    .Y(\reg_module/_03495_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10779_  (.A(\reg_module/gprf[716] ),
    .B(net599),
    .Y(\reg_module/_03496_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10780_  (.A(\reg_module/_03495_ ),
    .B(\reg_module/_03187_ ),
    .C(\reg_module/_03496_ ),
    .Y(\reg_module/_03497_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10781_  (.A(\reg_module/_03494_ ),
    .B(\reg_module/_03497_ ),
    .Y(\reg_module/_03498_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10782_  (.A(\reg_module/_03498_ ),
    .B(\reg_module/_03269_ ),
    .Y(\reg_module/_03499_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10783_  (.A(\reg_module/_02545_ ),
    .X(\reg_module/_03500_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10784_  (.A(\reg_module/_03500_ ),
    .B(\reg_module/gprf[556] ),
    .Y(\reg_module/_03501_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10785_  (.A(\reg_module/gprf[524] ),
    .B(net626),
    .Y(\reg_module/_03502_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10786_  (.A(\reg_module/_03501_ ),
    .B(net500),
    .C(\reg_module/_03502_ ),
    .Y(\reg_module/_03503_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10787_  (.A(\reg_module/_03195_ ),
    .B(\reg_module/gprf[620] ),
    .Y(\reg_module/_03504_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10788_  (.A(\reg_module/_02553_ ),
    .X(\reg_module/_03505_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10789_  (.A(\reg_module/gprf[588] ),
    .B(net619),
    .Y(\reg_module/_03506_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10790_  (.A(\reg_module/_03504_ ),
    .B(\reg_module/_03505_ ),
    .C(\reg_module/_03506_ ),
    .Y(\reg_module/_03507_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10791_  (.A(\reg_module/_03503_ ),
    .B(\reg_module/_03507_ ),
    .Y(\reg_module/_03508_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10792_  (.A(\reg_module/_03508_ ),
    .B(net433),
    .Y(\reg_module/_03509_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10793_  (.A(\reg_module/_03499_ ),
    .B(\reg_module/_03509_ ),
    .C(net400),
    .Y(\reg_module/_03510_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10794_  (.A(\reg_module/_03491_ ),
    .B(\reg_module/_03510_ ),
    .Y(\reg_module/_03511_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10795_  (.A(\reg_module/_02562_ ),
    .X(\reg_module/_03512_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10796_  (.A(\reg_module/_03511_ ),
    .B(\reg_module/_03512_ ),
    .Y(\reg_module/_03513_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10797_  (.A(\reg_module/_03357_ ),
    .B(\reg_module/gprf[300] ),
    .Y(\reg_module/_03514_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10798_  (.A(\reg_module/gprf[268] ),
    .B(net624),
    .Y(\reg_module/_03515_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10799_  (.A(\reg_module/_03514_ ),
    .B(net498),
    .C(\reg_module/_03515_ ),
    .Y(\reg_module/_03516_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10800_  (.A(\reg_module/_03361_ ),
    .B(\reg_module/gprf[364] ),
    .Y(\reg_module/_03517_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10801_  (.A(\reg_module/gprf[332] ),
    .B(net623),
    .Y(\reg_module/_03518_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10802_  (.A(\reg_module/_03517_ ),
    .B(\reg_module/_03363_ ),
    .C(\reg_module/_03518_ ),
    .Y(\reg_module/_03519_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10803_  (.A(\reg_module/_03516_ ),
    .B(\reg_module/_03519_ ),
    .Y(\reg_module/_03520_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10804_  (.A(\reg_module/_03520_ ),
    .B(net433),
    .Y(\reg_module/_03521_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10805_  (.A(\reg_module/_03212_ ),
    .B(\reg_module/gprf[428] ),
    .Y(\reg_module/_03522_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10806_  (.A(\reg_module/gprf[396] ),
    .B(net602),
    .Y(\reg_module/_03523_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10807_  (.A(\reg_module/_03522_ ),
    .B(net490),
    .C(\reg_module/_03523_ ),
    .Y(\reg_module/_03524_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10808_  (.A(\reg_module/_03371_ ),
    .B(\reg_module/gprf[492] ),
    .Y(\reg_module/_03525_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10809_  (.A(\reg_module/gprf[460] ),
    .B(net603),
    .Y(\reg_module/_03526_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10810_  (.A(\reg_module/_03525_ ),
    .B(\reg_module/_03217_ ),
    .C(\reg_module/_03526_ ),
    .Y(\reg_module/_03527_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10811_  (.A(\reg_module/_03524_ ),
    .B(\reg_module/_03527_ ),
    .Y(\reg_module/_03528_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_10812_  (.A(\reg_module/_02735_ ),
    .X(\reg_module/_03529_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10813_  (.A(\reg_module/_03528_ ),
    .B(\reg_module/_03529_ ),
    .Y(\reg_module/_03530_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10814_  (.A(\reg_module/_03521_ ),
    .B(\reg_module/_03530_ ),
    .C(\reg_module/_03222_ ),
    .Y(\reg_module/_03531_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10815_  (.A(\reg_module/_03361_ ),
    .B(\reg_module/gprf[44] ),
    .Y(\reg_module/_03532_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10816_  (.A(\reg_module/gprf[12] ),
    .B(net627),
    .Y(\reg_module/_03533_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10817_  (.A(\reg_module/_03532_ ),
    .B(net500),
    .C(\reg_module/_03533_ ),
    .Y(\reg_module/_03534_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10818_  (.A(\reg_module/_03227_ ),
    .B(\reg_module/gprf[108] ),
    .Y(\reg_module/_03535_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10819_  (.A(\reg_module/gprf[76] ),
    .B(net627),
    .Y(\reg_module/_03536_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10820_  (.A(\reg_module/_03535_ ),
    .B(\reg_module/_03382_ ),
    .C(\reg_module/_03536_ ),
    .Y(\reg_module/_03537_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10821_  (.A(\reg_module/_03534_ ),
    .B(\reg_module/_03537_ ),
    .Y(\reg_module/_03538_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10822_  (.A(\reg_module/_03538_ ),
    .B(net434),
    .Y(\reg_module/_03539_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10823_  (.A(\reg_module/_02584_ ),
    .X(\reg_module/_03540_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10824_  (.A(\reg_module/_03540_ ),
    .B(\reg_module/gprf[172] ),
    .Y(\reg_module/_03541_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10825_  (.A(\reg_module/gprf[140] ),
    .B(net617),
    .Y(\reg_module/_03542_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10826_  (.A(\reg_module/_03541_ ),
    .B(net495),
    .C(\reg_module/_03542_ ),
    .Y(\reg_module/_03543_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10827_  (.A(\reg_module/_02491_ ),
    .X(\reg_module/_03544_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10828_  (.A(\reg_module/_03544_ ),
    .B(\reg_module/gprf[236] ),
    .Y(\reg_module/_03545_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10829_  (.A(\reg_module/gprf[204] ),
    .B(net617),
    .Y(\reg_module/_03546_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10830_  (.A(\reg_module/_03545_ ),
    .B(\reg_module/_03391_ ),
    .C(\reg_module/_03546_ ),
    .Y(\reg_module/_03547_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10831_  (.A(\reg_module/_03543_ ),
    .B(\reg_module/_03547_ ),
    .Y(\reg_module/_03548_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_10832_  (.A(\reg_module/_02522_ ),
    .X(\reg_module/_03549_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10833_  (.A(\reg_module/_03548_ ),
    .B(\reg_module/_03549_ ),
    .Y(\reg_module/_03550_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10834_  (.A(\reg_module/_03539_ ),
    .B(\reg_module/_03550_ ),
    .C(net401),
    .Y(\reg_module/_03551_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10835_  (.A(\reg_module/_03531_ ),
    .B(\reg_module/_03551_ ),
    .Y(\reg_module/_03552_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10836_  (.A(\reg_module/_03552_ ),
    .B(net384),
    .Y(\reg_module/_03553_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_10837_  (.A(\reg_module/_03513_ ),
    .B(\reg_module/_03553_ ),
    .Y(\wRs2Data[12] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10838_  (.A(\reg_module/_03471_ ),
    .B(\reg_module/gprf[813] ),
    .Y(\reg_module/_03554_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10839_  (.A(\reg_module/gprf[781] ),
    .B(net622),
    .Y(\reg_module/_03555_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10840_  (.A(\reg_module/_03554_ ),
    .B(net498),
    .C(\reg_module/_03555_ ),
    .Y(\reg_module/_03556_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10841_  (.A(\reg_module/_03475_ ),
    .B(\reg_module/gprf[877] ),
    .Y(\reg_module/_03557_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10842_  (.A(\reg_module/gprf[845] ),
    .B(net614),
    .Y(\reg_module/_03558_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10843_  (.A(\reg_module/_03557_ ),
    .B(\reg_module/_03477_ ),
    .C(\reg_module/_03558_ ),
    .Y(\reg_module/_03559_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10844_  (.A(\reg_module/_03556_ ),
    .B(\reg_module/_03559_ ),
    .Y(\reg_module/_03560_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10845_  (.A(\reg_module/_03560_ ),
    .B(net433),
    .Y(\reg_module/_03561_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10846_  (.A(\reg_module/_03326_ ),
    .B(\reg_module/gprf[941] ),
    .Y(\reg_module/_03562_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10847_  (.A(\reg_module/gprf[909] ),
    .B(net598),
    .Y(\reg_module/_03563_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10848_  (.A(\reg_module/_03562_ ),
    .B(net487),
    .C(\reg_module/_03563_ ),
    .Y(\reg_module/_03564_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10849_  (.A(\reg_module/_03330_ ),
    .B(\reg_module/gprf[1005] ),
    .Y(\reg_module/_03565_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10850_  (.A(\reg_module/gprf[973] ),
    .B(net598),
    .Y(\reg_module/_03566_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10851_  (.A(\reg_module/_03565_ ),
    .B(\reg_module/_03486_ ),
    .C(\reg_module/_03566_ ),
    .Y(\reg_module/_03567_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10852_  (.A(\reg_module/_03564_ ),
    .B(\reg_module/_03567_ ),
    .Y(\reg_module/_03568_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10853_  (.A(\reg_module/_03568_ ),
    .B(\reg_module/_03179_ ),
    .Y(\reg_module/_03569_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10854_  (.A(\reg_module/_03561_ ),
    .B(\reg_module/_03569_ ),
    .C(\reg_module/_03260_ ),
    .Y(\reg_module/_03570_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10855_  (.A(\reg_module/_03182_ ),
    .B(\reg_module/gprf[685] ),
    .Y(\reg_module/_03571_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10856_  (.A(\reg_module/gprf[653] ),
    .B(net621),
    .Y(\reg_module/_03572_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10857_  (.A(\reg_module/_03571_ ),
    .B(net494),
    .C(\reg_module/_03572_ ),
    .Y(\reg_module/_03573_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10858_  (.A(\reg_module/_03340_ ),
    .B(\reg_module/gprf[749] ),
    .Y(\reg_module/_03574_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10859_  (.A(\reg_module/gprf[717] ),
    .B(net599),
    .Y(\reg_module/_03575_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10860_  (.A(\reg_module/_03574_ ),
    .B(\reg_module/_03187_ ),
    .C(\reg_module/_03575_ ),
    .Y(\reg_module/_03576_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10861_  (.A(\reg_module/_03573_ ),
    .B(\reg_module/_03576_ ),
    .Y(\reg_module/_03577_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10862_  (.A(\reg_module/_03577_ ),
    .B(\reg_module/_03269_ ),
    .Y(\reg_module/_03578_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10863_  (.A(\reg_module/_03500_ ),
    .B(\reg_module/gprf[557] ),
    .Y(\reg_module/_03579_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10864_  (.A(\reg_module/gprf[525] ),
    .B(net626),
    .Y(\reg_module/_03580_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10865_  (.A(\reg_module/_03579_ ),
    .B(net500),
    .C(\reg_module/_03580_ ),
    .Y(\reg_module/_03581_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10866_  (.A(\reg_module/_03195_ ),
    .B(\reg_module/gprf[621] ),
    .Y(\reg_module/_03582_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10867_  (.A(\reg_module/gprf[589] ),
    .B(net619),
    .Y(\reg_module/_03583_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10868_  (.A(\reg_module/_03582_ ),
    .B(\reg_module/_03505_ ),
    .C(\reg_module/_03583_ ),
    .Y(\reg_module/_03584_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10869_  (.A(\reg_module/_03581_ ),
    .B(\reg_module/_03584_ ),
    .Y(\reg_module/_03585_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10870_  (.A(\reg_module/_03585_ ),
    .B(net434),
    .Y(\reg_module/_03586_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10871_  (.A(\reg_module/_03578_ ),
    .B(\reg_module/_03586_ ),
    .C(net401),
    .Y(\reg_module/_03587_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10872_  (.A(\reg_module/_03570_ ),
    .B(\reg_module/_03587_ ),
    .Y(\reg_module/_03588_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10873_  (.A(\reg_module/_03588_ ),
    .B(\reg_module/_03512_ ),
    .Y(\reg_module/_03589_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10874_  (.A(\reg_module/_03357_ ),
    .B(\reg_module/gprf[301] ),
    .Y(\reg_module/_03590_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10875_  (.A(\reg_module/gprf[269] ),
    .B(net624),
    .Y(\reg_module/_03591_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10876_  (.A(\reg_module/_03590_ ),
    .B(net498),
    .C(\reg_module/_03591_ ),
    .Y(\reg_module/_03592_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10877_  (.A(\reg_module/_02897_ ),
    .X(\reg_module/_03593_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10878_  (.A(\reg_module/_03593_ ),
    .B(\reg_module/gprf[365] ),
    .Y(\reg_module/_03594_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10879_  (.A(\reg_module/gprf[333] ),
    .B(net624),
    .Y(\reg_module/_03595_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10880_  (.A(\reg_module/_03594_ ),
    .B(\reg_module/_03363_ ),
    .C(\reg_module/_03595_ ),
    .Y(\reg_module/_03596_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10881_  (.A(\reg_module/_03592_ ),
    .B(\reg_module/_03596_ ),
    .Y(\reg_module/_03597_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10882_  (.A(\reg_module/_03597_ ),
    .B(net436),
    .Y(\reg_module/_03598_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10883_  (.A(\reg_module/_03212_ ),
    .B(\reg_module/gprf[429] ),
    .Y(\reg_module/_03599_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10884_  (.A(\reg_module/gprf[397] ),
    .B(net604),
    .Y(\reg_module/_03600_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10885_  (.A(\reg_module/_03599_ ),
    .B(net489),
    .C(\reg_module/_03600_ ),
    .Y(\reg_module/_03601_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10886_  (.A(\reg_module/_03371_ ),
    .B(\reg_module/gprf[493] ),
    .Y(\reg_module/_03602_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10887_  (.A(\reg_module/gprf[461] ),
    .B(net603),
    .Y(\reg_module/_03603_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10888_  (.A(\reg_module/_03602_ ),
    .B(\reg_module/_03217_ ),
    .C(\reg_module/_03603_ ),
    .Y(\reg_module/_03604_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10889_  (.A(\reg_module/_03601_ ),
    .B(\reg_module/_03604_ ),
    .Y(\reg_module/_03605_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10890_  (.A(\reg_module/_03605_ ),
    .B(\reg_module/_03529_ ),
    .Y(\reg_module/_03606_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10891_  (.A(\reg_module/_03598_ ),
    .B(\reg_module/_03606_ ),
    .C(\reg_module/_03222_ ),
    .Y(\reg_module/_03607_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10892_  (.A(\reg_module/_03593_ ),
    .B(\reg_module/gprf[45] ),
    .Y(\reg_module/_03608_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10893_  (.A(\reg_module/gprf[13] ),
    .B(net628),
    .Y(\reg_module/_03609_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10894_  (.A(\reg_module/_03608_ ),
    .B(net501),
    .C(\reg_module/_03609_ ),
    .Y(\reg_module/_03610_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10895_  (.A(\reg_module/_03227_ ),
    .B(\reg_module/gprf[109] ),
    .Y(\reg_module/_03611_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10896_  (.A(\reg_module/gprf[77] ),
    .B(net627),
    .Y(\reg_module/_03612_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10897_  (.A(\reg_module/_03611_ ),
    .B(\reg_module/_03382_ ),
    .C(\reg_module/_03612_ ),
    .Y(\reg_module/_03613_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10898_  (.A(\reg_module/_03610_ ),
    .B(\reg_module/_03613_ ),
    .Y(\reg_module/_03614_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10899_  (.A(\reg_module/_03614_ ),
    .B(net435),
    .Y(\reg_module/_03615_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10900_  (.A(\reg_module/_03540_ ),
    .B(\reg_module/gprf[173] ),
    .Y(\reg_module/_03616_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10901_  (.A(\reg_module/gprf[141] ),
    .B(net627),
    .Y(\reg_module/_03617_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10902_  (.A(\reg_module/_03616_ ),
    .B(net500),
    .C(\reg_module/_03617_ ),
    .Y(\reg_module/_03618_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10903_  (.A(\reg_module/_03544_ ),
    .B(\reg_module/gprf[237] ),
    .Y(\reg_module/_03619_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10904_  (.A(\reg_module/gprf[205] ),
    .B(net618),
    .Y(\reg_module/_03620_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10905_  (.A(\reg_module/_03619_ ),
    .B(\reg_module/_03391_ ),
    .C(\reg_module/_03620_ ),
    .Y(\reg_module/_03621_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10906_  (.A(\reg_module/_03618_ ),
    .B(\reg_module/_03621_ ),
    .Y(\reg_module/_03622_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10907_  (.A(\reg_module/_03622_ ),
    .B(\reg_module/_03549_ ),
    .Y(\reg_module/_03623_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10908_  (.A(\reg_module/_03615_ ),
    .B(\reg_module/_03623_ ),
    .C(net402),
    .Y(\reg_module/_03624_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10909_  (.A(\reg_module/_03607_ ),
    .B(\reg_module/_03624_ ),
    .Y(\reg_module/_03625_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10910_  (.A(\reg_module/_03625_ ),
    .B(net384),
    .Y(\reg_module/_03626_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_10911_  (.A(\reg_module/_03589_ ),
    .B(\reg_module/_03626_ ),
    .Y(\wRs2Data[13] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10912_  (.A(\reg_module/_03471_ ),
    .B(\reg_module/gprf[558] ),
    .Y(\reg_module/_03627_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10913_  (.A(\reg_module/gprf[526] ),
    .B(net623),
    .Y(\reg_module/_03628_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10914_  (.A(\reg_module/_03627_ ),
    .B(net498),
    .C(\reg_module/_03628_ ),
    .Y(\reg_module/_03629_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10915_  (.A(\reg_module/_03475_ ),
    .B(\reg_module/gprf[622] ),
    .Y(\reg_module/_03630_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10916_  (.A(\reg_module/gprf[590] ),
    .B(net623),
    .Y(\reg_module/_03631_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10917_  (.A(\reg_module/_03630_ ),
    .B(\reg_module/_03477_ ),
    .C(\reg_module/_03631_ ),
    .Y(\reg_module/_03632_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10918_  (.A(\reg_module/_03629_ ),
    .B(\reg_module/_03632_ ),
    .Y(\reg_module/_03633_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10919_  (.A(\reg_module/_03633_ ),
    .B(net433),
    .Y(\reg_module/_03634_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10920_  (.A(\reg_module/_03326_ ),
    .B(\reg_module/gprf[686] ),
    .Y(\reg_module/_03635_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10921_  (.A(\reg_module/gprf[654] ),
    .B(net598),
    .Y(\reg_module/_03636_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10922_  (.A(\reg_module/_03635_ ),
    .B(net487),
    .C(\reg_module/_03636_ ),
    .Y(\reg_module/_03637_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10923_  (.A(\reg_module/_03330_ ),
    .B(\reg_module/gprf[750] ),
    .Y(\reg_module/_03638_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10924_  (.A(\reg_module/gprf[718] ),
    .B(net598),
    .Y(\reg_module/_03639_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10925_  (.A(\reg_module/_03638_ ),
    .B(\reg_module/_03486_ ),
    .C(\reg_module/_03639_ ),
    .Y(\reg_module/_03640_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10926_  (.A(\reg_module/_03637_ ),
    .B(\reg_module/_03640_ ),
    .Y(\reg_module/_03641_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10927_  (.A(\reg_module/_02592_ ),
    .X(\reg_module/_03642_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10928_  (.A(\reg_module/_03641_ ),
    .B(\reg_module/_03642_ ),
    .Y(\reg_module/_03643_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10929_  (.A(\reg_module/_03634_ ),
    .B(\reg_module/_03643_ ),
    .C(net399),
    .Y(\reg_module/_03644_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10930_  (.A(\reg_module/_02530_ ),
    .X(\reg_module/_03645_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10931_  (.A(\reg_module/_03645_ ),
    .B(\reg_module/gprf[814] ),
    .Y(\reg_module/_03646_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10932_  (.A(\reg_module/gprf[782] ),
    .B(net609),
    .Y(\reg_module/_03647_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10933_  (.A(\reg_module/_03646_ ),
    .B(net491),
    .C(\reg_module/_03647_ ),
    .Y(\reg_module/_03648_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10934_  (.A(\reg_module/_03340_ ),
    .B(\reg_module/gprf[878] ),
    .Y(\reg_module/_03649_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10935_  (.A(\reg_module/_02538_ ),
    .X(\reg_module/_03650_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10936_  (.A(\reg_module/gprf[846] ),
    .B(net608),
    .Y(\reg_module/_03651_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10937_  (.A(\reg_module/_03649_ ),
    .B(\reg_module/_03650_ ),
    .C(\reg_module/_03651_ ),
    .Y(\reg_module/_03652_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10938_  (.A(\reg_module/_03648_ ),
    .B(\reg_module/_03652_ ),
    .Y(\reg_module/_03653_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10939_  (.A(\reg_module/_03653_ ),
    .B(net428),
    .Y(\reg_module/_03654_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10940_  (.A(\reg_module/_03500_ ),
    .B(\reg_module/gprf[942] ),
    .Y(\reg_module/_03655_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10941_  (.A(\reg_module/gprf[910] ),
    .B(net608),
    .Y(\reg_module/_03656_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10942_  (.A(\reg_module/_03655_ ),
    .B(net491),
    .C(\reg_module/_03656_ ),
    .Y(\reg_module/_03657_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_10943_  (.A(\reg_module/_02614_ ),
    .X(\reg_module/_03658_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10944_  (.A(\reg_module/_03658_ ),
    .B(\reg_module/gprf[1006] ),
    .Y(\reg_module/_03659_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10945_  (.A(\reg_module/gprf[974] ),
    .B(net608),
    .Y(\reg_module/_03660_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10946_  (.A(\reg_module/_03659_ ),
    .B(\reg_module/_03505_ ),
    .C(\reg_module/_03660_ ),
    .Y(\reg_module/_03661_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10947_  (.A(\reg_module/_03657_ ),
    .B(\reg_module/_03661_ ),
    .Y(\reg_module/_03662_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_10948_  (.A(\reg_module/_02735_ ),
    .X(\reg_module/_03663_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10949_  (.A(\reg_module/_03662_ ),
    .B(\reg_module/_03663_ ),
    .Y(\reg_module/_03664_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10950_  (.A(\reg_module/_03654_ ),
    .B(\reg_module/_03664_ ),
    .C(\reg_module/_02738_ ),
    .Y(\reg_module/_03665_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10951_  (.A(\reg_module/_03644_ ),
    .B(\reg_module/_03665_ ),
    .Y(\reg_module/_03666_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10952_  (.A(\reg_module/_03666_ ),
    .B(\reg_module/_03512_ ),
    .Y(\reg_module/_03667_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10953_  (.A(\reg_module/_03357_ ),
    .B(\reg_module/gprf[302] ),
    .Y(\reg_module/_03668_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10954_  (.A(\reg_module/gprf[270] ),
    .B(net624),
    .Y(\reg_module/_03669_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10955_  (.A(\reg_module/_03668_ ),
    .B(net499),
    .C(\reg_module/_03669_ ),
    .Y(\reg_module/_03670_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10956_  (.A(\reg_module/_03593_ ),
    .B(\reg_module/gprf[366] ),
    .Y(\reg_module/_03671_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10957_  (.A(\reg_module/gprf[334] ),
    .B(net625),
    .Y(\reg_module/_03672_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10958_  (.A(\reg_module/_03671_ ),
    .B(\reg_module/_03363_ ),
    .C(\reg_module/_03672_ ),
    .Y(\reg_module/_03673_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10959_  (.A(\reg_module/_03670_ ),
    .B(\reg_module/_03673_ ),
    .Y(\reg_module/_03674_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10960_  (.A(\reg_module/_03674_ ),
    .B(net428),
    .Y(\reg_module/_03675_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10961_  (.A(\reg_module/_02579_ ),
    .X(\reg_module/_03676_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10962_  (.A(\reg_module/_03676_ ),
    .B(\reg_module/gprf[430] ),
    .Y(\reg_module/_03677_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10963_  (.A(\reg_module/gprf[398] ),
    .B(net604),
    .Y(\reg_module/_03678_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10964_  (.A(\reg_module/_03677_ ),
    .B(net490),
    .C(\reg_module/_03678_ ),
    .Y(\reg_module/_03679_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10965_  (.A(\reg_module/_03371_ ),
    .B(\reg_module/gprf[494] ),
    .Y(\reg_module/_03680_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10966_  (.A(\reg_module/_02587_ ),
    .X(\reg_module/_03681_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10967_  (.A(\reg_module/gprf[462] ),
    .B(net602),
    .Y(\reg_module/_03682_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10968_  (.A(\reg_module/_03680_ ),
    .B(\reg_module/_03681_ ),
    .C(\reg_module/_03682_ ),
    .Y(\reg_module/_03683_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10969_  (.A(\reg_module/_03679_ ),
    .B(\reg_module/_03683_ ),
    .Y(\reg_module/_03684_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10970_  (.A(\reg_module/_03684_ ),
    .B(\reg_module/_03529_ ),
    .Y(\reg_module/_03685_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_10971_  (.A(\reg_module/_02595_ ),
    .X(\reg_module/_03686_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10972_  (.A(\reg_module/_03675_ ),
    .B(\reg_module/_03685_ ),
    .C(\reg_module/_03686_ ),
    .Y(\reg_module/_03687_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10973_  (.A(\reg_module/_03593_ ),
    .B(\reg_module/gprf[46] ),
    .Y(\reg_module/_03688_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10974_  (.A(\reg_module/gprf[14] ),
    .B(net629),
    .Y(\reg_module/_03689_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10975_  (.A(\reg_module/_03688_ ),
    .B(net501),
    .C(\reg_module/_03689_ ),
    .Y(\reg_module/_03690_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_10976_  (.A(\reg_module/_02601_ ),
    .X(\reg_module/_03691_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10977_  (.A(\reg_module/_03691_ ),
    .B(\reg_module/gprf[110] ),
    .Y(\reg_module/_03692_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10978_  (.A(\reg_module/gprf[78] ),
    .B(net627),
    .Y(\reg_module/_03693_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10979_  (.A(\reg_module/_03692_ ),
    .B(\reg_module/_03382_ ),
    .C(\reg_module/_03693_ ),
    .Y(\reg_module/_03694_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10980_  (.A(\reg_module/_03690_ ),
    .B(\reg_module/_03694_ ),
    .Y(\reg_module/_03695_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10981_  (.A(\reg_module/_03695_ ),
    .B(net435),
    .Y(\reg_module/_03696_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10982_  (.A(\reg_module/_03540_ ),
    .B(\reg_module/gprf[174] ),
    .Y(\reg_module/_03697_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10983_  (.A(\reg_module/gprf[142] ),
    .B(net618),
    .Y(\reg_module/_03698_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10984_  (.A(\reg_module/_03697_ ),
    .B(net496),
    .C(\reg_module/_03698_ ),
    .Y(\reg_module/_03699_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10985_  (.A(\reg_module/_03544_ ),
    .B(\reg_module/gprf[238] ),
    .Y(\reg_module/_03700_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10986_  (.A(\reg_module/gprf[206] ),
    .B(net617),
    .Y(\reg_module/_03701_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10987_  (.A(\reg_module/_03700_ ),
    .B(\reg_module/_03391_ ),
    .C(\reg_module/_03701_ ),
    .Y(\reg_module/_03702_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10988_  (.A(\reg_module/_03699_ ),
    .B(\reg_module/_03702_ ),
    .Y(\reg_module/_03703_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10989_  (.A(\reg_module/_03703_ ),
    .B(\reg_module/_03549_ ),
    .Y(\reg_module/_03704_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10990_  (.A(\reg_module/_03696_ ),
    .B(\reg_module/_03704_ ),
    .C(net401),
    .Y(\reg_module/_03705_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10991_  (.A(\reg_module/_03687_ ),
    .B(\reg_module/_03705_ ),
    .Y(\reg_module/_03706_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10992_  (.A(\reg_module/_03706_ ),
    .B(net384),
    .Y(\reg_module/_03707_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10993_  (.A(\reg_module/_03667_ ),
    .B(\reg_module/_03707_ ),
    .Y(\wRs2Data[14] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10994_  (.A(\reg_module/_03471_ ),
    .B(\reg_module/gprf[815] ),
    .Y(\reg_module/_03708_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10995_  (.A(\reg_module/gprf[783] ),
    .B(net624),
    .Y(\reg_module/_03709_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10996_  (.A(\reg_module/_03708_ ),
    .B(net499),
    .C(\reg_module/_03709_ ),
    .Y(\reg_module/_03710_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10997_  (.A(\reg_module/_03475_ ),
    .B(\reg_module/gprf[879] ),
    .Y(\reg_module/_03711_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_10998_  (.A(\reg_module/gprf[847] ),
    .B(net622),
    .Y(\reg_module/_03712_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_10999_  (.A(\reg_module/_03711_ ),
    .B(\reg_module/_03477_ ),
    .C(\reg_module/_03712_ ),
    .Y(\reg_module/_03713_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11000_  (.A(\reg_module/_03710_ ),
    .B(\reg_module/_03713_ ),
    .Y(\reg_module/_03714_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11001_  (.A(\reg_module/_03714_ ),
    .B(net433),
    .Y(\reg_module/_03715_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11002_  (.A(\reg_module/_03326_ ),
    .B(\reg_module/gprf[943] ),
    .Y(\reg_module/_03716_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11003_  (.A(\reg_module/gprf[911] ),
    .B(net607),
    .Y(\reg_module/_03717_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11004_  (.A(\reg_module/_03716_ ),
    .B(net491),
    .C(\reg_module/_03717_ ),
    .Y(\reg_module/_03718_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11005_  (.A(\reg_module/_03330_ ),
    .B(\reg_module/gprf[1007] ),
    .Y(\reg_module/_03719_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11006_  (.A(\reg_module/gprf[975] ),
    .B(net607),
    .Y(\reg_module/_03720_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11007_  (.A(\reg_module/_03719_ ),
    .B(\reg_module/_03486_ ),
    .C(\reg_module/_03720_ ),
    .Y(\reg_module/_03721_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11008_  (.A(\reg_module/_03718_ ),
    .B(\reg_module/_03721_ ),
    .Y(\reg_module/_03722_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11009_  (.A(\reg_module/_03722_ ),
    .B(\reg_module/_03642_ ),
    .Y(\reg_module/_03723_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11010_  (.A(\reg_module/_03715_ ),
    .B(\reg_module/_03723_ ),
    .C(\reg_module/_03260_ ),
    .Y(\reg_module/_03724_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11011_  (.A(\reg_module/_03645_ ),
    .B(\reg_module/gprf[687] ),
    .Y(\reg_module/_03725_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11012_  (.A(\reg_module/gprf[655] ),
    .B(net599),
    .Y(\reg_module/_03726_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11013_  (.A(\reg_module/_03725_ ),
    .B(net486),
    .C(\reg_module/_03726_ ),
    .Y(\reg_module/_03727_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11014_  (.A(\reg_module/_03340_ ),
    .B(\reg_module/gprf[751] ),
    .Y(\reg_module/_03728_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11015_  (.A(\reg_module/gprf[719] ),
    .B(net599),
    .Y(\reg_module/_03729_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11016_  (.A(\reg_module/_03728_ ),
    .B(\reg_module/_03650_ ),
    .C(\reg_module/_03729_ ),
    .Y(\reg_module/_03730_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11017_  (.A(\reg_module/_03727_ ),
    .B(\reg_module/_03730_ ),
    .Y(\reg_module/_03731_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11018_  (.A(\reg_module/_03731_ ),
    .B(\reg_module/_03269_ ),
    .Y(\reg_module/_03732_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11019_  (.A(\reg_module/_03500_ ),
    .B(\reg_module/gprf[559] ),
    .Y(\reg_module/_03733_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11020_  (.A(\reg_module/gprf[527] ),
    .B(net626),
    .Y(\reg_module/_03734_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11021_  (.A(\reg_module/_03733_ ),
    .B(net500),
    .C(\reg_module/_03734_ ),
    .Y(\reg_module/_03735_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11022_  (.A(\reg_module/_03658_ ),
    .B(\reg_module/gprf[623] ),
    .Y(\reg_module/_03736_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11023_  (.A(\reg_module/gprf[591] ),
    .B(net626),
    .Y(\reg_module/_03737_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11024_  (.A(\reg_module/_03736_ ),
    .B(\reg_module/_03505_ ),
    .C(\reg_module/_03737_ ),
    .Y(\reg_module/_03738_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11025_  (.A(\reg_module/_03735_ ),
    .B(\reg_module/_03738_ ),
    .Y(\reg_module/_03739_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11026_  (.A(\reg_module/_03739_ ),
    .B(net434),
    .Y(\reg_module/_03740_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11027_  (.A(\reg_module/_03732_ ),
    .B(\reg_module/_03740_ ),
    .C(net400),
    .Y(\reg_module/_03741_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11028_  (.A(\reg_module/_03724_ ),
    .B(\reg_module/_03741_ ),
    .Y(\reg_module/_03742_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11029_  (.A(\reg_module/_03742_ ),
    .B(\reg_module/_03512_ ),
    .Y(\reg_module/_03743_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11030_  (.A(\reg_module/_03357_ ),
    .B(\reg_module/gprf[303] ),
    .Y(\reg_module/_03744_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11031_  (.A(\reg_module/gprf[271] ),
    .B(net624),
    .Y(\reg_module/_03745_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11032_  (.A(\reg_module/_03744_ ),
    .B(net499),
    .C(\reg_module/_03745_ ),
    .Y(\reg_module/_03746_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11033_  (.A(\reg_module/_03593_ ),
    .B(\reg_module/gprf[367] ),
    .Y(\reg_module/_03747_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11034_  (.A(\reg_module/gprf[335] ),
    .B(net625),
    .Y(\reg_module/_03748_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11035_  (.A(\reg_module/_03747_ ),
    .B(\reg_module/_03363_ ),
    .C(\reg_module/_03748_ ),
    .Y(\reg_module/_03749_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11036_  (.A(\reg_module/_03746_ ),
    .B(\reg_module/_03749_ ),
    .Y(\reg_module/_03750_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11037_  (.A(\reg_module/_03750_ ),
    .B(net436),
    .Y(\reg_module/_03751_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11038_  (.A(\reg_module/_03676_ ),
    .B(\reg_module/gprf[431] ),
    .Y(\reg_module/_03752_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11039_  (.A(\reg_module/gprf[399] ),
    .B(net604),
    .Y(\reg_module/_03753_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11040_  (.A(\reg_module/_03752_ ),
    .B(net489),
    .C(\reg_module/_03753_ ),
    .Y(\reg_module/_03754_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11041_  (.A(\reg_module/_03371_ ),
    .B(\reg_module/gprf[495] ),
    .Y(\reg_module/_03755_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11042_  (.A(\reg_module/gprf[463] ),
    .B(net604),
    .Y(\reg_module/_03756_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11043_  (.A(\reg_module/_03755_ ),
    .B(\reg_module/_03681_ ),
    .C(\reg_module/_03756_ ),
    .Y(\reg_module/_03757_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11044_  (.A(\reg_module/_03754_ ),
    .B(\reg_module/_03757_ ),
    .Y(\reg_module/_03758_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11045_  (.A(\reg_module/_03758_ ),
    .B(\reg_module/_03529_ ),
    .Y(\reg_module/_03759_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11046_  (.A(\reg_module/_03751_ ),
    .B(\reg_module/_03759_ ),
    .C(\reg_module/_03686_ ),
    .Y(\reg_module/_03760_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11047_  (.A(\reg_module/_03593_ ),
    .B(\reg_module/gprf[47] ),
    .Y(\reg_module/_03761_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11048_  (.A(\reg_module/gprf[15] ),
    .B(net628),
    .Y(\reg_module/_03762_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11049_  (.A(\reg_module/_03761_ ),
    .B(net501),
    .C(\reg_module/_03762_ ),
    .Y(\reg_module/_03763_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11050_  (.A(\reg_module/_03691_ ),
    .B(\reg_module/gprf[111] ),
    .Y(\reg_module/_03764_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11051_  (.A(\reg_module/gprf[79] ),
    .B(net627),
    .Y(\reg_module/_03765_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11052_  (.A(\reg_module/_03764_ ),
    .B(\reg_module/_03382_ ),
    .C(\reg_module/_03765_ ),
    .Y(\reg_module/_03766_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11053_  (.A(\reg_module/_03763_ ),
    .B(\reg_module/_03766_ ),
    .Y(\reg_module/_03767_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11054_  (.A(\reg_module/_03767_ ),
    .B(net435),
    .Y(\reg_module/_03768_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11055_  (.A(\reg_module/_03540_ ),
    .B(\reg_module/gprf[175] ),
    .Y(\reg_module/_03769_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11056_  (.A(\reg_module/gprf[143] ),
    .B(net617),
    .Y(\reg_module/_03770_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11057_  (.A(\reg_module/_03769_ ),
    .B(net496),
    .C(\reg_module/_03770_ ),
    .Y(\reg_module/_03771_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11058_  (.A(\reg_module/_03544_ ),
    .B(\reg_module/gprf[239] ),
    .Y(\reg_module/_03772_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11059_  (.A(\reg_module/gprf[207] ),
    .B(net618),
    .Y(\reg_module/_03773_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11060_  (.A(\reg_module/_03772_ ),
    .B(\reg_module/_03391_ ),
    .C(\reg_module/_03773_ ),
    .Y(\reg_module/_03774_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11061_  (.A(\reg_module/_03771_ ),
    .B(\reg_module/_03774_ ),
    .Y(\reg_module/_03775_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11062_  (.A(\reg_module/_03775_ ),
    .B(\reg_module/_03549_ ),
    .Y(\reg_module/_03776_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11063_  (.A(\reg_module/_03768_ ),
    .B(\reg_module/_03776_ ),
    .C(net401),
    .Y(\reg_module/_03777_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11064_  (.A(\reg_module/_03760_ ),
    .B(\reg_module/_03777_ ),
    .Y(\reg_module/_03778_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11065_  (.A(\reg_module/_03778_ ),
    .B(net385),
    .Y(\reg_module/_03779_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11066_  (.A(\reg_module/_03743_ ),
    .B(\reg_module/_03779_ ),
    .Y(\wRs2Data[15] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11067_  (.A(\reg_module/_03471_ ),
    .B(\reg_module/gprf[816] ),
    .Y(\reg_module/_03780_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11068_  (.A(\reg_module/gprf[784] ),
    .B(net609),
    .Y(\reg_module/_03781_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11069_  (.A(\reg_module/_03780_ ),
    .B(net492),
    .C(\reg_module/_03781_ ),
    .Y(\reg_module/_03782_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11070_  (.A(\reg_module/_03475_ ),
    .B(\reg_module/gprf[880] ),
    .Y(\reg_module/_03783_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11071_  (.A(\reg_module/gprf[848] ),
    .B(net622),
    .Y(\reg_module/_03784_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11072_  (.A(\reg_module/_03783_ ),
    .B(\reg_module/_03477_ ),
    .C(\reg_module/_03784_ ),
    .Y(\reg_module/_03785_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11073_  (.A(\reg_module/_03782_ ),
    .B(\reg_module/_03785_ ),
    .Y(\reg_module/_03786_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11074_  (.A(\reg_module/_03786_ ),
    .B(net428),
    .Y(\reg_module/_03787_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11075_  (.A(\reg_module/_02570_ ),
    .X(\reg_module/_03788_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11076_  (.A(\reg_module/_03788_ ),
    .B(\reg_module/gprf[944] ),
    .Y(\reg_module/_03789_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11077_  (.A(\reg_module/gprf[912] ),
    .B(net607),
    .Y(\reg_module/_03790_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11078_  (.A(\reg_module/_03789_ ),
    .B(net491),
    .C(\reg_module/_03790_ ),
    .Y(\reg_module/_03791_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11079_  (.A(\reg_module/_02513_ ),
    .X(\reg_module/_03792_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11080_  (.A(\reg_module/_03792_ ),
    .B(\reg_module/gprf[1008] ),
    .Y(\reg_module/_03793_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11081_  (.A(\reg_module/gprf[976] ),
    .B(net607),
    .Y(\reg_module/_03794_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11082_  (.A(\reg_module/_03793_ ),
    .B(\reg_module/_03486_ ),
    .C(\reg_module/_03794_ ),
    .Y(\reg_module/_03795_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11083_  (.A(\reg_module/_03791_ ),
    .B(\reg_module/_03795_ ),
    .Y(\reg_module/_03796_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11084_  (.A(\reg_module/_03796_ ),
    .B(\reg_module/_03642_ ),
    .Y(\reg_module/_03797_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11085_  (.A(\reg_module/_03787_ ),
    .B(\reg_module/_03797_ ),
    .C(\reg_module/_03260_ ),
    .Y(\reg_module/_03798_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11086_  (.A(\reg_module/_03645_ ),
    .B(\reg_module/gprf[688] ),
    .Y(\reg_module/_03799_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11087_  (.A(\reg_module/gprf[656] ),
    .B(net594),
    .Y(\reg_module/_03800_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11088_  (.A(\reg_module/_03799_ ),
    .B(net485),
    .C(\reg_module/_03800_ ),
    .Y(\reg_module/_03801_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_11089_  (.A(\reg_module/_02579_ ),
    .X(\reg_module/_03802_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11090_  (.A(\reg_module/_03802_ ),
    .B(\reg_module/gprf[752] ),
    .Y(\reg_module/_03803_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11091_  (.A(\reg_module/gprf[720] ),
    .B(net600),
    .Y(\reg_module/_03804_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11092_  (.A(\reg_module/_03803_ ),
    .B(\reg_module/_03650_ ),
    .C(\reg_module/_03804_ ),
    .Y(\reg_module/_03805_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11093_  (.A(\reg_module/_03801_ ),
    .B(\reg_module/_03805_ ),
    .Y(\reg_module/_03806_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11094_  (.A(\reg_module/_03806_ ),
    .B(\reg_module/_03269_ ),
    .Y(\reg_module/_03807_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11095_  (.A(\reg_module/_03500_ ),
    .B(\reg_module/gprf[560] ),
    .Y(\reg_module/_03808_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11096_  (.A(\reg_module/gprf[528] ),
    .B(net626),
    .Y(\reg_module/_03809_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11097_  (.A(\reg_module/_03808_ ),
    .B(net500),
    .C(\reg_module/_03809_ ),
    .Y(\reg_module/_03810_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11098_  (.A(\reg_module/_03658_ ),
    .B(\reg_module/gprf[624] ),
    .Y(\reg_module/_03811_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11099_  (.A(\reg_module/gprf[592] ),
    .B(net626),
    .Y(\reg_module/_03812_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11100_  (.A(\reg_module/_03811_ ),
    .B(\reg_module/_03505_ ),
    .C(\reg_module/_03812_ ),
    .Y(\reg_module/_03813_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11101_  (.A(\reg_module/_03810_ ),
    .B(\reg_module/_03813_ ),
    .Y(\reg_module/_03814_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11102_  (.A(\reg_module/_03814_ ),
    .B(net434),
    .Y(\reg_module/_03815_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11103_  (.A(\reg_module/_03807_ ),
    .B(\reg_module/_03815_ ),
    .C(net399),
    .Y(\reg_module/_03816_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11104_  (.A(\reg_module/_03798_ ),
    .B(\reg_module/_03816_ ),
    .Y(\reg_module/_03817_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11105_  (.A(\reg_module/_03817_ ),
    .B(\reg_module/_03512_ ),
    .Y(\reg_module/_03818_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11106_  (.A(\reg_module/_02565_ ),
    .X(\reg_module/_03819_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11107_  (.A(\reg_module/_03819_ ),
    .B(\reg_module/gprf[304] ),
    .Y(\reg_module/_03820_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11108_  (.A(\reg_module/gprf[272] ),
    .B(net609),
    .Y(\reg_module/_03821_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11109_  (.A(\reg_module/_03820_ ),
    .B(net491),
    .C(\reg_module/_03821_ ),
    .Y(\reg_module/_03822_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11110_  (.A(\reg_module/_02897_ ),
    .X(\reg_module/_03823_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11111_  (.A(\reg_module/_03823_ ),
    .B(\reg_module/gprf[368] ),
    .Y(\reg_module/_03824_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11112_  (.A(\reg_module/_02538_ ),
    .X(\reg_module/_03825_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11113_  (.A(\reg_module/gprf[336] ),
    .B(net609),
    .Y(\reg_module/_03826_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11114_  (.A(\reg_module/_03824_ ),
    .B(\reg_module/_03825_ ),
    .C(\reg_module/_03826_ ),
    .Y(\reg_module/_03827_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11115_  (.A(\reg_module/_03822_ ),
    .B(\reg_module/_03827_ ),
    .Y(\reg_module/_03828_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11116_  (.A(\reg_module/_03828_ ),
    .B(net428),
    .Y(\reg_module/_03829_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11117_  (.A(\reg_module/_03676_ ),
    .B(\reg_module/gprf[432] ),
    .Y(\reg_module/_03830_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11118_  (.A(\reg_module/gprf[400] ),
    .B(net606),
    .Y(\reg_module/_03831_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11119_  (.A(\reg_module/_03830_ ),
    .B(net490),
    .C(\reg_module/_03831_ ),
    .Y(\reg_module/_03832_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11120_  (.A(\reg_module/_02550_ ),
    .X(\reg_module/_03833_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11121_  (.A(\reg_module/_03833_ ),
    .B(\reg_module/gprf[496] ),
    .Y(\reg_module/_03834_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11122_  (.A(\reg_module/gprf[464] ),
    .B(net603),
    .Y(\reg_module/_03835_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11123_  (.A(\reg_module/_03834_ ),
    .B(\reg_module/_03681_ ),
    .C(\reg_module/_03835_ ),
    .Y(\reg_module/_03836_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11124_  (.A(\reg_module/_03832_ ),
    .B(\reg_module/_03836_ ),
    .Y(\reg_module/_03837_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11125_  (.A(\reg_module/_03837_ ),
    .B(\reg_module/_03529_ ),
    .Y(\reg_module/_03838_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11126_  (.A(\reg_module/_03829_ ),
    .B(\reg_module/_03838_ ),
    .C(\reg_module/_03686_ ),
    .Y(\reg_module/_03839_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11127_  (.A(\reg_module/_03823_ ),
    .B(\reg_module/gprf[48] ),
    .Y(\reg_module/_03840_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11128_  (.A(\reg_module/gprf[16] ),
    .B(net628),
    .Y(\reg_module/_03841_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11129_  (.A(\reg_module/_03840_ ),
    .B(net501),
    .C(\reg_module/_03841_ ),
    .Y(\reg_module/_03842_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11130_  (.A(\reg_module/_03691_ ),
    .B(\reg_module/gprf[112] ),
    .Y(\reg_module/_03843_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11131_  (.A(\reg_module/_02604_ ),
    .X(\reg_module/_03844_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11132_  (.A(\reg_module/gprf[80] ),
    .B(net628),
    .Y(\reg_module/_03845_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11133_  (.A(\reg_module/_03843_ ),
    .B(\reg_module/_03844_ ),
    .C(\reg_module/_03845_ ),
    .Y(\reg_module/_03846_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11134_  (.A(\reg_module/_03842_ ),
    .B(\reg_module/_03846_ ),
    .Y(\reg_module/_03847_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11135_  (.A(\reg_module/_03847_ ),
    .B(net434),
    .Y(\reg_module/_03848_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11136_  (.A(\reg_module/_03540_ ),
    .B(\reg_module/gprf[176] ),
    .Y(\reg_module/_03849_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11137_  (.A(\reg_module/gprf[144] ),
    .B(net617),
    .Y(\reg_module/_03850_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11138_  (.A(\reg_module/_03849_ ),
    .B(net495),
    .C(\reg_module/_03850_ ),
    .Y(\reg_module/_03851_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11139_  (.A(\reg_module/_03544_ ),
    .B(\reg_module/gprf[240] ),
    .Y(\reg_module/_03852_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_11140_  (.A(\reg_module/_02502_ ),
    .X(\reg_module/_03853_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11141_  (.A(\reg_module/gprf[208] ),
    .B(net615),
    .Y(\reg_module/_03854_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11142_  (.A(\reg_module/_03852_ ),
    .B(\reg_module/_03853_ ),
    .C(\reg_module/_03854_ ),
    .Y(\reg_module/_03855_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11143_  (.A(\reg_module/_03851_ ),
    .B(\reg_module/_03855_ ),
    .Y(\reg_module/_03856_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11144_  (.A(\reg_module/_03856_ ),
    .B(\reg_module/_03549_ ),
    .Y(\reg_module/_03857_ ));
 sky130_fd_sc_hd__nand3_2 \reg_module/_11145_  (.A(\reg_module/_03848_ ),
    .B(\reg_module/_03857_ ),
    .C(net401),
    .Y(\reg_module/_03858_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11146_  (.A(\reg_module/_03839_ ),
    .B(\reg_module/_03858_ ),
    .Y(\reg_module/_03859_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11147_  (.A(\reg_module/_03859_ ),
    .B(net385),
    .Y(\reg_module/_03860_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11148_  (.A(\reg_module/_03818_ ),
    .B(\reg_module/_03860_ ),
    .Y(\wRs2Data[16] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11149_  (.A(\reg_module/_03471_ ),
    .B(\reg_module/gprf[561] ),
    .Y(\reg_module/_03861_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11150_  (.A(\reg_module/gprf[529] ),
    .B(net622),
    .Y(\reg_module/_03862_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11151_  (.A(\reg_module/_03861_ ),
    .B(net498),
    .C(\reg_module/_03862_ ),
    .Y(\reg_module/_03863_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11152_  (.A(\reg_module/_03475_ ),
    .B(\reg_module/gprf[625] ),
    .Y(\reg_module/_03864_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11153_  (.A(\reg_module/gprf[593] ),
    .B(net623),
    .Y(\reg_module/_03865_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11154_  (.A(\reg_module/_03864_ ),
    .B(\reg_module/_03477_ ),
    .C(\reg_module/_03865_ ),
    .Y(\reg_module/_03866_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11155_  (.A(\reg_module/_03863_ ),
    .B(\reg_module/_03866_ ),
    .Y(\reg_module/_03867_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11156_  (.A(\reg_module/_03867_ ),
    .B(net429),
    .Y(\reg_module/_03868_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11157_  (.A(\reg_module/_03788_ ),
    .B(\reg_module/gprf[689] ),
    .Y(\reg_module/_03869_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11158_  (.A(\reg_module/gprf[657] ),
    .B(net595),
    .Y(\reg_module/_03870_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11159_  (.A(\reg_module/_03869_ ),
    .B(net488),
    .C(\reg_module/_03870_ ),
    .Y(\reg_module/_03871_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11160_  (.A(\reg_module/_03792_ ),
    .B(\reg_module/gprf[753] ),
    .Y(\reg_module/_03872_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11161_  (.A(\reg_module/gprf[721] ),
    .B(net599),
    .Y(\reg_module/_03873_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11162_  (.A(\reg_module/_03872_ ),
    .B(\reg_module/_03486_ ),
    .C(\reg_module/_03873_ ),
    .Y(\reg_module/_03874_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11163_  (.A(\reg_module/_03871_ ),
    .B(\reg_module/_03874_ ),
    .Y(\reg_module/_03875_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11164_  (.A(\reg_module/_03875_ ),
    .B(\reg_module/_03642_ ),
    .Y(\reg_module/_03876_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11165_  (.A(\reg_module/_03868_ ),
    .B(\reg_module/_03876_ ),
    .C(net399),
    .Y(\reg_module/_03877_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11166_  (.A(\reg_module/_03645_ ),
    .B(\reg_module/gprf[817] ),
    .Y(\reg_module/_03878_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11167_  (.A(\reg_module/gprf[785] ),
    .B(net610),
    .Y(\reg_module/_03879_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11168_  (.A(\reg_module/_03878_ ),
    .B(net492),
    .C(\reg_module/_03879_ ),
    .Y(\reg_module/_03880_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11169_  (.A(\reg_module/_03802_ ),
    .B(\reg_module/gprf[881] ),
    .Y(\reg_module/_03881_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11170_  (.A(\reg_module/gprf[849] ),
    .B(net608),
    .Y(\reg_module/_03882_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11171_  (.A(\reg_module/_03881_ ),
    .B(\reg_module/_03650_ ),
    .C(\reg_module/_03882_ ),
    .Y(\reg_module/_03883_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11172_  (.A(\reg_module/_03880_ ),
    .B(\reg_module/_03883_ ),
    .Y(\reg_module/_03884_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11173_  (.A(\reg_module/_03884_ ),
    .B(net428),
    .Y(\reg_module/_03885_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11174_  (.A(\reg_module/_03500_ ),
    .B(\reg_module/gprf[945] ),
    .Y(\reg_module/_03886_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11175_  (.A(\reg_module/gprf[913] ),
    .B(net607),
    .Y(\reg_module/_03887_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11176_  (.A(\reg_module/_03886_ ),
    .B(net491),
    .C(\reg_module/_03887_ ),
    .Y(\reg_module/_03888_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11177_  (.A(\reg_module/_03658_ ),
    .B(\reg_module/gprf[1009] ),
    .Y(\reg_module/_03889_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11178_  (.A(\reg_module/gprf[977] ),
    .B(net607),
    .Y(\reg_module/_03890_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11179_  (.A(\reg_module/_03889_ ),
    .B(\reg_module/_03505_ ),
    .C(\reg_module/_03890_ ),
    .Y(\reg_module/_03891_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11180_  (.A(\reg_module/_03888_ ),
    .B(\reg_module/_03891_ ),
    .Y(\reg_module/_03892_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11181_  (.A(\reg_module/_03892_ ),
    .B(\reg_module/_03663_ ),
    .Y(\reg_module/_03893_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11182_  (.A(\reg_module/_03885_ ),
    .B(\reg_module/_03893_ ),
    .C(\reg_module/_02738_ ),
    .Y(\reg_module/_03894_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11183_  (.A(\reg_module/_03877_ ),
    .B(\reg_module/_03894_ ),
    .Y(\reg_module/_03895_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11184_  (.A(\reg_module/_03895_ ),
    .B(\reg_module/_03512_ ),
    .Y(\reg_module/_03896_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11185_  (.A(\reg_module/_03819_ ),
    .B(\reg_module/gprf[305] ),
    .Y(\reg_module/_03897_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11186_  (.A(\reg_module/gprf[273] ),
    .B(net609),
    .Y(\reg_module/_03898_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11187_  (.A(\reg_module/_03897_ ),
    .B(net492),
    .C(\reg_module/_03898_ ),
    .Y(\reg_module/_03899_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11188_  (.A(\reg_module/_03823_ ),
    .B(\reg_module/gprf[369] ),
    .Y(\reg_module/_03900_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11189_  (.A(\reg_module/gprf[337] ),
    .B(net609),
    .Y(\reg_module/_03901_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11190_  (.A(\reg_module/_03900_ ),
    .B(\reg_module/_03825_ ),
    .C(\reg_module/_03901_ ),
    .Y(\reg_module/_03902_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11191_  (.A(\reg_module/_03899_ ),
    .B(\reg_module/_03902_ ),
    .Y(\reg_module/_03903_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11192_  (.A(\reg_module/_03903_ ),
    .B(net428),
    .Y(\reg_module/_03904_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11193_  (.A(\reg_module/_03676_ ),
    .B(\reg_module/gprf[433] ),
    .Y(\reg_module/_03905_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11194_  (.A(\reg_module/gprf[401] ),
    .B(net604),
    .Y(\reg_module/_03906_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11195_  (.A(\reg_module/_03905_ ),
    .B(net489),
    .C(\reg_module/_03906_ ),
    .Y(\reg_module/_03907_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11196_  (.A(\reg_module/_03833_ ),
    .B(\reg_module/gprf[497] ),
    .Y(\reg_module/_03908_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11197_  (.A(\reg_module/gprf[465] ),
    .B(net604),
    .Y(\reg_module/_03909_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11198_  (.A(\reg_module/_03908_ ),
    .B(\reg_module/_03681_ ),
    .C(\reg_module/_03909_ ),
    .Y(\reg_module/_03910_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11199_  (.A(\reg_module/_03907_ ),
    .B(\reg_module/_03910_ ),
    .Y(\reg_module/_03911_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11200_  (.A(\reg_module/_03911_ ),
    .B(\reg_module/_03529_ ),
    .Y(\reg_module/_03912_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11201_  (.A(\reg_module/_03904_ ),
    .B(\reg_module/_03912_ ),
    .C(\reg_module/_03686_ ),
    .Y(\reg_module/_03913_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11202_  (.A(\reg_module/_03823_ ),
    .B(\reg_module/gprf[49] ),
    .Y(\reg_module/_03914_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11203_  (.A(\reg_module/gprf[17] ),
    .B(net628),
    .Y(\reg_module/_03915_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11204_  (.A(\reg_module/_03914_ ),
    .B(net501),
    .C(\reg_module/_03915_ ),
    .Y(\reg_module/_03916_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11205_  (.A(\reg_module/_03691_ ),
    .B(\reg_module/gprf[113] ),
    .Y(\reg_module/_03917_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11206_  (.A(\reg_module/gprf[81] ),
    .B(net628),
    .Y(\reg_module/_03918_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11207_  (.A(\reg_module/_03917_ ),
    .B(\reg_module/_03844_ ),
    .C(\reg_module/_03918_ ),
    .Y(\reg_module/_03919_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11208_  (.A(\reg_module/_03916_ ),
    .B(\reg_module/_03919_ ),
    .Y(\reg_module/_03920_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11209_  (.A(\reg_module/_03920_ ),
    .B(net434),
    .Y(\reg_module/_03921_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11210_  (.A(\reg_module/_03540_ ),
    .B(\reg_module/gprf[177] ),
    .Y(\reg_module/_03922_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11211_  (.A(\reg_module/gprf[145] ),
    .B(net617),
    .Y(\reg_module/_03923_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11212_  (.A(\reg_module/_03922_ ),
    .B(net496),
    .C(\reg_module/_03923_ ),
    .Y(\reg_module/_03924_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11213_  (.A(\reg_module/_03544_ ),
    .B(\reg_module/gprf[241] ),
    .Y(\reg_module/_03925_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11214_  (.A(\reg_module/gprf[209] ),
    .B(net619),
    .Y(\reg_module/_03926_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11215_  (.A(\reg_module/_03925_ ),
    .B(\reg_module/_03853_ ),
    .C(\reg_module/_03926_ ),
    .Y(\reg_module/_03927_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11216_  (.A(\reg_module/_03924_ ),
    .B(\reg_module/_03927_ ),
    .Y(\reg_module/_03928_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11217_  (.A(\reg_module/_03928_ ),
    .B(\reg_module/_03549_ ),
    .Y(\reg_module/_03929_ ));
 sky130_fd_sc_hd__nand3_2 \reg_module/_11218_  (.A(\reg_module/_03921_ ),
    .B(\reg_module/_03929_ ),
    .C(net401),
    .Y(\reg_module/_03930_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11219_  (.A(\reg_module/_03913_ ),
    .B(\reg_module/_03930_ ),
    .Y(\reg_module/_03931_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11220_  (.A(\reg_module/_03931_ ),
    .B(net384),
    .Y(\reg_module/_03932_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11221_  (.A(\reg_module/_03896_ ),
    .B(\reg_module/_03932_ ),
    .Y(\wRs2Data[17] ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11222_  (.A(\reg_module/_02492_ ),
    .X(\reg_module/_03933_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11223_  (.A(\reg_module/_03933_ ),
    .B(\reg_module/gprf[818] ),
    .Y(\reg_module/_03934_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11224_  (.A(\reg_module/gprf[786] ),
    .B(net556),
    .Y(\reg_module/_03935_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11225_  (.A(\reg_module/_03934_ ),
    .B(net465),
    .C(\reg_module/_03935_ ),
    .Y(\reg_module/_03936_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11226_  (.A(\reg_module/_02498_ ),
    .X(\reg_module/_03937_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11227_  (.A(\reg_module/_03937_ ),
    .B(\reg_module/gprf[882] ),
    .Y(\reg_module/_03938_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11228_  (.A(\reg_module/_02573_ ),
    .X(\reg_module/_03939_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11229_  (.A(\reg_module/gprf[850] ),
    .B(net556),
    .Y(\reg_module/_03940_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11230_  (.A(\reg_module/_03938_ ),
    .B(\reg_module/_03939_ ),
    .C(\reg_module/_03940_ ),
    .Y(\reg_module/_03941_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11231_  (.A(\reg_module/_03936_ ),
    .B(\reg_module/_03941_ ),
    .Y(\reg_module/_03942_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11232_  (.A(\reg_module/_03942_ ),
    .B(net417),
    .Y(\reg_module/_03943_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11233_  (.A(\reg_module/_03788_ ),
    .B(\reg_module/gprf[946] ),
    .Y(\reg_module/_03944_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11234_  (.A(\reg_module/gprf[914] ),
    .B(net548),
    .Y(\reg_module/_03945_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11235_  (.A(\reg_module/_03944_ ),
    .B(net461),
    .C(\reg_module/_03945_ ),
    .Y(\reg_module/_03946_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11236_  (.A(\reg_module/_03792_ ),
    .B(\reg_module/gprf[1010] ),
    .Y(\reg_module/_03947_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11237_  (.A(\reg_module/_02516_ ),
    .X(\reg_module/_03948_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11238_  (.A(\reg_module/gprf[978] ),
    .B(net595),
    .Y(\reg_module/_03949_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11239_  (.A(\reg_module/_03947_ ),
    .B(\reg_module/_03948_ ),
    .C(\reg_module/_03949_ ),
    .Y(\reg_module/_03950_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11240_  (.A(\reg_module/_03946_ ),
    .B(\reg_module/_03950_ ),
    .Y(\reg_module/_03951_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11241_  (.A(\reg_module/_03951_ ),
    .B(\reg_module/_03642_ ),
    .Y(\reg_module/_03952_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11242_  (.A(\reg_module/_02595_ ),
    .X(\reg_module/_03953_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11243_  (.A(\reg_module/_03943_ ),
    .B(\reg_module/_03952_ ),
    .C(\reg_module/_03953_ ),
    .Y(\reg_module/_03954_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11244_  (.A(\reg_module/_03645_ ),
    .B(\reg_module/gprf[690] ),
    .Y(\reg_module/_03955_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11245_  (.A(\reg_module/gprf[658] ),
    .B(net594),
    .Y(\reg_module/_03956_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11246_  (.A(\reg_module/_03955_ ),
    .B(net485),
    .C(\reg_module/_03956_ ),
    .Y(\reg_module/_03957_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11247_  (.A(\reg_module/_03802_ ),
    .B(\reg_module/gprf[754] ),
    .Y(\reg_module/_03958_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11248_  (.A(\reg_module/gprf[722] ),
    .B(net595),
    .Y(\reg_module/_03959_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11249_  (.A(\reg_module/_03958_ ),
    .B(\reg_module/_03650_ ),
    .C(\reg_module/_03959_ ),
    .Y(\reg_module/_03960_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11250_  (.A(\reg_module/_03957_ ),
    .B(\reg_module/_03960_ ),
    .Y(\reg_module/_03961_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11251_  (.A(\reg_module/_02523_ ),
    .X(\reg_module/_03962_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11252_  (.A(\reg_module/_03961_ ),
    .B(\reg_module/_03962_ ),
    .Y(\reg_module/_03963_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11253_  (.A(\reg_module/_02545_ ),
    .X(\reg_module/_03964_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11254_  (.A(\reg_module/_03964_ ),
    .B(\reg_module/gprf[562] ),
    .Y(\reg_module/_03965_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11255_  (.A(\reg_module/gprf[530] ),
    .B(net555),
    .Y(\reg_module/_03966_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11256_  (.A(\reg_module/_03965_ ),
    .B(net465),
    .C(\reg_module/_03966_ ),
    .Y(\reg_module/_03967_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11257_  (.A(\reg_module/_03658_ ),
    .B(\reg_module/gprf[626] ),
    .Y(\reg_module/_03968_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11258_  (.A(\reg_module/_02553_ ),
    .X(\reg_module/_03969_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11259_  (.A(\reg_module/gprf[594] ),
    .B(net556),
    .Y(\reg_module/_03970_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11260_  (.A(\reg_module/_03968_ ),
    .B(\reg_module/_03969_ ),
    .C(\reg_module/_03970_ ),
    .Y(\reg_module/_03971_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11261_  (.A(\reg_module/_03967_ ),
    .B(\reg_module/_03971_ ),
    .Y(\reg_module/_03972_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11262_  (.A(\reg_module/_03972_ ),
    .B(net417),
    .Y(\reg_module/_03973_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11263_  (.A(\reg_module/_03963_ ),
    .B(\reg_module/_03973_ ),
    .C(net392),
    .Y(\reg_module/_03974_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11264_  (.A(\reg_module/_03954_ ),
    .B(\reg_module/_03974_ ),
    .Y(\reg_module/_03975_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11265_  (.A(\reg_module/_02562_ ),
    .X(\reg_module/_03976_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11266_  (.A(\reg_module/_03975_ ),
    .B(\reg_module/_03976_ ),
    .Y(\reg_module/_03977_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11267_  (.A(\reg_module/_03819_ ),
    .B(\reg_module/gprf[306] ),
    .Y(\reg_module/_03978_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11268_  (.A(\reg_module/gprf[274] ),
    .B(net605),
    .Y(\reg_module/_03979_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11269_  (.A(\reg_module/_03978_ ),
    .B(net489),
    .C(\reg_module/_03979_ ),
    .Y(\reg_module/_03980_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11270_  (.A(\reg_module/_03823_ ),
    .B(\reg_module/gprf[370] ),
    .Y(\reg_module/_03981_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11271_  (.A(\reg_module/gprf[338] ),
    .B(net605),
    .Y(\reg_module/_03982_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11272_  (.A(\reg_module/_03981_ ),
    .B(\reg_module/_03825_ ),
    .C(\reg_module/_03982_ ),
    .Y(\reg_module/_03983_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11273_  (.A(\reg_module/_03980_ ),
    .B(\reg_module/_03983_ ),
    .Y(\reg_module/_03984_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11274_  (.A(\reg_module/_03984_ ),
    .B(net429),
    .Y(\reg_module/_03985_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11275_  (.A(\reg_module/_03676_ ),
    .B(\reg_module/gprf[434] ),
    .Y(\reg_module/_03986_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11276_  (.A(\reg_module/gprf[402] ),
    .B(net602),
    .Y(\reg_module/_03987_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11277_  (.A(\reg_module/_03986_ ),
    .B(net490),
    .C(\reg_module/_03987_ ),
    .Y(\reg_module/_03988_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11278_  (.A(\reg_module/_03833_ ),
    .B(\reg_module/gprf[498] ),
    .Y(\reg_module/_03989_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11279_  (.A(\reg_module/gprf[466] ),
    .B(net602),
    .Y(\reg_module/_03990_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11280_  (.A(\reg_module/_03989_ ),
    .B(\reg_module/_03681_ ),
    .C(\reg_module/_03990_ ),
    .Y(\reg_module/_03991_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11281_  (.A(\reg_module/_03988_ ),
    .B(\reg_module/_03991_ ),
    .Y(\reg_module/_03992_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11282_  (.A(\reg_module/_02735_ ),
    .X(\reg_module/_03993_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11283_  (.A(\reg_module/_03992_ ),
    .B(\reg_module/_03993_ ),
    .Y(\reg_module/_03994_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11284_  (.A(\reg_module/_03985_ ),
    .B(\reg_module/_03994_ ),
    .C(\reg_module/_03686_ ),
    .Y(\reg_module/_03995_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11285_  (.A(\reg_module/_03823_ ),
    .B(\reg_module/gprf[50] ),
    .Y(\reg_module/_03996_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11286_  (.A(\reg_module/gprf[18] ),
    .B(net605),
    .Y(\reg_module/_03997_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11287_  (.A(\reg_module/_03996_ ),
    .B(net489),
    .C(\reg_module/_03997_ ),
    .Y(\reg_module/_03998_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11288_  (.A(\reg_module/_03691_ ),
    .B(\reg_module/gprf[114] ),
    .Y(\reg_module/_03999_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11289_  (.A(\reg_module/gprf[82] ),
    .B(net605),
    .Y(\reg_module/_04000_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11290_  (.A(\reg_module/_03999_ ),
    .B(\reg_module/_03844_ ),
    .C(\reg_module/_04000_ ),
    .Y(\reg_module/_04001_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11291_  (.A(\reg_module/_03998_ ),
    .B(\reg_module/_04001_ ),
    .Y(\reg_module/_04002_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11292_  (.A(\reg_module/_04002_ ),
    .B(net429),
    .Y(\reg_module/_04003_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11293_  (.A(\reg_module/_02584_ ),
    .X(\reg_module/_04004_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11294_  (.A(\reg_module/_04004_ ),
    .B(\reg_module/gprf[178] ),
    .Y(\reg_module/_04005_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11295_  (.A(\reg_module/gprf[146] ),
    .B(net593),
    .Y(\reg_module/_04006_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11296_  (.A(\reg_module/_04005_ ),
    .B(net485),
    .C(\reg_module/_04006_ ),
    .Y(\reg_module/_04007_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11297_  (.A(\reg_module/_02491_ ),
    .X(\reg_module/_04008_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11298_  (.A(\reg_module/_04008_ ),
    .B(\reg_module/gprf[242] ),
    .Y(\reg_module/_04009_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11299_  (.A(\reg_module/gprf[210] ),
    .B(net593),
    .Y(\reg_module/_04010_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11300_  (.A(\reg_module/_04009_ ),
    .B(\reg_module/_03853_ ),
    .C(\reg_module/_04010_ ),
    .Y(\reg_module/_04011_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11301_  (.A(\reg_module/_04007_ ),
    .B(\reg_module/_04011_ ),
    .Y(\reg_module/_04012_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11302_  (.A(\reg_module/_02522_ ),
    .X(\reg_module/_04013_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11303_  (.A(\reg_module/_04012_ ),
    .B(\reg_module/_04013_ ),
    .Y(\reg_module/_04014_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11304_  (.A(\reg_module/_04003_ ),
    .B(\reg_module/_04014_ ),
    .C(net400),
    .Y(\reg_module/_04015_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11305_  (.A(\reg_module/_03995_ ),
    .B(\reg_module/_04015_ ),
    .Y(\reg_module/_04016_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11306_  (.A(\reg_module/_04016_ ),
    .B(net384),
    .Y(\reg_module/_04017_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11307_  (.A(\reg_module/_03977_ ),
    .B(\reg_module/_04017_ ),
    .Y(\wRs2Data[18] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11308_  (.A(\reg_module/_03933_ ),
    .B(\reg_module/gprf[819] ),
    .Y(\reg_module/_04018_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11309_  (.A(\reg_module/gprf[787] ),
    .B(net558),
    .Y(\reg_module/_04019_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11310_  (.A(\reg_module/_04018_ ),
    .B(net466),
    .C(\reg_module/_04019_ ),
    .Y(\reg_module/_04020_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11311_  (.A(\reg_module/_03937_ ),
    .B(\reg_module/gprf[883] ),
    .Y(\reg_module/_04021_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11312_  (.A(\reg_module/gprf[851] ),
    .B(net556),
    .Y(\reg_module/_04022_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11313_  (.A(\reg_module/_04021_ ),
    .B(\reg_module/_03939_ ),
    .C(\reg_module/_04022_ ),
    .Y(\reg_module/_04023_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11314_  (.A(\reg_module/_04020_ ),
    .B(\reg_module/_04023_ ),
    .Y(\reg_module/_04024_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11315_  (.A(\reg_module/_04024_ ),
    .B(net417),
    .Y(\reg_module/_04025_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11316_  (.A(\reg_module/_03788_ ),
    .B(\reg_module/gprf[947] ),
    .Y(\reg_module/_04026_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11317_  (.A(\reg_module/gprf[915] ),
    .B(net549),
    .Y(\reg_module/_04027_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11318_  (.A(\reg_module/_04026_ ),
    .B(net461),
    .C(\reg_module/_04027_ ),
    .Y(\reg_module/_04028_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11319_  (.A(\reg_module/_03792_ ),
    .B(\reg_module/gprf[1011] ),
    .Y(\reg_module/_04029_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11320_  (.A(\reg_module/gprf[979] ),
    .B(net548),
    .Y(\reg_module/_04030_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11321_  (.A(\reg_module/_04029_ ),
    .B(\reg_module/_03948_ ),
    .C(\reg_module/_04030_ ),
    .Y(\reg_module/_04031_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11322_  (.A(\reg_module/_04028_ ),
    .B(\reg_module/_04031_ ),
    .Y(\reg_module/_04032_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11323_  (.A(\reg_module/_04032_ ),
    .B(\reg_module/_03642_ ),
    .Y(\reg_module/_04033_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11324_  (.A(\reg_module/_04025_ ),
    .B(\reg_module/_04033_ ),
    .C(\reg_module/_03953_ ),
    .Y(\reg_module/_04034_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11325_  (.A(\reg_module/_03645_ ),
    .B(\reg_module/gprf[691] ),
    .Y(\reg_module/_04035_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11326_  (.A(\reg_module/gprf[659] ),
    .B(net594),
    .Y(\reg_module/_04036_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11327_  (.A(\reg_module/_04035_ ),
    .B(net485),
    .C(\reg_module/_04036_ ),
    .Y(\reg_module/_04037_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11328_  (.A(\reg_module/_03802_ ),
    .B(\reg_module/gprf[755] ),
    .Y(\reg_module/_04038_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11329_  (.A(\reg_module/gprf[723] ),
    .B(net549),
    .Y(\reg_module/_04039_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11330_  (.A(\reg_module/_04038_ ),
    .B(\reg_module/_03650_ ),
    .C(\reg_module/_04039_ ),
    .Y(\reg_module/_04040_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11331_  (.A(\reg_module/_04037_ ),
    .B(\reg_module/_04040_ ),
    .Y(\reg_module/_04041_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11332_  (.A(\reg_module/_04041_ ),
    .B(\reg_module/_03962_ ),
    .Y(\reg_module/_04042_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11333_  (.A(\reg_module/_03964_ ),
    .B(\reg_module/gprf[563] ),
    .Y(\reg_module/_04043_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11334_  (.A(\reg_module/gprf[531] ),
    .B(net555),
    .Y(\reg_module/_04044_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11335_  (.A(\reg_module/_04043_ ),
    .B(net465),
    .C(\reg_module/_04044_ ),
    .Y(\reg_module/_04045_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11336_  (.A(\reg_module/_03658_ ),
    .B(\reg_module/gprf[627] ),
    .Y(\reg_module/_04046_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11337_  (.A(\reg_module/gprf[595] ),
    .B(net555),
    .Y(\reg_module/_04047_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11338_  (.A(\reg_module/_04046_ ),
    .B(\reg_module/_03969_ ),
    .C(\reg_module/_04047_ ),
    .Y(\reg_module/_04048_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11339_  (.A(\reg_module/_04045_ ),
    .B(\reg_module/_04048_ ),
    .Y(\reg_module/_04049_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11340_  (.A(\reg_module/_04049_ ),
    .B(net417),
    .Y(\reg_module/_04050_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11341_  (.A(\reg_module/_04042_ ),
    .B(\reg_module/_04050_ ),
    .C(net392),
    .Y(\reg_module/_04051_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11342_  (.A(\reg_module/_04034_ ),
    .B(\reg_module/_04051_ ),
    .Y(\reg_module/_04052_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11343_  (.A(\reg_module/_04052_ ),
    .B(\reg_module/_03976_ ),
    .Y(\reg_module/_04053_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11344_  (.A(\reg_module/_03819_ ),
    .B(\reg_module/gprf[307] ),
    .Y(\reg_module/_04054_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11345_  (.A(\reg_module/gprf[275] ),
    .B(net557),
    .Y(\reg_module/_04055_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11346_  (.A(\reg_module/_04054_ ),
    .B(net466),
    .C(\reg_module/_04055_ ),
    .Y(\reg_module/_04056_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11347_  (.A(\reg_module/_02897_ ),
    .X(\reg_module/_04057_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11348_  (.A(\reg_module/_04057_ ),
    .B(\reg_module/gprf[371] ),
    .Y(\reg_module/_04058_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11349_  (.A(\reg_module/gprf[339] ),
    .B(net557),
    .Y(\reg_module/_04059_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11350_  (.A(\reg_module/_04058_ ),
    .B(\reg_module/_03825_ ),
    .C(\reg_module/_04059_ ),
    .Y(\reg_module/_04060_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11351_  (.A(\reg_module/_04056_ ),
    .B(\reg_module/_04060_ ),
    .Y(\reg_module/_04061_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11352_  (.A(\reg_module/_04061_ ),
    .B(net417),
    .Y(\reg_module/_04062_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11353_  (.A(\reg_module/_03676_ ),
    .B(\reg_module/gprf[435] ),
    .Y(\reg_module/_04063_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11354_  (.A(\reg_module/gprf[403] ),
    .B(net602),
    .Y(\reg_module/_04064_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11355_  (.A(\reg_module/_04063_ ),
    .B(net490),
    .C(\reg_module/_04064_ ),
    .Y(\reg_module/_04065_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11356_  (.A(\reg_module/_03833_ ),
    .B(\reg_module/gprf[499] ),
    .Y(\reg_module/_04066_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11357_  (.A(\reg_module/gprf[467] ),
    .B(net602),
    .Y(\reg_module/_04067_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11358_  (.A(\reg_module/_04066_ ),
    .B(\reg_module/_03681_ ),
    .C(\reg_module/_04067_ ),
    .Y(\reg_module/_04068_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11359_  (.A(\reg_module/_04065_ ),
    .B(\reg_module/_04068_ ),
    .Y(\reg_module/_04069_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11360_  (.A(\reg_module/_04069_ ),
    .B(\reg_module/_03993_ ),
    .Y(\reg_module/_04070_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11361_  (.A(\reg_module/_04062_ ),
    .B(\reg_module/_04070_ ),
    .C(\reg_module/_03686_ ),
    .Y(\reg_module/_04071_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11362_  (.A(\reg_module/_04057_ ),
    .B(\reg_module/gprf[51] ),
    .Y(\reg_module/_04072_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11363_  (.A(\reg_module/gprf[19] ),
    .B(net605),
    .Y(\reg_module/_04073_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11364_  (.A(\reg_module/_04072_ ),
    .B(net489),
    .C(\reg_module/_04073_ ),
    .Y(\reg_module/_04074_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11365_  (.A(\reg_module/_03691_ ),
    .B(\reg_module/gprf[115] ),
    .Y(\reg_module/_04075_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11366_  (.A(\reg_module/gprf[83] ),
    .B(net605),
    .Y(\reg_module/_04076_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11367_  (.A(\reg_module/_04075_ ),
    .B(\reg_module/_03844_ ),
    .C(\reg_module/_04076_ ),
    .Y(\reg_module/_04077_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11368_  (.A(\reg_module/_04074_ ),
    .B(\reg_module/_04077_ ),
    .Y(\reg_module/_04078_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11369_  (.A(\reg_module/_04078_ ),
    .B(net418),
    .Y(\reg_module/_04079_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11370_  (.A(\reg_module/_04004_ ),
    .B(\reg_module/gprf[179] ),
    .Y(\reg_module/_04080_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11371_  (.A(\reg_module/gprf[147] ),
    .B(net546),
    .Y(\reg_module/_04081_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11372_  (.A(\reg_module/_04080_ ),
    .B(net460),
    .C(\reg_module/_04081_ ),
    .Y(\reg_module/_04082_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11373_  (.A(\reg_module/_04008_ ),
    .B(\reg_module/gprf[243] ),
    .Y(\reg_module/_04083_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11374_  (.A(\reg_module/gprf[211] ),
    .B(net593),
    .Y(\reg_module/_04084_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11375_  (.A(\reg_module/_04083_ ),
    .B(\reg_module/_03853_ ),
    .C(\reg_module/_04084_ ),
    .Y(\reg_module/_04085_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11376_  (.A(\reg_module/_04082_ ),
    .B(\reg_module/_04085_ ),
    .Y(\reg_module/_04086_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11377_  (.A(\reg_module/_04086_ ),
    .B(\reg_module/_04013_ ),
    .Y(\reg_module/_04087_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11378_  (.A(\reg_module/_04079_ ),
    .B(\reg_module/_04087_ ),
    .C(net391),
    .Y(\reg_module/_04088_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11379_  (.A(\reg_module/_04071_ ),
    .B(\reg_module/_04088_ ),
    .Y(\reg_module/_04089_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11380_  (.A(\reg_module/_04089_ ),
    .B(net384),
    .Y(\reg_module/_04090_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11381_  (.A(\reg_module/_04053_ ),
    .B(\reg_module/_04090_ ),
    .Y(\wRs2Data[19] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11382_  (.A(\reg_module/_03933_ ),
    .B(\reg_module/gprf[564] ),
    .Y(\reg_module/_04091_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11383_  (.A(\reg_module/gprf[532] ),
    .B(net555),
    .Y(\reg_module/_04092_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11384_  (.A(\reg_module/_04091_ ),
    .B(net465),
    .C(\reg_module/_04092_ ),
    .Y(\reg_module/_04093_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11385_  (.A(\reg_module/_03937_ ),
    .B(\reg_module/gprf[628] ),
    .Y(\reg_module/_04094_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11386_  (.A(\reg_module/gprf[596] ),
    .B(net556),
    .Y(\reg_module/_04095_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11387_  (.A(\reg_module/_04094_ ),
    .B(\reg_module/_03939_ ),
    .C(\reg_module/_04095_ ),
    .Y(\reg_module/_04096_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11388_  (.A(\reg_module/_04093_ ),
    .B(\reg_module/_04096_ ),
    .Y(\reg_module/_04097_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11389_  (.A(\reg_module/_04097_ ),
    .B(net416),
    .Y(\reg_module/_04098_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11390_  (.A(\reg_module/_03788_ ),
    .B(\reg_module/gprf[692] ),
    .Y(\reg_module/_04099_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11391_  (.A(\reg_module/gprf[660] ),
    .B(net549),
    .Y(\reg_module/_04100_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11392_  (.A(\reg_module/_04099_ ),
    .B(net461),
    .C(\reg_module/_04100_ ),
    .Y(\reg_module/_04101_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11393_  (.A(\reg_module/_03792_ ),
    .B(\reg_module/gprf[756] ),
    .Y(\reg_module/_04102_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11394_  (.A(\reg_module/gprf[724] ),
    .B(net549),
    .Y(\reg_module/_04103_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11395_  (.A(\reg_module/_04102_ ),
    .B(\reg_module/_03948_ ),
    .C(\reg_module/_04103_ ),
    .Y(\reg_module/_04104_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11396_  (.A(\reg_module/_04101_ ),
    .B(\reg_module/_04104_ ),
    .Y(\reg_module/_04105_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11397_  (.A(\reg_module/_02592_ ),
    .X(\reg_module/_04106_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11398_  (.A(\reg_module/_04105_ ),
    .B(\reg_module/_04106_ ),
    .Y(\reg_module/_04107_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11399_  (.A(\reg_module/_04098_ ),
    .B(\reg_module/_04107_ ),
    .C(net391),
    .Y(\reg_module/_04108_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11400_  (.A(\reg_module/_02530_ ),
    .X(\reg_module/_04109_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11401_  (.A(\reg_module/_04109_ ),
    .B(\reg_module/gprf[820] ),
    .Y(\reg_module/_04110_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11402_  (.A(\reg_module/gprf[788] ),
    .B(net552),
    .Y(\reg_module/_04111_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11403_  (.A(\reg_module/_04110_ ),
    .B(net465),
    .C(\reg_module/_04111_ ),
    .Y(\reg_module/_04112_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11404_  (.A(\reg_module/_03802_ ),
    .B(\reg_module/gprf[884] ),
    .Y(\reg_module/_04113_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11405_  (.A(\reg_module/_02516_ ),
    .X(\reg_module/_04114_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11406_  (.A(\reg_module/gprf[852] ),
    .B(net555),
    .Y(\reg_module/_04115_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11407_  (.A(\reg_module/_04113_ ),
    .B(\reg_module/_04114_ ),
    .C(\reg_module/_04115_ ),
    .Y(\reg_module/_04116_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11408_  (.A(\reg_module/_04112_ ),
    .B(\reg_module/_04116_ ),
    .Y(\reg_module/_04117_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11409_  (.A(\reg_module/_04117_ ),
    .B(net416),
    .Y(\reg_module/_04118_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11410_  (.A(\reg_module/_03964_ ),
    .B(\reg_module/gprf[948] ),
    .Y(\reg_module/_04119_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11411_  (.A(\reg_module/gprf[916] ),
    .B(net555),
    .Y(\reg_module/_04120_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11412_  (.A(\reg_module/_04119_ ),
    .B(net465),
    .C(\reg_module/_04120_ ),
    .Y(\reg_module/_04121_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11413_  (.A(\reg_module/_02614_ ),
    .X(\reg_module/_04122_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11414_  (.A(\reg_module/_04122_ ),
    .B(\reg_module/gprf[1012] ),
    .Y(\reg_module/_04123_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11415_  (.A(\reg_module/gprf[980] ),
    .B(net551),
    .Y(\reg_module/_04124_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11416_  (.A(\reg_module/_04123_ ),
    .B(\reg_module/_03969_ ),
    .C(\reg_module/_04124_ ),
    .Y(\reg_module/_04125_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11417_  (.A(\reg_module/_04121_ ),
    .B(\reg_module/_04125_ ),
    .Y(\reg_module/_04126_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11418_  (.A(\reg_module/_04126_ ),
    .B(\reg_module/_03663_ ),
    .Y(\reg_module/_04127_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11419_  (.A(\reg_module/_04118_ ),
    .B(\reg_module/_04127_ ),
    .C(\reg_module/_02527_ ),
    .Y(\reg_module/_04128_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11420_  (.A(\reg_module/_04108_ ),
    .B(\reg_module/_04128_ ),
    .Y(\reg_module/_04129_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11421_  (.A(\reg_module/_04129_ ),
    .B(\reg_module/_03976_ ),
    .Y(\reg_module/_04130_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11422_  (.A(\reg_module/_03819_ ),
    .B(\reg_module/gprf[308] ),
    .Y(\reg_module/_04131_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11423_  (.A(\reg_module/gprf[276] ),
    .B(net554),
    .Y(\reg_module/_04132_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11424_  (.A(\reg_module/_04131_ ),
    .B(net464),
    .C(\reg_module/_04132_ ),
    .Y(\reg_module/_04133_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11425_  (.A(\reg_module/_04057_ ),
    .B(\reg_module/gprf[372] ),
    .Y(\reg_module/_04134_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11426_  (.A(\reg_module/gprf[340] ),
    .B(net554),
    .Y(\reg_module/_04135_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11427_  (.A(\reg_module/_04134_ ),
    .B(\reg_module/_03825_ ),
    .C(\reg_module/_04135_ ),
    .Y(\reg_module/_04136_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11428_  (.A(\reg_module/_04133_ ),
    .B(\reg_module/_04136_ ),
    .Y(\reg_module/_04137_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11429_  (.A(\reg_module/_04137_ ),
    .B(net416),
    .Y(\reg_module/_04138_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11430_  (.A(\reg_module/_02545_ ),
    .X(\reg_module/_04139_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11431_  (.A(\reg_module/_04139_ ),
    .B(\reg_module/gprf[436] ),
    .Y(\reg_module/_04140_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11432_  (.A(\reg_module/gprf[404] ),
    .B(net539),
    .Y(\reg_module/_04141_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11433_  (.A(\reg_module/_04140_ ),
    .B(net458),
    .C(\reg_module/_04141_ ),
    .Y(\reg_module/_04142_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11434_  (.A(\reg_module/_03833_ ),
    .B(\reg_module/gprf[500] ),
    .Y(\reg_module/_04143_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11435_  (.A(\reg_module/_02587_ ),
    .X(\reg_module/_04144_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11436_  (.A(\reg_module/gprf[468] ),
    .B(net539),
    .Y(\reg_module/_04145_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11437_  (.A(\reg_module/_04143_ ),
    .B(\reg_module/_04144_ ),
    .C(\reg_module/_04145_ ),
    .Y(\reg_module/_04146_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11438_  (.A(\reg_module/_04142_ ),
    .B(\reg_module/_04146_ ),
    .Y(\reg_module/_04147_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11439_  (.A(\reg_module/_04147_ ),
    .B(\reg_module/_03993_ ),
    .Y(\reg_module/_04148_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11440_  (.A(\reg_module/_02595_ ),
    .X(\reg_module/_04149_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11441_  (.A(\reg_module/_04138_ ),
    .B(\reg_module/_04148_ ),
    .C(\reg_module/_04149_ ),
    .Y(\reg_module/_04150_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11442_  (.A(\reg_module/_04057_ ),
    .B(\reg_module/gprf[52] ),
    .Y(\reg_module/_04151_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11443_  (.A(\reg_module/gprf[20] ),
    .B(net557),
    .Y(\reg_module/_04152_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11444_  (.A(\reg_module/_04151_ ),
    .B(net466),
    .C(\reg_module/_04152_ ),
    .Y(\reg_module/_04153_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_11445_  (.A(\reg_module/_02601_ ),
    .X(\reg_module/_04154_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11446_  (.A(\reg_module/_04154_ ),
    .B(\reg_module/gprf[116] ),
    .Y(\reg_module/_04155_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11447_  (.A(\reg_module/gprf[84] ),
    .B(net557),
    .Y(\reg_module/_04156_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11448_  (.A(\reg_module/_04155_ ),
    .B(\reg_module/_03844_ ),
    .C(\reg_module/_04156_ ),
    .Y(\reg_module/_04157_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11449_  (.A(\reg_module/_04153_ ),
    .B(\reg_module/_04157_ ),
    .Y(\reg_module/_04158_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11450_  (.A(\reg_module/_04158_ ),
    .B(net417),
    .Y(\reg_module/_04159_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11451_  (.A(\reg_module/_04004_ ),
    .B(\reg_module/gprf[180] ),
    .Y(\reg_module/_04160_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11452_  (.A(\reg_module/gprf[148] ),
    .B(net546),
    .Y(\reg_module/_04161_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11453_  (.A(\reg_module/_04160_ ),
    .B(net460),
    .C(\reg_module/_04161_ ),
    .Y(\reg_module/_04162_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11454_  (.A(\reg_module/_04008_ ),
    .B(\reg_module/gprf[244] ),
    .Y(\reg_module/_04163_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11455_  (.A(\reg_module/gprf[212] ),
    .B(net547),
    .Y(\reg_module/_04164_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11456_  (.A(\reg_module/_04163_ ),
    .B(\reg_module/_03853_ ),
    .C(\reg_module/_04164_ ),
    .Y(\reg_module/_04165_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11457_  (.A(\reg_module/_04162_ ),
    .B(\reg_module/_04165_ ),
    .Y(\reg_module/_04166_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11458_  (.A(\reg_module/_04166_ ),
    .B(\reg_module/_04013_ ),
    .Y(\reg_module/_04167_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11459_  (.A(\reg_module/_04159_ ),
    .B(\reg_module/_04167_ ),
    .C(net392),
    .Y(\reg_module/_04168_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11460_  (.A(\reg_module/_04150_ ),
    .B(\reg_module/_04168_ ),
    .Y(\reg_module/_04169_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11461_  (.A(\reg_module/_04169_ ),
    .B(net383),
    .Y(\reg_module/_04170_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11462_  (.A(\reg_module/_04130_ ),
    .B(\reg_module/_04170_ ),
    .Y(\wRs2Data[20] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11463_  (.A(\reg_module/_03933_ ),
    .B(\reg_module/gprf[821] ),
    .Y(\reg_module/_04171_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11464_  (.A(\reg_module/gprf[789] ),
    .B(net552),
    .Y(\reg_module/_04172_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11465_  (.A(\reg_module/_04171_ ),
    .B(net463),
    .C(\reg_module/_04172_ ),
    .Y(\reg_module/_04173_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11466_  (.A(\reg_module/_03937_ ),
    .B(\reg_module/gprf[885] ),
    .Y(\reg_module/_04174_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11467_  (.A(\reg_module/gprf[853] ),
    .B(net552),
    .Y(\reg_module/_04175_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11468_  (.A(\reg_module/_04174_ ),
    .B(\reg_module/_03939_ ),
    .C(\reg_module/_04175_ ),
    .Y(\reg_module/_04176_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11469_  (.A(\reg_module/_04173_ ),
    .B(\reg_module/_04176_ ),
    .Y(\reg_module/_04177_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11470_  (.A(\reg_module/_04177_ ),
    .B(net415),
    .Y(\reg_module/_04178_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11471_  (.A(\reg_module/_03788_ ),
    .B(\reg_module/gprf[949] ),
    .Y(\reg_module/_04179_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11472_  (.A(\reg_module/gprf[917] ),
    .B(net548),
    .Y(\reg_module/_04180_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11473_  (.A(\reg_module/_04179_ ),
    .B(net461),
    .C(\reg_module/_04180_ ),
    .Y(\reg_module/_04181_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11474_  (.A(\reg_module/_03792_ ),
    .B(\reg_module/gprf[1013] ),
    .Y(\reg_module/_04182_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11475_  (.A(\reg_module/gprf[981] ),
    .B(net544),
    .Y(\reg_module/_04183_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11476_  (.A(\reg_module/_04182_ ),
    .B(\reg_module/_03948_ ),
    .C(\reg_module/_04183_ ),
    .Y(\reg_module/_04184_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11477_  (.A(\reg_module/_04181_ ),
    .B(\reg_module/_04184_ ),
    .Y(\reg_module/_04185_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11478_  (.A(\reg_module/_04185_ ),
    .B(\reg_module/_04106_ ),
    .Y(\reg_module/_04186_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11479_  (.A(\reg_module/_04178_ ),
    .B(\reg_module/_04186_ ),
    .C(\reg_module/_03953_ ),
    .Y(\reg_module/_04187_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11480_  (.A(\reg_module/_04109_ ),
    .B(\reg_module/gprf[693] ),
    .Y(\reg_module/_04188_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11481_  (.A(\reg_module/gprf[661] ),
    .B(net548),
    .Y(\reg_module/_04189_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11482_  (.A(\reg_module/_04188_ ),
    .B(net461),
    .C(\reg_module/_04189_ ),
    .Y(\reg_module/_04190_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11483_  (.A(\reg_module/_03802_ ),
    .B(\reg_module/gprf[757] ),
    .Y(\reg_module/_04191_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11484_  (.A(\reg_module/gprf[725] ),
    .B(net548),
    .Y(\reg_module/_04192_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11485_  (.A(\reg_module/_04191_ ),
    .B(\reg_module/_04114_ ),
    .C(\reg_module/_04192_ ),
    .Y(\reg_module/_04193_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11486_  (.A(\reg_module/_04190_ ),
    .B(\reg_module/_04193_ ),
    .Y(\reg_module/_04194_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11487_  (.A(\reg_module/_04194_ ),
    .B(\reg_module/_03962_ ),
    .Y(\reg_module/_04195_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11488_  (.A(\reg_module/_03964_ ),
    .B(\reg_module/gprf[565] ),
    .Y(\reg_module/_04196_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11489_  (.A(\reg_module/gprf[533] ),
    .B(net551),
    .Y(\reg_module/_04197_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11490_  (.A(\reg_module/_04196_ ),
    .B(net463),
    .C(\reg_module/_04197_ ),
    .Y(\reg_module/_04198_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11491_  (.A(\reg_module/_04122_ ),
    .B(\reg_module/gprf[629] ),
    .Y(\reg_module/_04199_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11492_  (.A(\reg_module/gprf[597] ),
    .B(net551),
    .Y(\reg_module/_04200_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11493_  (.A(\reg_module/_04199_ ),
    .B(\reg_module/_03969_ ),
    .C(\reg_module/_04200_ ),
    .Y(\reg_module/_04201_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11494_  (.A(\reg_module/_04198_ ),
    .B(\reg_module/_04201_ ),
    .Y(\reg_module/_04202_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11495_  (.A(\reg_module/_04202_ ),
    .B(net415),
    .Y(\reg_module/_04203_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11496_  (.A(\reg_module/_04195_ ),
    .B(\reg_module/_04203_ ),
    .C(net391),
    .Y(\reg_module/_04204_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11497_  (.A(\reg_module/_04187_ ),
    .B(\reg_module/_04204_ ),
    .Y(\reg_module/_04205_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11498_  (.A(\reg_module/_04205_ ),
    .B(\reg_module/_03976_ ),
    .Y(\reg_module/_04206_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11499_  (.A(\reg_module/_03819_ ),
    .B(\reg_module/gprf[309] ),
    .Y(\reg_module/_04207_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11500_  (.A(\reg_module/gprf[277] ),
    .B(net554),
    .Y(\reg_module/_04208_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11501_  (.A(\reg_module/_04207_ ),
    .B(net464),
    .C(\reg_module/_04208_ ),
    .Y(\reg_module/_04209_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11502_  (.A(\reg_module/_04057_ ),
    .B(\reg_module/gprf[373] ),
    .Y(\reg_module/_04210_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11503_  (.A(\reg_module/gprf[341] ),
    .B(net554),
    .Y(\reg_module/_04211_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11504_  (.A(\reg_module/_04210_ ),
    .B(\reg_module/_03825_ ),
    .C(\reg_module/_04211_ ),
    .Y(\reg_module/_04212_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11505_  (.A(\reg_module/_04209_ ),
    .B(\reg_module/_04212_ ),
    .Y(\reg_module/_04213_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11506_  (.A(\reg_module/_04213_ ),
    .B(net416),
    .Y(\reg_module/_04214_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11507_  (.A(\reg_module/_04139_ ),
    .B(\reg_module/gprf[437] ),
    .Y(\reg_module/_04215_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11508_  (.A(\reg_module/gprf[405] ),
    .B(net539),
    .Y(\reg_module/_04216_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11509_  (.A(\reg_module/_04215_ ),
    .B(net459),
    .C(\reg_module/_04216_ ),
    .Y(\reg_module/_04217_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11510_  (.A(\reg_module/_03833_ ),
    .B(\reg_module/gprf[501] ),
    .Y(\reg_module/_04218_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11511_  (.A(\reg_module/gprf[469] ),
    .B(net539),
    .Y(\reg_module/_04219_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11512_  (.A(\reg_module/_04218_ ),
    .B(\reg_module/_04144_ ),
    .C(\reg_module/_04219_ ),
    .Y(\reg_module/_04220_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11513_  (.A(\reg_module/_04217_ ),
    .B(\reg_module/_04220_ ),
    .Y(\reg_module/_04221_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11514_  (.A(\reg_module/_04221_ ),
    .B(\reg_module/_03993_ ),
    .Y(\reg_module/_04222_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11515_  (.A(\reg_module/_04214_ ),
    .B(\reg_module/_04222_ ),
    .C(\reg_module/_04149_ ),
    .Y(\reg_module/_04223_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11516_  (.A(\reg_module/_04057_ ),
    .B(\reg_module/gprf[53] ),
    .Y(\reg_module/_04224_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11517_  (.A(\reg_module/gprf[21] ),
    .B(net557),
    .Y(\reg_module/_04225_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11518_  (.A(\reg_module/_04224_ ),
    .B(net466),
    .C(\reg_module/_04225_ ),
    .Y(\reg_module/_04226_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11519_  (.A(\reg_module/_04154_ ),
    .B(\reg_module/gprf[117] ),
    .Y(\reg_module/_04227_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11520_  (.A(\reg_module/gprf[85] ),
    .B(net557),
    .Y(\reg_module/_04228_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11521_  (.A(\reg_module/_04227_ ),
    .B(\reg_module/_03844_ ),
    .C(\reg_module/_04228_ ),
    .Y(\reg_module/_04229_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11522_  (.A(\reg_module/_04226_ ),
    .B(\reg_module/_04229_ ),
    .Y(\reg_module/_04230_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11523_  (.A(\reg_module/_04230_ ),
    .B(net418),
    .Y(\reg_module/_04231_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11524_  (.A(\reg_module/_04004_ ),
    .B(\reg_module/gprf[181] ),
    .Y(\reg_module/_04232_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11525_  (.A(\reg_module/gprf[149] ),
    .B(net546),
    .Y(\reg_module/_04233_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11526_  (.A(\reg_module/_04232_ ),
    .B(net460),
    .C(\reg_module/_04233_ ),
    .Y(\reg_module/_04234_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11527_  (.A(\reg_module/_04008_ ),
    .B(\reg_module/gprf[245] ),
    .Y(\reg_module/_04235_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11528_  (.A(\reg_module/gprf[213] ),
    .B(net546),
    .Y(\reg_module/_04236_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11529_  (.A(\reg_module/_04235_ ),
    .B(\reg_module/_03853_ ),
    .C(\reg_module/_04236_ ),
    .Y(\reg_module/_04237_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11530_  (.A(\reg_module/_04234_ ),
    .B(\reg_module/_04237_ ),
    .Y(\reg_module/_04238_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11531_  (.A(\reg_module/_04238_ ),
    .B(\reg_module/_04013_ ),
    .Y(\reg_module/_04239_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11532_  (.A(\reg_module/_04231_ ),
    .B(\reg_module/_04239_ ),
    .C(net391),
    .Y(\reg_module/_04240_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11533_  (.A(\reg_module/_04223_ ),
    .B(\reg_module/_04240_ ),
    .Y(\reg_module/_04241_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11534_  (.A(\reg_module/_04241_ ),
    .B(net383),
    .Y(\reg_module/_04242_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11535_  (.A(\reg_module/_04206_ ),
    .B(\reg_module/_04242_ ),
    .Y(\wRs2Data[21] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11536_  (.A(\reg_module/_03933_ ),
    .B(\reg_module/gprf[822] ),
    .Y(\reg_module/_04243_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11537_  (.A(\reg_module/gprf[790] ),
    .B(net553),
    .Y(\reg_module/_04244_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11538_  (.A(\reg_module/_04243_ ),
    .B(net463),
    .C(\reg_module/_04244_ ),
    .Y(\reg_module/_04245_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11539_  (.A(\reg_module/_03937_ ),
    .B(\reg_module/gprf[886] ),
    .Y(\reg_module/_04246_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11540_  (.A(\reg_module/gprf[854] ),
    .B(net553),
    .Y(\reg_module/_04247_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11541_  (.A(\reg_module/_04246_ ),
    .B(\reg_module/_03939_ ),
    .C(\reg_module/_04247_ ),
    .Y(\reg_module/_04248_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11542_  (.A(\reg_module/_04245_ ),
    .B(\reg_module/_04248_ ),
    .Y(\reg_module/_04249_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11543_  (.A(\reg_module/_04249_ ),
    .B(net415),
    .Y(\reg_module/_04250_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_11544_  (.A(\reg_module/_02570_ ),
    .X(\reg_module/_04251_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11545_  (.A(\reg_module/_04251_ ),
    .B(\reg_module/gprf[950] ),
    .Y(\reg_module/_04252_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11546_  (.A(\reg_module/gprf[918] ),
    .B(net536),
    .Y(\reg_module/_04253_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11547_  (.A(\reg_module/_04252_ ),
    .B(net456),
    .C(\reg_module/_04253_ ),
    .Y(\reg_module/_04254_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11548_  (.A(\reg_module/_02513_ ),
    .X(\reg_module/_04255_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11549_  (.A(\reg_module/_04255_ ),
    .B(\reg_module/gprf[1014] ),
    .Y(\reg_module/_04256_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11550_  (.A(\reg_module/gprf[982] ),
    .B(net536),
    .Y(\reg_module/_04257_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11551_  (.A(\reg_module/_04256_ ),
    .B(\reg_module/_03948_ ),
    .C(\reg_module/_04257_ ),
    .Y(\reg_module/_04258_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11552_  (.A(\reg_module/_04254_ ),
    .B(\reg_module/_04258_ ),
    .Y(\reg_module/_04259_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11553_  (.A(\reg_module/_04259_ ),
    .B(\reg_module/_04106_ ),
    .Y(\reg_module/_04260_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11554_  (.A(\reg_module/_04250_ ),
    .B(\reg_module/_04260_ ),
    .C(\reg_module/_03953_ ),
    .Y(\reg_module/_04261_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11555_  (.A(\reg_module/_04109_ ),
    .B(\reg_module/gprf[694] ),
    .Y(\reg_module/_04262_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11556_  (.A(\reg_module/gprf[662] ),
    .B(net548),
    .Y(\reg_module/_04263_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11557_  (.A(\reg_module/_04262_ ),
    .B(net462),
    .C(\reg_module/_04263_ ),
    .Y(\reg_module/_04264_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11558_  (.A(\reg_module/_02579_ ),
    .X(\reg_module/_04265_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11559_  (.A(\reg_module/_04265_ ),
    .B(\reg_module/gprf[758] ),
    .Y(\reg_module/_04266_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11560_  (.A(\reg_module/gprf[726] ),
    .B(net545),
    .Y(\reg_module/_04267_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11561_  (.A(\reg_module/_04266_ ),
    .B(\reg_module/_04114_ ),
    .C(\reg_module/_04267_ ),
    .Y(\reg_module/_04268_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11562_  (.A(\reg_module/_04264_ ),
    .B(\reg_module/_04268_ ),
    .Y(\reg_module/_04269_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11563_  (.A(\reg_module/_04269_ ),
    .B(\reg_module/_03962_ ),
    .Y(\reg_module/_04270_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11564_  (.A(\reg_module/_03964_ ),
    .B(\reg_module/gprf[566] ),
    .Y(\reg_module/_04271_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11565_  (.A(\reg_module/gprf[534] ),
    .B(net552),
    .Y(\reg_module/_04272_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11566_  (.A(\reg_module/_04271_ ),
    .B(net463),
    .C(\reg_module/_04272_ ),
    .Y(\reg_module/_04273_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11567_  (.A(\reg_module/_04122_ ),
    .B(\reg_module/gprf[630] ),
    .Y(\reg_module/_04274_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11568_  (.A(\reg_module/gprf[598] ),
    .B(net551),
    .Y(\reg_module/_04275_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11569_  (.A(\reg_module/_04274_ ),
    .B(\reg_module/_03969_ ),
    .C(\reg_module/_04275_ ),
    .Y(\reg_module/_04276_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11570_  (.A(\reg_module/_04273_ ),
    .B(\reg_module/_04276_ ),
    .Y(\reg_module/_04277_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11571_  (.A(\reg_module/_04277_ ),
    .B(net415),
    .Y(\reg_module/_04278_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11572_  (.A(\reg_module/_04270_ ),
    .B(\reg_module/_04278_ ),
    .C(net391),
    .Y(\reg_module/_04279_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11573_  (.A(\reg_module/_04261_ ),
    .B(\reg_module/_04279_ ),
    .Y(\reg_module/_04280_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11574_  (.A(\reg_module/_04280_ ),
    .B(\reg_module/_03976_ ),
    .Y(\reg_module/_04281_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11575_  (.A(\reg_module/_02565_ ),
    .X(\reg_module/_04282_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11576_  (.A(\reg_module/_04282_ ),
    .B(\reg_module/gprf[310] ),
    .Y(\reg_module/_04283_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11577_  (.A(\reg_module/gprf[278] ),
    .B(net540),
    .Y(\reg_module/_04284_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11578_  (.A(\reg_module/_04283_ ),
    .B(net458),
    .C(\reg_module/_04284_ ),
    .Y(\reg_module/_04285_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11579_  (.A(\reg_module/_02535_ ),
    .X(\reg_module/_04286_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11580_  (.A(\reg_module/_04286_ ),
    .B(\reg_module/gprf[374] ),
    .Y(\reg_module/_04287_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11581_  (.A(\reg_module/_02538_ ),
    .X(\reg_module/_04288_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11582_  (.A(\reg_module/gprf[342] ),
    .B(net540),
    .Y(\reg_module/_04289_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11583_  (.A(\reg_module/_04287_ ),
    .B(\reg_module/_04288_ ),
    .C(\reg_module/_04289_ ),
    .Y(\reg_module/_04290_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11584_  (.A(\reg_module/_04285_ ),
    .B(\reg_module/_04290_ ),
    .Y(\reg_module/_04291_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11585_  (.A(\reg_module/_04291_ ),
    .B(net414),
    .Y(\reg_module/_04292_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11586_  (.A(\reg_module/_04139_ ),
    .B(\reg_module/gprf[438] ),
    .Y(\reg_module/_04293_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11587_  (.A(\reg_module/gprf[406] ),
    .B(net539),
    .Y(\reg_module/_04294_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11588_  (.A(\reg_module/_04293_ ),
    .B(net458),
    .C(\reg_module/_04294_ ),
    .Y(\reg_module/_04295_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11589_  (.A(\reg_module/_02550_ ),
    .X(\reg_module/_04296_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11590_  (.A(\reg_module/_04296_ ),
    .B(\reg_module/gprf[502] ),
    .Y(\reg_module/_04297_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11591_  (.A(\reg_module/gprf[470] ),
    .B(net541),
    .Y(\reg_module/_04298_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11592_  (.A(\reg_module/_04297_ ),
    .B(\reg_module/_04144_ ),
    .C(\reg_module/_04298_ ),
    .Y(\reg_module/_04299_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11593_  (.A(\reg_module/_04295_ ),
    .B(\reg_module/_04299_ ),
    .Y(\reg_module/_04300_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11594_  (.A(\reg_module/_04300_ ),
    .B(\reg_module/_03993_ ),
    .Y(\reg_module/_04301_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11595_  (.A(\reg_module/_04292_ ),
    .B(\reg_module/_04301_ ),
    .C(\reg_module/_04149_ ),
    .Y(\reg_module/_04302_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11596_  (.A(\reg_module/_04286_ ),
    .B(\reg_module/gprf[54] ),
    .Y(\reg_module/_04303_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11597_  (.A(\reg_module/gprf[22] ),
    .B(net539),
    .Y(\reg_module/_04304_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11598_  (.A(\reg_module/_04303_ ),
    .B(net459),
    .C(\reg_module/_04304_ ),
    .Y(\reg_module/_04305_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11599_  (.A(\reg_module/_04154_ ),
    .B(\reg_module/gprf[118] ),
    .Y(\reg_module/_04306_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11600_  (.A(\reg_module/_02604_ ),
    .X(\reg_module/_04307_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11601_  (.A(\reg_module/gprf[86] ),
    .B(net540),
    .Y(\reg_module/_04308_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11602_  (.A(\reg_module/_04306_ ),
    .B(\reg_module/_04307_ ),
    .C(\reg_module/_04308_ ),
    .Y(\reg_module/_04309_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11603_  (.A(\reg_module/_04305_ ),
    .B(\reg_module/_04309_ ),
    .Y(\reg_module/_04310_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11604_  (.A(\reg_module/_04310_ ),
    .B(net414),
    .Y(\reg_module/_04311_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11605_  (.A(\reg_module/_04004_ ),
    .B(\reg_module/gprf[182] ),
    .Y(\reg_module/_04312_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11606_  (.A(\reg_module/gprf[150] ),
    .B(net546),
    .Y(\reg_module/_04313_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11607_  (.A(\reg_module/_04312_ ),
    .B(net460),
    .C(\reg_module/_04313_ ),
    .Y(\reg_module/_04314_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11608_  (.A(\reg_module/_04008_ ),
    .B(\reg_module/gprf[246] ),
    .Y(\reg_module/_04315_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_11609_  (.A(\reg_module/_02502_ ),
    .X(\reg_module/_04316_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11610_  (.A(\reg_module/gprf[214] ),
    .B(net547),
    .Y(\reg_module/_04317_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11611_  (.A(\reg_module/_04315_ ),
    .B(\reg_module/_04316_ ),
    .C(\reg_module/_04317_ ),
    .Y(\reg_module/_04318_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11612_  (.A(\reg_module/_04314_ ),
    .B(\reg_module/_04318_ ),
    .Y(\reg_module/_04319_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_11613_  (.A(\reg_module/_04319_ ),
    .B(\reg_module/_04013_ ),
    .Y(\reg_module/_04320_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11614_  (.A(\reg_module/_04311_ ),
    .B(\reg_module/_04320_ ),
    .C(net394),
    .Y(\reg_module/_04321_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11615_  (.A(\reg_module/_04302_ ),
    .B(\reg_module/_04321_ ),
    .Y(\reg_module/_04322_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11616_  (.A(\reg_module/_04322_ ),
    .B(net383),
    .Y(\reg_module/_04323_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11617_  (.A(\reg_module/_04281_ ),
    .B(\reg_module/_04323_ ),
    .Y(\wRs2Data[22] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11618_  (.A(\reg_module/_03933_ ),
    .B(\reg_module/gprf[567] ),
    .Y(\reg_module/_04324_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11619_  (.A(\reg_module/gprf[535] ),
    .B(net551),
    .Y(\reg_module/_04325_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11620_  (.A(\reg_module/_04324_ ),
    .B(net463),
    .C(\reg_module/_04325_ ),
    .Y(\reg_module/_04326_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11621_  (.A(\reg_module/_03937_ ),
    .B(\reg_module/gprf[631] ),
    .Y(\reg_module/_04327_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11622_  (.A(\reg_module/gprf[599] ),
    .B(net552),
    .Y(\reg_module/_04328_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11623_  (.A(\reg_module/_04327_ ),
    .B(\reg_module/_03939_ ),
    .C(\reg_module/_04328_ ),
    .Y(\reg_module/_04329_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11624_  (.A(\reg_module/_04326_ ),
    .B(\reg_module/_04329_ ),
    .Y(\reg_module/_04330_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11625_  (.A(\reg_module/_04330_ ),
    .B(net415),
    .Y(\reg_module/_04331_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11626_  (.A(\reg_module/_04251_ ),
    .B(\reg_module/gprf[695] ),
    .Y(\reg_module/_04332_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11627_  (.A(\reg_module/gprf[663] ),
    .B(net545),
    .Y(\reg_module/_04333_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11628_  (.A(\reg_module/_04332_ ),
    .B(net462),
    .C(\reg_module/_04333_ ),
    .Y(\reg_module/_04334_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11629_  (.A(\reg_module/_04255_ ),
    .B(\reg_module/gprf[759] ),
    .Y(\reg_module/_04335_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11630_  (.A(\reg_module/gprf[727] ),
    .B(net544),
    .Y(\reg_module/_04336_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11631_  (.A(\reg_module/_04335_ ),
    .B(\reg_module/_03948_ ),
    .C(\reg_module/_04336_ ),
    .Y(\reg_module/_04337_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11632_  (.A(\reg_module/_04334_ ),
    .B(\reg_module/_04337_ ),
    .Y(\reg_module/_04338_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11633_  (.A(\reg_module/_04338_ ),
    .B(\reg_module/_04106_ ),
    .Y(\reg_module/_04339_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11634_  (.A(\reg_module/_04331_ ),
    .B(\reg_module/_04339_ ),
    .C(net391),
    .Y(\reg_module/_04340_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11635_  (.A(\reg_module/_04109_ ),
    .B(\reg_module/gprf[823] ),
    .Y(\reg_module/_04341_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11636_  (.A(\reg_module/gprf[791] ),
    .B(net553),
    .Y(\reg_module/_04342_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11637_  (.A(\reg_module/_04341_ ),
    .B(net464),
    .C(\reg_module/_04342_ ),
    .Y(\reg_module/_04343_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11638_  (.A(\reg_module/_04265_ ),
    .B(\reg_module/gprf[887] ),
    .Y(\reg_module/_04344_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11639_  (.A(\reg_module/gprf[855] ),
    .B(net544),
    .Y(\reg_module/_04345_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11640_  (.A(\reg_module/_04344_ ),
    .B(\reg_module/_04114_ ),
    .C(\reg_module/_04345_ ),
    .Y(\reg_module/_04346_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11641_  (.A(\reg_module/_04343_ ),
    .B(\reg_module/_04346_ ),
    .Y(\reg_module/_04347_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11642_  (.A(\reg_module/_04347_ ),
    .B(net415),
    .Y(\reg_module/_04348_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11643_  (.A(\reg_module/_03964_ ),
    .B(\reg_module/gprf[951] ),
    .Y(\reg_module/_04349_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11644_  (.A(\reg_module/gprf[919] ),
    .B(net551),
    .Y(\reg_module/_04350_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11645_  (.A(\reg_module/_04349_ ),
    .B(net463),
    .C(\reg_module/_04350_ ),
    .Y(\reg_module/_04351_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11646_  (.A(\reg_module/_04122_ ),
    .B(\reg_module/gprf[1015] ),
    .Y(\reg_module/_04352_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11647_  (.A(\reg_module/gprf[983] ),
    .B(net544),
    .Y(\reg_module/_04353_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11648_  (.A(\reg_module/_04352_ ),
    .B(\reg_module/_03969_ ),
    .C(\reg_module/_04353_ ),
    .Y(\reg_module/_04354_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11649_  (.A(\reg_module/_04351_ ),
    .B(\reg_module/_04354_ ),
    .Y(\reg_module/_04355_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11650_  (.A(\reg_module/_04355_ ),
    .B(\reg_module/_03663_ ),
    .Y(\reg_module/_04356_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11651_  (.A(\reg_module/_04348_ ),
    .B(\reg_module/_04356_ ),
    .C(\reg_module/_02527_ ),
    .Y(\reg_module/_04357_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11652_  (.A(\reg_module/_04340_ ),
    .B(\reg_module/_04357_ ),
    .Y(\reg_module/_04358_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11653_  (.A(\reg_module/_04358_ ),
    .B(\reg_module/_03976_ ),
    .Y(\reg_module/_04359_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11654_  (.A(\reg_module/_04282_ ),
    .B(\reg_module/gprf[311] ),
    .Y(\reg_module/_04360_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11655_  (.A(\reg_module/gprf[279] ),
    .B(net540),
    .Y(\reg_module/_04361_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11656_  (.A(\reg_module/_04360_ ),
    .B(net458),
    .C(\reg_module/_04361_ ),
    .Y(\reg_module/_04362_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11657_  (.A(\reg_module/_04286_ ),
    .B(\reg_module/gprf[375] ),
    .Y(\reg_module/_04363_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11658_  (.A(\reg_module/gprf[343] ),
    .B(net540),
    .Y(\reg_module/_04364_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11659_  (.A(\reg_module/_04363_ ),
    .B(\reg_module/_04288_ ),
    .C(\reg_module/_04364_ ),
    .Y(\reg_module/_04365_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11660_  (.A(\reg_module/_04362_ ),
    .B(\reg_module/_04365_ ),
    .Y(\reg_module/_04366_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11661_  (.A(\reg_module/_04366_ ),
    .B(net414),
    .Y(\reg_module/_04367_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11662_  (.A(\reg_module/_04139_ ),
    .B(\reg_module/gprf[439] ),
    .Y(\reg_module/_04368_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11663_  (.A(\reg_module/gprf[407] ),
    .B(net541),
    .Y(\reg_module/_04369_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11664_  (.A(\reg_module/_04368_ ),
    .B(net458),
    .C(\reg_module/_04369_ ),
    .Y(\reg_module/_04370_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11665_  (.A(\reg_module/_04296_ ),
    .B(\reg_module/gprf[503] ),
    .Y(\reg_module/_04371_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11666_  (.A(\reg_module/gprf[471] ),
    .B(net541),
    .Y(\reg_module/_04372_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11667_  (.A(\reg_module/_04371_ ),
    .B(\reg_module/_04144_ ),
    .C(\reg_module/_04372_ ),
    .Y(\reg_module/_04373_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11668_  (.A(\reg_module/_04370_ ),
    .B(\reg_module/_04373_ ),
    .Y(\reg_module/_04374_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11669_  (.A(\reg_module/_04374_ ),
    .B(\reg_module/_03993_ ),
    .Y(\reg_module/_04375_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11670_  (.A(\reg_module/_04367_ ),
    .B(\reg_module/_04375_ ),
    .C(\reg_module/_04149_ ),
    .Y(\reg_module/_04376_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11671_  (.A(\reg_module/_04286_ ),
    .B(\reg_module/gprf[55] ),
    .Y(\reg_module/_04377_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11672_  (.A(\reg_module/gprf[23] ),
    .B(net541),
    .Y(\reg_module/_04378_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11673_  (.A(\reg_module/_04377_ ),
    .B(net458),
    .C(\reg_module/_04378_ ),
    .Y(\reg_module/_04379_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11674_  (.A(\reg_module/_04154_ ),
    .B(\reg_module/gprf[119] ),
    .Y(\reg_module/_04380_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11675_  (.A(\reg_module/gprf[87] ),
    .B(net541),
    .Y(\reg_module/_04381_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11676_  (.A(\reg_module/_04380_ ),
    .B(\reg_module/_04307_ ),
    .C(\reg_module/_04381_ ),
    .Y(\reg_module/_04382_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11677_  (.A(\reg_module/_04379_ ),
    .B(\reg_module/_04382_ ),
    .Y(\reg_module/_04383_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11678_  (.A(\reg_module/_04383_ ),
    .B(net414),
    .Y(\reg_module/_04384_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11679_  (.A(\reg_module/_04004_ ),
    .B(\reg_module/gprf[183] ),
    .Y(\reg_module/_04385_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11680_  (.A(\reg_module/gprf[151] ),
    .B(net546),
    .Y(\reg_module/_04386_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11681_  (.A(\reg_module/_04385_ ),
    .B(net460),
    .C(\reg_module/_04386_ ),
    .Y(\reg_module/_04387_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11682_  (.A(\reg_module/_04008_ ),
    .B(\reg_module/gprf[247] ),
    .Y(\reg_module/_04388_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11683_  (.A(\reg_module/gprf[215] ),
    .B(net547),
    .Y(\reg_module/_04389_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11684_  (.A(\reg_module/_04388_ ),
    .B(\reg_module/_04316_ ),
    .C(\reg_module/_04389_ ),
    .Y(\reg_module/_04390_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11685_  (.A(\reg_module/_04387_ ),
    .B(\reg_module/_04390_ ),
    .Y(\reg_module/_04391_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_11686_  (.A(\reg_module/_04391_ ),
    .B(\reg_module/_04013_ ),
    .Y(\reg_module/_04392_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11687_  (.A(\reg_module/_04384_ ),
    .B(\reg_module/_04392_ ),
    .C(net394),
    .Y(\reg_module/_04393_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11688_  (.A(\reg_module/_04376_ ),
    .B(\reg_module/_04393_ ),
    .Y(\reg_module/_04394_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11689_  (.A(\reg_module/_04394_ ),
    .B(net386),
    .Y(\reg_module/_04395_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11690_  (.A(\reg_module/_04359_ ),
    .B(\reg_module/_04395_ ),
    .Y(\wRs2Data[23] ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11691_  (.A(\reg_module/_02565_ ),
    .X(\reg_module/_04396_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11692_  (.A(\reg_module/_04396_ ),
    .B(\reg_module/gprf[824] ),
    .Y(\reg_module/_04397_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11693_  (.A(\reg_module/gprf[792] ),
    .B(net545),
    .Y(\reg_module/_04398_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11694_  (.A(\reg_module/_04397_ ),
    .B(net462),
    .C(\reg_module/_04398_ ),
    .Y(\reg_module/_04399_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11695_  (.A(\reg_module/_02498_ ),
    .X(\reg_module/_04400_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11696_  (.A(\reg_module/_04400_ ),
    .B(\reg_module/gprf[888] ),
    .Y(\reg_module/_04401_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11697_  (.A(\reg_module/_02573_ ),
    .X(\reg_module/_04402_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11698_  (.A(\reg_module/gprf[856] ),
    .B(net545),
    .Y(\reg_module/_04403_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11699_  (.A(\reg_module/_04401_ ),
    .B(\reg_module/_04402_ ),
    .C(\reg_module/_04403_ ),
    .Y(\reg_module/_04404_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11700_  (.A(\reg_module/_04399_ ),
    .B(\reg_module/_04404_ ),
    .Y(\reg_module/_04405_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11701_  (.A(\reg_module/_04405_ ),
    .B(net419),
    .Y(\reg_module/_04406_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11702_  (.A(\reg_module/_04251_ ),
    .B(\reg_module/gprf[952] ),
    .Y(\reg_module/_04407_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11703_  (.A(\reg_module/gprf[920] ),
    .B(net537),
    .Y(\reg_module/_04408_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11704_  (.A(\reg_module/_04407_ ),
    .B(net456),
    .C(\reg_module/_04408_ ),
    .Y(\reg_module/_04409_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11705_  (.A(\reg_module/_04255_ ),
    .B(\reg_module/gprf[1016] ),
    .Y(\reg_module/_04410_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11706_  (.A(\reg_module/_02604_ ),
    .X(\reg_module/_04411_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11707_  (.A(\reg_module/gprf[984] ),
    .B(net538),
    .Y(\reg_module/_04412_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11708_  (.A(\reg_module/_04410_ ),
    .B(\reg_module/_04411_ ),
    .C(\reg_module/_04412_ ),
    .Y(\reg_module/_04413_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11709_  (.A(\reg_module/_04409_ ),
    .B(\reg_module/_04413_ ),
    .Y(\reg_module/_04414_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11710_  (.A(\reg_module/_04414_ ),
    .B(\reg_module/_04106_ ),
    .Y(\reg_module/_04415_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11711_  (.A(\reg_module/_04406_ ),
    .B(\reg_module/_04415_ ),
    .C(\reg_module/_03953_ ),
    .Y(\reg_module/_04416_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11712_  (.A(\reg_module/_04109_ ),
    .B(\reg_module/gprf[696] ),
    .Y(\reg_module/_04417_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11713_  (.A(\reg_module/gprf[664] ),
    .B(net536),
    .Y(\reg_module/_04418_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11714_  (.A(\reg_module/_04417_ ),
    .B(net456),
    .C(\reg_module/_04418_ ),
    .Y(\reg_module/_04419_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11715_  (.A(\reg_module/_04265_ ),
    .B(\reg_module/gprf[760] ),
    .Y(\reg_module/_04420_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11716_  (.A(\reg_module/gprf[728] ),
    .B(net544),
    .Y(\reg_module/_04421_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11717_  (.A(\reg_module/_04420_ ),
    .B(\reg_module/_04114_ ),
    .C(\reg_module/_04421_ ),
    .Y(\reg_module/_04422_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11718_  (.A(\reg_module/_04419_ ),
    .B(\reg_module/_04422_ ),
    .Y(\reg_module/_04423_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11719_  (.A(\reg_module/_04423_ ),
    .B(\reg_module/_03962_ ),
    .Y(\reg_module/_04424_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11720_  (.A(\reg_module/_02513_ ),
    .X(\reg_module/_04425_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11721_  (.A(\reg_module/_04425_ ),
    .B(\reg_module/gprf[568] ),
    .Y(\reg_module/_04426_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11722_  (.A(\reg_module/gprf[536] ),
    .B(net543),
    .Y(\reg_module/_04427_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11723_  (.A(\reg_module/_04426_ ),
    .B(net462),
    .C(\reg_module/_04427_ ),
    .Y(\reg_module/_04428_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11724_  (.A(\reg_module/_04122_ ),
    .B(\reg_module/gprf[632] ),
    .Y(\reg_module/_04429_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11725_  (.A(\reg_module/_02553_ ),
    .X(\reg_module/_04430_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11726_  (.A(\reg_module/gprf[600] ),
    .B(net543),
    .Y(\reg_module/_04431_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11727_  (.A(\reg_module/_04429_ ),
    .B(\reg_module/_04430_ ),
    .C(\reg_module/_04431_ ),
    .Y(\reg_module/_04432_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11728_  (.A(\reg_module/_04428_ ),
    .B(\reg_module/_04432_ ),
    .Y(\reg_module/_04433_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11729_  (.A(\reg_module/_04433_ ),
    .B(net419),
    .Y(\reg_module/_04434_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11730_  (.A(\reg_module/_04424_ ),
    .B(\reg_module/_04434_ ),
    .C(net393),
    .Y(\reg_module/_04435_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11731_  (.A(\reg_module/_04416_ ),
    .B(\reg_module/_04435_ ),
    .Y(\reg_module/_04436_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11732_  (.A(\reg_module/_02561_ ),
    .X(\reg_module/_04437_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11733_  (.A(\reg_module/_04436_ ),
    .B(\reg_module/_04437_ ),
    .Y(\reg_module/_04438_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11734_  (.A(\reg_module/_04282_ ),
    .B(\reg_module/gprf[312] ),
    .Y(\reg_module/_04439_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11735_  (.A(\reg_module/gprf[280] ),
    .B(net536),
    .Y(\reg_module/_04440_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11736_  (.A(\reg_module/_04439_ ),
    .B(net457),
    .C(\reg_module/_04440_ ),
    .Y(\reg_module/_04441_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11737_  (.A(\reg_module/_04286_ ),
    .B(\reg_module/gprf[376] ),
    .Y(\reg_module/_04442_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11738_  (.A(\reg_module/gprf[344] ),
    .B(net536),
    .Y(\reg_module/_04443_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11739_  (.A(\reg_module/_04442_ ),
    .B(\reg_module/_04288_ ),
    .C(\reg_module/_04443_ ),
    .Y(\reg_module/_04444_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11740_  (.A(\reg_module/_04441_ ),
    .B(\reg_module/_04444_ ),
    .Y(\reg_module/_04445_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11741_  (.A(\reg_module/_04445_ ),
    .B(net413),
    .Y(\reg_module/_04446_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11742_  (.A(\reg_module/_04139_ ),
    .B(\reg_module/gprf[440] ),
    .Y(\reg_module/_04447_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11743_  (.A(\reg_module/gprf[408] ),
    .B(net535),
    .Y(\reg_module/_04448_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11744_  (.A(\reg_module/_04447_ ),
    .B(net455),
    .C(\reg_module/_04448_ ),
    .Y(\reg_module/_04449_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11745_  (.A(\reg_module/_04296_ ),
    .B(\reg_module/gprf[504] ),
    .Y(\reg_module/_04450_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11746_  (.A(\reg_module/gprf[472] ),
    .B(net535),
    .Y(\reg_module/_04451_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11747_  (.A(\reg_module/_04450_ ),
    .B(\reg_module/_04144_ ),
    .C(\reg_module/_04451_ ),
    .Y(\reg_module/_04452_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11748_  (.A(\reg_module/_04449_ ),
    .B(\reg_module/_04452_ ),
    .Y(\reg_module/_04453_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11749_  (.A(\reg_module/_02735_ ),
    .X(\reg_module/_04454_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11750_  (.A(\reg_module/_04453_ ),
    .B(\reg_module/_04454_ ),
    .Y(\reg_module/_04455_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11751_  (.A(\reg_module/_04446_ ),
    .B(\reg_module/_04455_ ),
    .C(\reg_module/_04149_ ),
    .Y(\reg_module/_04456_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11752_  (.A(\reg_module/_04286_ ),
    .B(\reg_module/gprf[56] ),
    .Y(\reg_module/_04457_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11753_  (.A(\reg_module/gprf[24] ),
    .B(net538),
    .Y(\reg_module/_04458_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11754_  (.A(\reg_module/_04457_ ),
    .B(net455),
    .C(\reg_module/_04458_ ),
    .Y(\reg_module/_04459_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11755_  (.A(\reg_module/_04154_ ),
    .B(\reg_module/gprf[120] ),
    .Y(\reg_module/_04460_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11756_  (.A(\reg_module/gprf[88] ),
    .B(net538),
    .Y(\reg_module/_04461_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11757_  (.A(\reg_module/_04460_ ),
    .B(\reg_module/_04307_ ),
    .C(\reg_module/_04461_ ),
    .Y(\reg_module/_04462_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11758_  (.A(\reg_module/_04459_ ),
    .B(\reg_module/_04462_ ),
    .Y(\reg_module/_04463_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11759_  (.A(\reg_module/_04463_ ),
    .B(net413),
    .Y(\reg_module/_04464_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11760_  (.A(\reg_module/_02584_ ),
    .X(\reg_module/_04465_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11761_  (.A(\reg_module/_04465_ ),
    .B(\reg_module/gprf[184] ),
    .Y(\reg_module/_04466_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11762_  (.A(\reg_module/gprf[152] ),
    .B(net533),
    .Y(\reg_module/_04467_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11763_  (.A(\reg_module/_04466_ ),
    .B(net454),
    .C(\reg_module/_04467_ ),
    .Y(\reg_module/_04468_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11764_  (.A(\reg_module/_02491_ ),
    .X(\reg_module/_04469_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11765_  (.A(\reg_module/_04469_ ),
    .B(\reg_module/gprf[248] ),
    .Y(\reg_module/_04470_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11766_  (.A(\reg_module/gprf[216] ),
    .B(net533),
    .Y(\reg_module/_04471_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11767_  (.A(\reg_module/_04470_ ),
    .B(\reg_module/_04316_ ),
    .C(\reg_module/_04471_ ),
    .Y(\reg_module/_04472_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11768_  (.A(\reg_module/_04468_ ),
    .B(\reg_module/_04472_ ),
    .Y(\reg_module/_04473_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11769_  (.A(\reg_module/_02522_ ),
    .X(\reg_module/_04474_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11770_  (.A(\reg_module/_04473_ ),
    .B(\reg_module/_04474_ ),
    .Y(\reg_module/_04475_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11771_  (.A(\reg_module/_04464_ ),
    .B(\reg_module/_04475_ ),
    .C(net394),
    .Y(\reg_module/_04476_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11772_  (.A(\reg_module/_04456_ ),
    .B(\reg_module/_04476_ ),
    .Y(\reg_module/_04477_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11773_  (.A(\reg_module/_04477_ ),
    .B(net383),
    .Y(\reg_module/_04478_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11774_  (.A(\reg_module/_04438_ ),
    .B(\reg_module/_04478_ ),
    .Y(\wRs2Data[24] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11775_  (.A(\reg_module/_04396_ ),
    .B(\reg_module/gprf[825] ),
    .Y(\reg_module/_04479_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11776_  (.A(\reg_module/gprf[793] ),
    .B(net547),
    .Y(\reg_module/_04480_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11777_  (.A(\reg_module/_04479_ ),
    .B(net460),
    .C(\reg_module/_04480_ ),
    .Y(\reg_module/_04481_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11778_  (.A(\reg_module/_04400_ ),
    .B(\reg_module/gprf[889] ),
    .Y(\reg_module/_04482_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11779_  (.A(\reg_module/gprf[857] ),
    .B(net547),
    .Y(\reg_module/_04483_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11780_  (.A(\reg_module/_04482_ ),
    .B(\reg_module/_04402_ ),
    .C(\reg_module/_04483_ ),
    .Y(\reg_module/_04484_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11781_  (.A(\reg_module/_04481_ ),
    .B(\reg_module/_04484_ ),
    .Y(\reg_module/_04485_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11782_  (.A(\reg_module/_04485_ ),
    .B(net419),
    .Y(\reg_module/_04486_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11783_  (.A(\reg_module/_04251_ ),
    .B(\reg_module/gprf[953] ),
    .Y(\reg_module/_04487_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11784_  (.A(\reg_module/gprf[921] ),
    .B(net537),
    .Y(\reg_module/_04488_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11785_  (.A(\reg_module/_04487_ ),
    .B(net456),
    .C(\reg_module/_04488_ ),
    .Y(\reg_module/_04489_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11786_  (.A(\reg_module/_04255_ ),
    .B(\reg_module/gprf[1017] ),
    .Y(\reg_module/_04490_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11787_  (.A(\reg_module/gprf[985] ),
    .B(net537),
    .Y(\reg_module/_04491_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11788_  (.A(\reg_module/_04490_ ),
    .B(\reg_module/_04411_ ),
    .C(\reg_module/_04491_ ),
    .Y(\reg_module/_04492_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11789_  (.A(\reg_module/_04489_ ),
    .B(\reg_module/_04492_ ),
    .Y(\reg_module/_04493_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11790_  (.A(\reg_module/_04493_ ),
    .B(\reg_module/_04106_ ),
    .Y(\reg_module/_04494_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11791_  (.A(\reg_module/_04486_ ),
    .B(\reg_module/_04494_ ),
    .C(\reg_module/_03953_ ),
    .Y(\reg_module/_04495_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11792_  (.A(\reg_module/_04109_ ),
    .B(\reg_module/gprf[697] ),
    .Y(\reg_module/_04496_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11793_  (.A(\reg_module/gprf[665] ),
    .B(net536),
    .Y(\reg_module/_04497_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11794_  (.A(\reg_module/_04496_ ),
    .B(net456),
    .C(\reg_module/_04497_ ),
    .Y(\reg_module/_04498_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11795_  (.A(\reg_module/_04265_ ),
    .B(\reg_module/gprf[761] ),
    .Y(\reg_module/_04499_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11796_  (.A(\reg_module/gprf[729] ),
    .B(net544),
    .Y(\reg_module/_04500_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11797_  (.A(\reg_module/_04499_ ),
    .B(\reg_module/_04114_ ),
    .C(\reg_module/_04500_ ),
    .Y(\reg_module/_04501_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11798_  (.A(\reg_module/_04498_ ),
    .B(\reg_module/_04501_ ),
    .Y(\reg_module/_04502_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11799_  (.A(\reg_module/_04502_ ),
    .B(\reg_module/_03962_ ),
    .Y(\reg_module/_04503_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11800_  (.A(\reg_module/_04425_ ),
    .B(\reg_module/gprf[569] ),
    .Y(\reg_module/_04504_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11801_  (.A(\reg_module/gprf[537] ),
    .B(net543),
    .Y(\reg_module/_04505_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11802_  (.A(\reg_module/_04504_ ),
    .B(net462),
    .C(\reg_module/_04505_ ),
    .Y(\reg_module/_04506_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11803_  (.A(\reg_module/_04122_ ),
    .B(\reg_module/gprf[633] ),
    .Y(\reg_module/_04507_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11804_  (.A(\reg_module/gprf[601] ),
    .B(net543),
    .Y(\reg_module/_04508_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11805_  (.A(\reg_module/_04507_ ),
    .B(\reg_module/_04430_ ),
    .C(\reg_module/_04508_ ),
    .Y(\reg_module/_04509_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11806_  (.A(\reg_module/_04506_ ),
    .B(\reg_module/_04509_ ),
    .Y(\reg_module/_04510_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11807_  (.A(\reg_module/_04510_ ),
    .B(net419),
    .Y(\reg_module/_04511_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11808_  (.A(\reg_module/_04503_ ),
    .B(\reg_module/_04511_ ),
    .C(net393),
    .Y(\reg_module/_04512_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11809_  (.A(\reg_module/_04495_ ),
    .B(\reg_module/_04512_ ),
    .Y(\reg_module/_04513_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11810_  (.A(\reg_module/_04513_ ),
    .B(\reg_module/_04437_ ),
    .Y(\reg_module/_04514_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11811_  (.A(\reg_module/_04282_ ),
    .B(\reg_module/gprf[313] ),
    .Y(\reg_module/_04515_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11812_  (.A(\reg_module/gprf[281] ),
    .B(net537),
    .Y(\reg_module/_04516_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11813_  (.A(\reg_module/_04515_ ),
    .B(net454),
    .C(\reg_module/_04516_ ),
    .Y(\reg_module/_04517_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11814_  (.A(\reg_module/_02535_ ),
    .X(\reg_module/_04518_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11815_  (.A(\reg_module/_04518_ ),
    .B(\reg_module/gprf[377] ),
    .Y(\reg_module/_04519_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11816_  (.A(\reg_module/gprf[345] ),
    .B(net534),
    .Y(\reg_module/_04520_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11817_  (.A(\reg_module/_04519_ ),
    .B(\reg_module/_04288_ ),
    .C(\reg_module/_04520_ ),
    .Y(\reg_module/_04521_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11818_  (.A(\reg_module/_04517_ ),
    .B(\reg_module/_04521_ ),
    .Y(\reg_module/_04522_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11819_  (.A(\reg_module/_04522_ ),
    .B(net413),
    .Y(\reg_module/_04523_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11820_  (.A(\reg_module/_04139_ ),
    .B(\reg_module/gprf[441] ),
    .Y(\reg_module/_04524_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11821_  (.A(\reg_module/gprf[409] ),
    .B(net535),
    .Y(\reg_module/_04525_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11822_  (.A(\reg_module/_04524_ ),
    .B(net455),
    .C(\reg_module/_04525_ ),
    .Y(\reg_module/_04526_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11823_  (.A(\reg_module/_04296_ ),
    .B(\reg_module/gprf[505] ),
    .Y(\reg_module/_04527_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11824_  (.A(\reg_module/gprf[473] ),
    .B(net535),
    .Y(\reg_module/_04528_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11825_  (.A(\reg_module/_04527_ ),
    .B(\reg_module/_04144_ ),
    .C(\reg_module/_04528_ ),
    .Y(\reg_module/_04529_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11826_  (.A(\reg_module/_04526_ ),
    .B(\reg_module/_04529_ ),
    .Y(\reg_module/_04530_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11827_  (.A(\reg_module/_04530_ ),
    .B(\reg_module/_04454_ ),
    .Y(\reg_module/_04531_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11828_  (.A(\reg_module/_04523_ ),
    .B(\reg_module/_04531_ ),
    .C(\reg_module/_04149_ ),
    .Y(\reg_module/_04532_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11829_  (.A(\reg_module/_04518_ ),
    .B(\reg_module/gprf[57] ),
    .Y(\reg_module/_04533_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11830_  (.A(\reg_module/gprf[25] ),
    .B(net533),
    .Y(\reg_module/_04534_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11831_  (.A(\reg_module/_04533_ ),
    .B(net454),
    .C(\reg_module/_04534_ ),
    .Y(\reg_module/_04535_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11832_  (.A(\reg_module/_04154_ ),
    .B(\reg_module/gprf[121] ),
    .Y(\reg_module/_04536_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11833_  (.A(\reg_module/gprf[89] ),
    .B(net534),
    .Y(\reg_module/_04537_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11834_  (.A(\reg_module/_04536_ ),
    .B(\reg_module/_04307_ ),
    .C(\reg_module/_04537_ ),
    .Y(\reg_module/_04538_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11835_  (.A(\reg_module/_04535_ ),
    .B(\reg_module/_04538_ ),
    .Y(\reg_module/_04539_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11836_  (.A(\reg_module/_04539_ ),
    .B(net413),
    .Y(\reg_module/_04540_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11837_  (.A(\reg_module/_04465_ ),
    .B(\reg_module/gprf[185] ),
    .Y(\reg_module/_04541_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11838_  (.A(\reg_module/gprf[153] ),
    .B(net533),
    .Y(\reg_module/_04542_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11839_  (.A(\reg_module/_04541_ ),
    .B(net454),
    .C(\reg_module/_04542_ ),
    .Y(\reg_module/_04543_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11840_  (.A(\reg_module/_04469_ ),
    .B(\reg_module/gprf[249] ),
    .Y(\reg_module/_04544_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11841_  (.A(\reg_module/gprf[217] ),
    .B(net533),
    .Y(\reg_module/_04545_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11842_  (.A(\reg_module/_04544_ ),
    .B(\reg_module/_04316_ ),
    .C(\reg_module/_04545_ ),
    .Y(\reg_module/_04546_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11843_  (.A(\reg_module/_04543_ ),
    .B(\reg_module/_04546_ ),
    .Y(\reg_module/_04547_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11844_  (.A(\reg_module/_04547_ ),
    .B(\reg_module/_04474_ ),
    .Y(\reg_module/_04548_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11845_  (.A(\reg_module/_04540_ ),
    .B(\reg_module/_04548_ ),
    .C(net394),
    .Y(\reg_module/_04549_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11846_  (.A(\reg_module/_04532_ ),
    .B(\reg_module/_04549_ ),
    .Y(\reg_module/_04550_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11847_  (.A(\reg_module/_04550_ ),
    .B(net383),
    .Y(\reg_module/_04551_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11848_  (.A(\reg_module/_04514_ ),
    .B(\reg_module/_04551_ ),
    .Y(\wRs2Data[25] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11849_  (.A(\reg_module/_04396_ ),
    .B(\reg_module/gprf[570] ),
    .Y(\reg_module/_04552_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11850_  (.A(\reg_module/gprf[538] ),
    .B(net527),
    .Y(\reg_module/_04553_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11851_  (.A(\reg_module/_04552_ ),
    .B(net452),
    .C(\reg_module/_04553_ ),
    .Y(\reg_module/_04554_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11852_  (.A(\reg_module/_04400_ ),
    .B(\reg_module/gprf[634] ),
    .Y(\reg_module/_04555_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11853_  (.A(\reg_module/gprf[602] ),
    .B(net528),
    .Y(\reg_module/_04556_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11854_  (.A(\reg_module/_04555_ ),
    .B(\reg_module/_04402_ ),
    .C(\reg_module/_04556_ ),
    .Y(\reg_module/_04557_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11855_  (.A(\reg_module/_04554_ ),
    .B(\reg_module/_04557_ ),
    .Y(\reg_module/_04558_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11856_  (.A(\reg_module/_04558_ ),
    .B(net409),
    .Y(\reg_module/_04559_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11857_  (.A(\reg_module/_04251_ ),
    .B(\reg_module/gprf[698] ),
    .Y(\reg_module/_04560_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11858_  (.A(\reg_module/gprf[666] ),
    .B(net537),
    .Y(\reg_module/_04561_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11859_  (.A(\reg_module/_04560_ ),
    .B(net456),
    .C(\reg_module/_04561_ ),
    .Y(\reg_module/_04562_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11860_  (.A(\reg_module/_04255_ ),
    .B(\reg_module/gprf[762] ),
    .Y(\reg_module/_04563_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11861_  (.A(\reg_module/gprf[730] ),
    .B(net537),
    .Y(\reg_module/_04564_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11862_  (.A(\reg_module/_04563_ ),
    .B(\reg_module/_04411_ ),
    .C(\reg_module/_04564_ ),
    .Y(\reg_module/_04565_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11863_  (.A(\reg_module/_04562_ ),
    .B(\reg_module/_04565_ ),
    .Y(\reg_module/_04566_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11864_  (.A(\reg_module/_02592_ ),
    .X(\reg_module/_04567_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11865_  (.A(\reg_module/_04566_ ),
    .B(\reg_module/_04567_ ),
    .Y(\reg_module/_04568_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11866_  (.A(\reg_module/_04559_ ),
    .B(\reg_module/_04568_ ),
    .C(net393),
    .Y(\reg_module/_04569_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_11867_  (.A(\reg_module/_02530_ ),
    .X(\reg_module/_04570_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11868_  (.A(\reg_module/_04570_ ),
    .B(\reg_module/gprf[826] ),
    .Y(\reg_module/_04571_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11869_  (.A(\reg_module/gprf[794] ),
    .B(net531),
    .Y(\reg_module/_04572_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11870_  (.A(\reg_module/_04571_ ),
    .B(net451),
    .C(\reg_module/_04572_ ),
    .Y(\reg_module/_04573_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11871_  (.A(\reg_module/_04265_ ),
    .B(\reg_module/gprf[890] ),
    .Y(\reg_module/_04574_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_11872_  (.A(\reg_module/_02516_ ),
    .X(\reg_module/_04575_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11873_  (.A(\reg_module/gprf[858] ),
    .B(net527),
    .Y(\reg_module/_04576_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11874_  (.A(\reg_module/_04574_ ),
    .B(\reg_module/_04575_ ),
    .C(\reg_module/_04576_ ),
    .Y(\reg_module/_04577_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11875_  (.A(\reg_module/_04573_ ),
    .B(\reg_module/_04577_ ),
    .Y(\reg_module/_04578_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11876_  (.A(\reg_module/_04578_ ),
    .B(net409),
    .Y(\reg_module/_04579_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11877_  (.A(\reg_module/_04425_ ),
    .B(\reg_module/gprf[954] ),
    .Y(\reg_module/_04580_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11878_  (.A(\reg_module/gprf[922] ),
    .B(net543),
    .Y(\reg_module/_04581_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11879_  (.A(\reg_module/_04580_ ),
    .B(net462),
    .C(\reg_module/_04581_ ),
    .Y(\reg_module/_04582_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_11880_  (.A(\reg_module/_02614_ ),
    .X(\reg_module/_04583_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11881_  (.A(\reg_module/_04583_ ),
    .B(\reg_module/gprf[1018] ),
    .Y(\reg_module/_04584_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11882_  (.A(\reg_module/gprf[986] ),
    .B(net543),
    .Y(\reg_module/_04585_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11883_  (.A(\reg_module/_04584_ ),
    .B(\reg_module/_04430_ ),
    .C(\reg_module/_04585_ ),
    .Y(\reg_module/_04586_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11884_  (.A(\reg_module/_04582_ ),
    .B(\reg_module/_04586_ ),
    .Y(\reg_module/_04587_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11885_  (.A(\reg_module/_04587_ ),
    .B(\reg_module/_03663_ ),
    .Y(\reg_module/_04588_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11886_  (.A(\reg_module/_04579_ ),
    .B(\reg_module/_04588_ ),
    .C(\reg_module/_02527_ ),
    .Y(\reg_module/_04589_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11887_  (.A(\reg_module/_04569_ ),
    .B(\reg_module/_04589_ ),
    .Y(\reg_module/_04590_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11888_  (.A(\reg_module/_04590_ ),
    .B(\reg_module/_04437_ ),
    .Y(\reg_module/_04591_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11889_  (.A(\reg_module/_04282_ ),
    .B(\reg_module/gprf[314] ),
    .Y(\reg_module/_04592_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11890_  (.A(\reg_module/gprf[282] ),
    .B(net534),
    .Y(\reg_module/_04593_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11891_  (.A(\reg_module/_04592_ ),
    .B(net454),
    .C(\reg_module/_04593_ ),
    .Y(\reg_module/_04594_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11892_  (.A(\reg_module/_04518_ ),
    .B(\reg_module/gprf[378] ),
    .Y(\reg_module/_04595_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11893_  (.A(\reg_module/gprf[346] ),
    .B(net534),
    .Y(\reg_module/_04596_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11894_  (.A(\reg_module/_04595_ ),
    .B(\reg_module/_04288_ ),
    .C(\reg_module/_04596_ ),
    .Y(\reg_module/_04597_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11895_  (.A(\reg_module/_04594_ ),
    .B(\reg_module/_04597_ ),
    .Y(\reg_module/_04598_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11896_  (.A(\reg_module/_04598_ ),
    .B(net413),
    .Y(\reg_module/_04599_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11897_  (.A(\reg_module/_02545_ ),
    .X(\reg_module/_04600_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11898_  (.A(\reg_module/_04600_ ),
    .B(\reg_module/gprf[442] ),
    .Y(\reg_module/_04601_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11899_  (.A(\reg_module/gprf[410] ),
    .B(net510),
    .Y(\reg_module/_04602_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11900_  (.A(\reg_module/_04601_ ),
    .B(net443),
    .C(\reg_module/_04602_ ),
    .Y(\reg_module/_04603_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11901_  (.A(\reg_module/_04296_ ),
    .B(\reg_module/gprf[506] ),
    .Y(\reg_module/_04604_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_11902_  (.A(\reg_module/_02587_ ),
    .X(\reg_module/_04605_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11903_  (.A(\reg_module/gprf[474] ),
    .B(net510),
    .Y(\reg_module/_04606_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11904_  (.A(\reg_module/_04604_ ),
    .B(\reg_module/_04605_ ),
    .C(\reg_module/_04606_ ),
    .Y(\reg_module/_04607_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11905_  (.A(\reg_module/_04603_ ),
    .B(\reg_module/_04607_ ),
    .Y(\reg_module/_04608_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11906_  (.A(\reg_module/_04608_ ),
    .B(\reg_module/_04454_ ),
    .Y(\reg_module/_04609_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_11907_  (.A(\reg_module/_02526_ ),
    .X(\reg_module/_04610_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11908_  (.A(\reg_module/_04599_ ),
    .B(\reg_module/_04609_ ),
    .C(\reg_module/_04610_ ),
    .Y(\reg_module/_04611_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11909_  (.A(\reg_module/_04518_ ),
    .B(\reg_module/gprf[58] ),
    .Y(\reg_module/_04612_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11910_  (.A(\reg_module/gprf[26] ),
    .B(net533),
    .Y(\reg_module/_04613_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11911_  (.A(\reg_module/_04612_ ),
    .B(net454),
    .C(\reg_module/_04613_ ),
    .Y(\reg_module/_04614_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_11912_  (.A(\reg_module/_02601_ ),
    .X(\reg_module/_04615_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11913_  (.A(\reg_module/_04615_ ),
    .B(\reg_module/gprf[122] ),
    .Y(\reg_module/_04616_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11914_  (.A(\reg_module/gprf[90] ),
    .B(net534),
    .Y(\reg_module/_04617_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11915_  (.A(\reg_module/_04616_ ),
    .B(\reg_module/_04307_ ),
    .C(\reg_module/_04617_ ),
    .Y(\reg_module/_04618_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11916_  (.A(\reg_module/_04614_ ),
    .B(\reg_module/_04618_ ),
    .Y(\reg_module/_04619_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11917_  (.A(\reg_module/_04619_ ),
    .B(net413),
    .Y(\reg_module/_04620_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11918_  (.A(\reg_module/_04465_ ),
    .B(\reg_module/gprf[186] ),
    .Y(\reg_module/_04621_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11919_  (.A(\reg_module/gprf[154] ),
    .B(net511),
    .Y(\reg_module/_04622_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11920_  (.A(\reg_module/_04621_ ),
    .B(net443),
    .C(\reg_module/_04622_ ),
    .Y(\reg_module/_04623_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11921_  (.A(\reg_module/_04469_ ),
    .B(\reg_module/gprf[250] ),
    .Y(\reg_module/_04624_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11922_  (.A(\reg_module/gprf[218] ),
    .B(net511),
    .Y(\reg_module/_04625_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11923_  (.A(\reg_module/_04624_ ),
    .B(\reg_module/_04316_ ),
    .C(\reg_module/_04625_ ),
    .Y(\reg_module/_04626_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11924_  (.A(\reg_module/_04623_ ),
    .B(\reg_module/_04626_ ),
    .Y(\reg_module/_04627_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11925_  (.A(\reg_module/_04627_ ),
    .B(\reg_module/_04474_ ),
    .Y(\reg_module/_04628_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11926_  (.A(\reg_module/_04620_ ),
    .B(\reg_module/_04628_ ),
    .C(net394),
    .Y(\reg_module/_04629_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11927_  (.A(\reg_module/_04611_ ),
    .B(\reg_module/_04629_ ),
    .Y(\reg_module/_04630_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11928_  (.A(\reg_module/_04630_ ),
    .B(net382),
    .Y(\reg_module/_04631_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_11929_  (.A(\reg_module/_04591_ ),
    .B(\reg_module/_04631_ ),
    .Y(\wRs2Data[26] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11930_  (.A(\reg_module/_04396_ ),
    .B(\reg_module/gprf[827] ),
    .Y(\reg_module/_04632_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11931_  (.A(\reg_module/gprf[795] ),
    .B(net531),
    .Y(\reg_module/_04633_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11932_  (.A(\reg_module/_04632_ ),
    .B(net452),
    .C(\reg_module/_04633_ ),
    .Y(\reg_module/_04634_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11933_  (.A(\reg_module/_04400_ ),
    .B(\reg_module/gprf[891] ),
    .Y(\reg_module/_04635_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11934_  (.A(\reg_module/gprf[859] ),
    .B(net531),
    .Y(\reg_module/_04636_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11935_  (.A(\reg_module/_04635_ ),
    .B(\reg_module/_04402_ ),
    .C(\reg_module/_04636_ ),
    .Y(\reg_module/_04637_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11936_  (.A(\reg_module/_04634_ ),
    .B(\reg_module/_04637_ ),
    .Y(\reg_module/_04638_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11937_  (.A(\reg_module/_04638_ ),
    .B(net410),
    .Y(\reg_module/_04639_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11938_  (.A(\reg_module/_04251_ ),
    .B(\reg_module/gprf[955] ),
    .Y(\reg_module/_04640_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11939_  (.A(\reg_module/gprf[923] ),
    .B(net514),
    .Y(\reg_module/_04641_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11940_  (.A(\reg_module/_04640_ ),
    .B(net444),
    .C(\reg_module/_04641_ ),
    .Y(\reg_module/_04642_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11941_  (.A(\reg_module/_04255_ ),
    .B(\reg_module/gprf[1019] ),
    .Y(\reg_module/_04643_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11942_  (.A(\reg_module/gprf[987] ),
    .B(net513),
    .Y(\reg_module/_04644_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11943_  (.A(\reg_module/_04643_ ),
    .B(\reg_module/_04411_ ),
    .C(\reg_module/_04644_ ),
    .Y(\reg_module/_04645_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11944_  (.A(\reg_module/_04642_ ),
    .B(\reg_module/_04645_ ),
    .Y(\reg_module/_04646_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11945_  (.A(\reg_module/_04646_ ),
    .B(\reg_module/_04567_ ),
    .Y(\reg_module/_04647_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11946_  (.A(\reg_module/_04639_ ),
    .B(\reg_module/_04647_ ),
    .C(\reg_module/_02596_ ),
    .Y(\reg_module/_04648_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11947_  (.A(\reg_module/_04570_ ),
    .B(\reg_module/gprf[699] ),
    .Y(\reg_module/_04649_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11948_  (.A(\reg_module/gprf[667] ),
    .B(net527),
    .Y(\reg_module/_04650_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11949_  (.A(\reg_module/_04649_ ),
    .B(net452),
    .C(\reg_module/_04650_ ),
    .Y(\reg_module/_04651_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11950_  (.A(\reg_module/_04265_ ),
    .B(\reg_module/gprf[763] ),
    .Y(\reg_module/_04652_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11951_  (.A(\reg_module/gprf[731] ),
    .B(net527),
    .Y(\reg_module/_04653_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11952_  (.A(\reg_module/_04652_ ),
    .B(\reg_module/_04575_ ),
    .C(\reg_module/_04653_ ),
    .Y(\reg_module/_04654_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11953_  (.A(\reg_module/_04651_ ),
    .B(\reg_module/_04654_ ),
    .Y(\reg_module/_04655_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11954_  (.A(\reg_module/_04655_ ),
    .B(\reg_module/_02524_ ),
    .Y(\reg_module/_04656_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11955_  (.A(\reg_module/_04425_ ),
    .B(\reg_module/gprf[571] ),
    .Y(\reg_module/_04657_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11956_  (.A(\reg_module/gprf[539] ),
    .B(net527),
    .Y(\reg_module/_04658_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11957_  (.A(\reg_module/_04657_ ),
    .B(net450),
    .C(\reg_module/_04658_ ),
    .Y(\reg_module/_04659_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11958_  (.A(\reg_module/_04583_ ),
    .B(\reg_module/gprf[635] ),
    .Y(\reg_module/_04660_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11959_  (.A(\reg_module/gprf[603] ),
    .B(net527),
    .Y(\reg_module/_04661_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11960_  (.A(\reg_module/_04660_ ),
    .B(\reg_module/_04430_ ),
    .C(\reg_module/_04661_ ),
    .Y(\reg_module/_04662_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11961_  (.A(\reg_module/_04659_ ),
    .B(\reg_module/_04662_ ),
    .Y(\reg_module/_04663_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11962_  (.A(\reg_module/_04663_ ),
    .B(net409),
    .Y(\reg_module/_04664_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11963_  (.A(\reg_module/_04656_ ),
    .B(\reg_module/_04664_ ),
    .C(net389),
    .Y(\reg_module/_04665_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11964_  (.A(\reg_module/_04648_ ),
    .B(\reg_module/_04665_ ),
    .Y(\reg_module/_04666_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11965_  (.A(\reg_module/_04666_ ),
    .B(\reg_module/_04437_ ),
    .Y(\reg_module/_04667_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11966_  (.A(\reg_module/_04282_ ),
    .B(\reg_module/gprf[315] ),
    .Y(\reg_module/_04668_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11967_  (.A(\reg_module/gprf[283] ),
    .B(net510),
    .Y(\reg_module/_04669_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11968_  (.A(\reg_module/_04668_ ),
    .B(net455),
    .C(\reg_module/_04669_ ),
    .Y(\reg_module/_04670_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11969_  (.A(\reg_module/_04518_ ),
    .B(\reg_module/gprf[379] ),
    .Y(\reg_module/_04671_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11970_  (.A(\reg_module/gprf[347] ),
    .B(net534),
    .Y(\reg_module/_04672_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11971_  (.A(\reg_module/_04671_ ),
    .B(\reg_module/_04288_ ),
    .C(\reg_module/_04672_ ),
    .Y(\reg_module/_04673_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11972_  (.A(\reg_module/_04670_ ),
    .B(\reg_module/_04673_ ),
    .Y(\reg_module/_04674_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11973_  (.A(\reg_module/_04674_ ),
    .B(net406),
    .Y(\reg_module/_04675_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11974_  (.A(\reg_module/_04600_ ),
    .B(\reg_module/gprf[443] ),
    .Y(\reg_module/_04676_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11975_  (.A(\reg_module/gprf[411] ),
    .B(net510),
    .Y(\reg_module/_04677_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11976_  (.A(\reg_module/_04676_ ),
    .B(net443),
    .C(\reg_module/_04677_ ),
    .Y(\reg_module/_04678_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11977_  (.A(\reg_module/_04296_ ),
    .B(\reg_module/gprf[507] ),
    .Y(\reg_module/_04679_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11978_  (.A(\reg_module/gprf[475] ),
    .B(net510),
    .Y(\reg_module/_04680_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11979_  (.A(\reg_module/_04679_ ),
    .B(\reg_module/_04605_ ),
    .C(\reg_module/_04680_ ),
    .Y(\reg_module/_04681_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11980_  (.A(\reg_module/_04678_ ),
    .B(\reg_module/_04681_ ),
    .Y(\reg_module/_04682_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11981_  (.A(\reg_module/_04682_ ),
    .B(\reg_module/_04454_ ),
    .Y(\reg_module/_04683_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11982_  (.A(\reg_module/_04675_ ),
    .B(\reg_module/_04683_ ),
    .C(\reg_module/_04610_ ),
    .Y(\reg_module/_04684_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11983_  (.A(\reg_module/_04518_ ),
    .B(\reg_module/gprf[59] ),
    .Y(\reg_module/_04685_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11984_  (.A(\reg_module/gprf[27] ),
    .B(net511),
    .Y(\reg_module/_04686_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11985_  (.A(\reg_module/_04685_ ),
    .B(net443),
    .C(\reg_module/_04686_ ),
    .Y(\reg_module/_04687_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11986_  (.A(\reg_module/_04615_ ),
    .B(\reg_module/gprf[123] ),
    .Y(\reg_module/_04688_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11987_  (.A(\reg_module/gprf[91] ),
    .B(net512),
    .Y(\reg_module/_04689_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11988_  (.A(\reg_module/_04688_ ),
    .B(\reg_module/_04307_ ),
    .C(\reg_module/_04689_ ),
    .Y(\reg_module/_04690_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11989_  (.A(\reg_module/_04687_ ),
    .B(\reg_module/_04690_ ),
    .Y(\reg_module/_04691_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11990_  (.A(\reg_module/_04691_ ),
    .B(net406),
    .Y(\reg_module/_04692_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11991_  (.A(\reg_module/_04465_ ),
    .B(\reg_module/gprf[187] ),
    .Y(\reg_module/_04693_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11992_  (.A(\reg_module/gprf[155] ),
    .B(net511),
    .Y(\reg_module/_04694_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11993_  (.A(\reg_module/_04693_ ),
    .B(net443),
    .C(\reg_module/_04694_ ),
    .Y(\reg_module/_04695_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11994_  (.A(\reg_module/_04469_ ),
    .B(\reg_module/gprf[251] ),
    .Y(\reg_module/_04696_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11995_  (.A(\reg_module/gprf[219] ),
    .B(net511),
    .Y(\reg_module/_04697_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11996_  (.A(\reg_module/_04696_ ),
    .B(\reg_module/_04316_ ),
    .C(\reg_module/_04697_ ),
    .Y(\reg_module/_04698_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11997_  (.A(\reg_module/_04695_ ),
    .B(\reg_module/_04698_ ),
    .Y(\reg_module/_04699_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_11998_  (.A(\reg_module/_04699_ ),
    .B(\reg_module/_04474_ ),
    .Y(\reg_module/_04700_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_11999_  (.A(\reg_module/_04692_ ),
    .B(\reg_module/_04700_ ),
    .C(net390),
    .Y(\reg_module/_04701_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12000_  (.A(\reg_module/_04684_ ),
    .B(\reg_module/_04701_ ),
    .Y(\reg_module/_04702_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12001_  (.A(\reg_module/_04702_ ),
    .B(net382),
    .Y(\reg_module/_04703_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_12002_  (.A(\reg_module/_04667_ ),
    .B(\reg_module/_04703_ ),
    .Y(\wRs2Data[27] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12003_  (.A(\reg_module/_04396_ ),
    .B(\reg_module/gprf[828] ),
    .Y(\reg_module/_04704_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12004_  (.A(\reg_module/gprf[796] ),
    .B(net529),
    .Y(\reg_module/_04705_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12005_  (.A(\reg_module/_04704_ ),
    .B(net451),
    .C(\reg_module/_04705_ ),
    .Y(\reg_module/_04706_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12006_  (.A(\reg_module/_04400_ ),
    .B(\reg_module/gprf[892] ),
    .Y(\reg_module/_04707_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12007_  (.A(\reg_module/gprf[860] ),
    .B(net529),
    .Y(\reg_module/_04708_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12008_  (.A(\reg_module/_04707_ ),
    .B(\reg_module/_04402_ ),
    .C(\reg_module/_04708_ ),
    .Y(\reg_module/_04709_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12009_  (.A(\reg_module/_04706_ ),
    .B(\reg_module/_04709_ ),
    .Y(\reg_module/_04710_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12010_  (.A(\reg_module/_04710_ ),
    .B(net410),
    .Y(\reg_module/_04711_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12011_  (.A(\reg_module/_02571_ ),
    .B(\reg_module/gprf[956] ),
    .Y(\reg_module/_04712_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12012_  (.A(\reg_module/gprf[924] ),
    .B(net513),
    .Y(\reg_module/_04713_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12013_  (.A(\reg_module/_04712_ ),
    .B(net444),
    .C(\reg_module/_04713_ ),
    .Y(\reg_module/_04714_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12014_  (.A(\reg_module/_02602_ ),
    .B(\reg_module/gprf[1020] ),
    .Y(\reg_module/_04715_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12015_  (.A(\reg_module/gprf[988] ),
    .B(net513),
    .Y(\reg_module/_04716_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12016_  (.A(\reg_module/_04715_ ),
    .B(\reg_module/_04411_ ),
    .C(\reg_module/_04716_ ),
    .Y(\reg_module/_04717_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12017_  (.A(\reg_module/_04714_ ),
    .B(\reg_module/_04717_ ),
    .Y(\reg_module/_04718_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12018_  (.A(\reg_module/_04718_ ),
    .B(\reg_module/_04567_ ),
    .Y(\reg_module/_04719_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12019_  (.A(\reg_module/_04711_ ),
    .B(\reg_module/_04719_ ),
    .C(\reg_module/_02596_ ),
    .Y(\reg_module/_04720_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12020_  (.A(\reg_module/_04570_ ),
    .B(\reg_module/gprf[700] ),
    .Y(\reg_module/_04721_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12021_  (.A(\reg_module/gprf[668] ),
    .B(net525),
    .Y(\reg_module/_04722_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12022_  (.A(\reg_module/_04721_ ),
    .B(net450),
    .C(\reg_module/_04722_ ),
    .Y(\reg_module/_04723_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12023_  (.A(\reg_module/_02580_ ),
    .B(\reg_module/gprf[764] ),
    .Y(\reg_module/_04724_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12024_  (.A(\reg_module/gprf[732] ),
    .B(net525),
    .Y(\reg_module/_04725_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12025_  (.A(\reg_module/_04724_ ),
    .B(\reg_module/_04575_ ),
    .C(\reg_module/_04725_ ),
    .Y(\reg_module/_04726_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12026_  (.A(\reg_module/_04723_ ),
    .B(\reg_module/_04726_ ),
    .Y(\reg_module/_04727_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12027_  (.A(\reg_module/_04727_ ),
    .B(\reg_module/_02524_ ),
    .Y(\reg_module/_04728_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12028_  (.A(\reg_module/_04425_ ),
    .B(\reg_module/gprf[572] ),
    .Y(\reg_module/_04729_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12029_  (.A(\reg_module/gprf[540] ),
    .B(net525),
    .Y(\reg_module/_04730_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12030_  (.A(\reg_module/_04729_ ),
    .B(net450),
    .C(\reg_module/_04730_ ),
    .Y(\reg_module/_04731_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12031_  (.A(\reg_module/_04583_ ),
    .B(\reg_module/gprf[636] ),
    .Y(\reg_module/_04732_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12032_  (.A(\reg_module/gprf[604] ),
    .B(net525),
    .Y(\reg_module/_04733_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12033_  (.A(\reg_module/_04732_ ),
    .B(\reg_module/_04430_ ),
    .C(\reg_module/_04733_ ),
    .Y(\reg_module/_04734_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12034_  (.A(\reg_module/_04731_ ),
    .B(\reg_module/_04734_ ),
    .Y(\reg_module/_04735_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12035_  (.A(\reg_module/_04735_ ),
    .B(net409),
    .Y(\reg_module/_04736_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12036_  (.A(\reg_module/_04728_ ),
    .B(\reg_module/_04736_ ),
    .C(net389),
    .Y(\reg_module/_04737_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12037_  (.A(\reg_module/_04720_ ),
    .B(\reg_module/_04737_ ),
    .Y(\reg_module/_04738_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12038_  (.A(\reg_module/_04738_ ),
    .B(\reg_module/_04437_ ),
    .Y(\reg_module/_04739_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12039_  (.A(\reg_module/_02531_ ),
    .B(\reg_module/gprf[316] ),
    .Y(\reg_module/_04740_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12040_  (.A(\reg_module/gprf[284] ),
    .B(net513),
    .Y(\reg_module/_04741_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12041_  (.A(\reg_module/_04740_ ),
    .B(net444),
    .C(\reg_module/_04741_ ),
    .Y(\reg_module/_04742_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12042_  (.A(\reg_module/_02535_ ),
    .X(\reg_module/_04743_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12043_  (.A(\reg_module/_04743_ ),
    .B(\reg_module/gprf[380] ),
    .Y(\reg_module/_04744_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12044_  (.A(\reg_module/gprf[348] ),
    .B(net509),
    .Y(\reg_module/_04745_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12045_  (.A(\reg_module/_04744_ ),
    .B(\reg_module/_02539_ ),
    .C(\reg_module/_04745_ ),
    .Y(\reg_module/_04746_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12046_  (.A(\reg_module/_04742_ ),
    .B(\reg_module/_04746_ ),
    .Y(\reg_module/_04747_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12047_  (.A(\reg_module/_04747_ ),
    .B(net405),
    .Y(\reg_module/_04748_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12048_  (.A(\reg_module/_04600_ ),
    .B(\reg_module/gprf[444] ),
    .Y(\reg_module/_04749_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12049_  (.A(\reg_module/gprf[412] ),
    .B(net510),
    .Y(\reg_module/_04750_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12050_  (.A(\reg_module/_04749_ ),
    .B(net442),
    .C(\reg_module/_04750_ ),
    .Y(\reg_module/_04751_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12051_  (.A(\reg_module/_02551_ ),
    .B(\reg_module/gprf[508] ),
    .Y(\reg_module/_04752_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12052_  (.A(\reg_module/gprf[476] ),
    .B(net509),
    .Y(\reg_module/_04753_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12053_  (.A(\reg_module/_04752_ ),
    .B(\reg_module/_04605_ ),
    .C(\reg_module/_04753_ ),
    .Y(\reg_module/_04754_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12054_  (.A(\reg_module/_04751_ ),
    .B(\reg_module/_04754_ ),
    .Y(\reg_module/_04755_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12055_  (.A(\reg_module/_04755_ ),
    .B(\reg_module/_04454_ ),
    .Y(\reg_module/_04756_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12056_  (.A(\reg_module/_04748_ ),
    .B(\reg_module/_04756_ ),
    .C(\reg_module/_04610_ ),
    .Y(\reg_module/_04757_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12057_  (.A(\reg_module/_04743_ ),
    .B(\reg_module/gprf[60] ),
    .Y(\reg_module/_04758_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12058_  (.A(\reg_module/gprf[28] ),
    .B(net508),
    .Y(\reg_module/_04759_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12059_  (.A(\reg_module/_04758_ ),
    .B(net442),
    .C(\reg_module/_04759_ ),
    .Y(\reg_module/_04760_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12060_  (.A(\reg_module/_04615_ ),
    .B(\reg_module/gprf[124] ),
    .Y(\reg_module/_04761_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12061_  (.A(\reg_module/gprf[92] ),
    .B(net509),
    .Y(\reg_module/_04762_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12062_  (.A(\reg_module/_04761_ ),
    .B(\reg_module/_02588_ ),
    .C(\reg_module/_04762_ ),
    .Y(\reg_module/_04763_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12063_  (.A(\reg_module/_04760_ ),
    .B(\reg_module/_04763_ ),
    .Y(\reg_module/_04764_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12064_  (.A(\reg_module/_04764_ ),
    .B(net406),
    .Y(\reg_module/_04765_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12065_  (.A(\reg_module/_04465_ ),
    .B(\reg_module/gprf[188] ),
    .Y(\reg_module/_04766_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12066_  (.A(\reg_module/gprf[156] ),
    .B(net508),
    .Y(\reg_module/_04767_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12067_  (.A(\reg_module/_04766_ ),
    .B(net442),
    .C(\reg_module/_04767_ ),
    .Y(\reg_module/_04768_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12068_  (.A(\reg_module/_04469_ ),
    .B(\reg_module/gprf[252] ),
    .Y(\reg_module/_04769_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12069_  (.A(\reg_module/gprf[220] ),
    .B(net508),
    .Y(\reg_module/_04770_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12070_  (.A(\reg_module/_04769_ ),
    .B(\reg_module/_02503_ ),
    .C(\reg_module/_04770_ ),
    .Y(\reg_module/_04771_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12071_  (.A(\reg_module/_04768_ ),
    .B(\reg_module/_04771_ ),
    .Y(\reg_module/_04772_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12072_  (.A(\reg_module/_04772_ ),
    .B(\reg_module/_04474_ ),
    .Y(\reg_module/_04773_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12073_  (.A(\reg_module/_04765_ ),
    .B(\reg_module/_04773_ ),
    .C(net390),
    .Y(\reg_module/_04774_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12074_  (.A(\reg_module/_04757_ ),
    .B(\reg_module/_04774_ ),
    .Y(\reg_module/_04775_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12075_  (.A(\reg_module/_04775_ ),
    .B(net382),
    .Y(\reg_module/_04776_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_12076_  (.A(\reg_module/_04739_ ),
    .B(\reg_module/_04776_ ),
    .Y(\wRs2Data[28] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12077_  (.A(\reg_module/_04396_ ),
    .B(\reg_module/gprf[573] ),
    .Y(\reg_module/_04777_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12078_  (.A(\reg_module/gprf[541] ),
    .B(net526),
    .Y(\reg_module/_04778_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12079_  (.A(\reg_module/_04777_ ),
    .B(net450),
    .C(\reg_module/_04778_ ),
    .Y(\reg_module/_04779_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12080_  (.A(\reg_module/_04400_ ),
    .B(\reg_module/gprf[637] ),
    .Y(\reg_module/_04780_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12081_  (.A(\reg_module/gprf[605] ),
    .B(net526),
    .Y(\reg_module/_04781_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12082_  (.A(\reg_module/_04780_ ),
    .B(\reg_module/_04402_ ),
    .C(\reg_module/_04781_ ),
    .Y(\reg_module/_04782_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12083_  (.A(\reg_module/_04779_ ),
    .B(\reg_module/_04782_ ),
    .Y(\reg_module/_04783_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12084_  (.A(\reg_module/_04783_ ),
    .B(net409),
    .Y(\reg_module/_04784_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12085_  (.A(\reg_module/_02571_ ),
    .B(\reg_module/gprf[701] ),
    .Y(\reg_module/_04785_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12086_  (.A(\reg_module/gprf[669] ),
    .B(net514),
    .Y(\reg_module/_04786_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12087_  (.A(\reg_module/_04785_ ),
    .B(net444),
    .C(\reg_module/_04786_ ),
    .Y(\reg_module/_04787_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12088_  (.A(\reg_module/_02602_ ),
    .B(\reg_module/gprf[765] ),
    .Y(\reg_module/_04788_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12089_  (.A(\reg_module/gprf[733] ),
    .B(net513),
    .Y(\reg_module/_04789_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12090_  (.A(\reg_module/_04788_ ),
    .B(\reg_module/_04411_ ),
    .C(\reg_module/_04789_ ),
    .Y(\reg_module/_04790_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12091_  (.A(\reg_module/_04787_ ),
    .B(\reg_module/_04790_ ),
    .Y(\reg_module/_04791_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12092_  (.A(\reg_module/_04791_ ),
    .B(\reg_module/_04567_ ),
    .Y(\reg_module/_04792_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12093_  (.A(\reg_module/_04784_ ),
    .B(\reg_module/_04792_ ),
    .C(net389),
    .Y(\reg_module/_04793_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12094_  (.A(\reg_module/_04570_ ),
    .B(\reg_module/gprf[829] ),
    .Y(\reg_module/_04794_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12095_  (.A(\reg_module/gprf[797] ),
    .B(net529),
    .Y(\reg_module/_04795_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12096_  (.A(\reg_module/_04794_ ),
    .B(net451),
    .C(\reg_module/_04795_ ),
    .Y(\reg_module/_04796_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12097_  (.A(\reg_module/_02580_ ),
    .B(\reg_module/gprf[893] ),
    .Y(\reg_module/_04797_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12098_  (.A(\reg_module/gprf[861] ),
    .B(net526),
    .Y(\reg_module/_04798_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12099_  (.A(\reg_module/_04797_ ),
    .B(\reg_module/_04575_ ),
    .C(\reg_module/_04798_ ),
    .Y(\reg_module/_04799_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12100_  (.A(\reg_module/_04796_ ),
    .B(\reg_module/_04799_ ),
    .Y(\reg_module/_04800_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12101_  (.A(\reg_module/_04800_ ),
    .B(net409),
    .Y(\reg_module/_04801_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12102_  (.A(\reg_module/_04425_ ),
    .B(\reg_module/gprf[957] ),
    .Y(\reg_module/_04802_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12103_  (.A(\reg_module/gprf[925] ),
    .B(net525),
    .Y(\reg_module/_04803_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12104_  (.A(\reg_module/_04802_ ),
    .B(net450),
    .C(\reg_module/_04803_ ),
    .Y(\reg_module/_04804_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12105_  (.A(\reg_module/_04583_ ),
    .B(\reg_module/gprf[1021] ),
    .Y(\reg_module/_04805_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12106_  (.A(\reg_module/gprf[989] ),
    .B(net525),
    .Y(\reg_module/_04806_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12107_  (.A(\reg_module/_04805_ ),
    .B(\reg_module/_04430_ ),
    .C(\reg_module/_04806_ ),
    .Y(\reg_module/_04807_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12108_  (.A(\reg_module/_04804_ ),
    .B(\reg_module/_04807_ ),
    .Y(\reg_module/_04808_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12109_  (.A(\reg_module/_04808_ ),
    .B(\reg_module/_03663_ ),
    .Y(\reg_module/_04809_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12110_  (.A(\reg_module/_04801_ ),
    .B(\reg_module/_04809_ ),
    .C(\reg_module/_02527_ ),
    .Y(\reg_module/_04810_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12111_  (.A(\reg_module/_04793_ ),
    .B(\reg_module/_04810_ ),
    .Y(\reg_module/_04811_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12112_  (.A(\reg_module/_04811_ ),
    .B(\reg_module/_04437_ ),
    .Y(\reg_module/_04812_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12113_  (.A(\reg_module/_02531_ ),
    .B(\reg_module/gprf[317] ),
    .Y(\reg_module/_04813_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12114_  (.A(\reg_module/gprf[285] ),
    .B(net513),
    .Y(\reg_module/_04814_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12115_  (.A(\reg_module/_04813_ ),
    .B(net445),
    .C(\reg_module/_04814_ ),
    .Y(\reg_module/_04815_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12116_  (.A(\reg_module/_04743_ ),
    .B(\reg_module/gprf[381] ),
    .Y(\reg_module/_04816_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12117_  (.A(\reg_module/gprf[349] ),
    .B(net512),
    .Y(\reg_module/_04817_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12118_  (.A(\reg_module/_04816_ ),
    .B(\reg_module/_02539_ ),
    .C(\reg_module/_04817_ ),
    .Y(\reg_module/_04818_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12119_  (.A(\reg_module/_04815_ ),
    .B(\reg_module/_04818_ ),
    .Y(\reg_module/_04819_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12120_  (.A(\reg_module/_04819_ ),
    .B(net406),
    .Y(\reg_module/_04820_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12121_  (.A(\reg_module/_04600_ ),
    .B(\reg_module/gprf[445] ),
    .Y(\reg_module/_04821_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12122_  (.A(\reg_module/gprf[413] ),
    .B(net509),
    .Y(\reg_module/_04822_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12123_  (.A(\reg_module/_04821_ ),
    .B(net442),
    .C(\reg_module/_04822_ ),
    .Y(\reg_module/_04823_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12124_  (.A(\reg_module/_02551_ ),
    .B(\reg_module/gprf[509] ),
    .Y(\reg_module/_04824_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12125_  (.A(\reg_module/gprf[477] ),
    .B(net509),
    .Y(\reg_module/_04825_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12126_  (.A(\reg_module/_04824_ ),
    .B(\reg_module/_04605_ ),
    .C(\reg_module/_04825_ ),
    .Y(\reg_module/_04826_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12127_  (.A(\reg_module/_04823_ ),
    .B(\reg_module/_04826_ ),
    .Y(\reg_module/_04827_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12128_  (.A(\reg_module/_04827_ ),
    .B(\reg_module/_04454_ ),
    .Y(\reg_module/_04828_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12129_  (.A(\reg_module/_04820_ ),
    .B(\reg_module/_04828_ ),
    .C(\reg_module/_04610_ ),
    .Y(\reg_module/_04829_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12130_  (.A(\reg_module/_04743_ ),
    .B(\reg_module/gprf[61] ),
    .Y(\reg_module/_04830_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12131_  (.A(\reg_module/gprf[29] ),
    .B(net508),
    .Y(\reg_module/_04831_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12132_  (.A(\reg_module/_04830_ ),
    .B(net442),
    .C(\reg_module/_04831_ ),
    .Y(\reg_module/_04832_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12133_  (.A(\reg_module/_04615_ ),
    .B(\reg_module/gprf[125] ),
    .Y(\reg_module/_04833_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12134_  (.A(\reg_module/gprf[93] ),
    .B(net507),
    .Y(\reg_module/_04834_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12135_  (.A(\reg_module/_04833_ ),
    .B(\reg_module/_02588_ ),
    .C(\reg_module/_04834_ ),
    .Y(\reg_module/_04835_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12136_  (.A(\reg_module/_04832_ ),
    .B(\reg_module/_04835_ ),
    .Y(\reg_module/_04836_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12137_  (.A(\reg_module/_04836_ ),
    .B(net405),
    .Y(\reg_module/_04837_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12138_  (.A(\reg_module/_04465_ ),
    .B(\reg_module/gprf[189] ),
    .Y(\reg_module/_04838_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12139_  (.A(\reg_module/gprf[157] ),
    .B(net508),
    .Y(\reg_module/_04839_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12140_  (.A(\reg_module/_04838_ ),
    .B(net442),
    .C(\reg_module/_04839_ ),
    .Y(\reg_module/_04840_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12141_  (.A(\reg_module/_04469_ ),
    .B(\reg_module/gprf[253] ),
    .Y(\reg_module/_04841_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12142_  (.A(\reg_module/gprf[221] ),
    .B(net508),
    .Y(\reg_module/_04842_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12143_  (.A(\reg_module/_04841_ ),
    .B(\reg_module/_02503_ ),
    .C(\reg_module/_04842_ ),
    .Y(\reg_module/_04843_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12144_  (.A(\reg_module/_04840_ ),
    .B(\reg_module/_04843_ ),
    .Y(\reg_module/_04844_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12145_  (.A(\reg_module/_04844_ ),
    .B(\reg_module/_04474_ ),
    .Y(\reg_module/_04845_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12146_  (.A(\reg_module/_04837_ ),
    .B(\reg_module/_04845_ ),
    .C(net390),
    .Y(\reg_module/_04846_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12147_  (.A(\reg_module/_04829_ ),
    .B(\reg_module/_04846_ ),
    .Y(\reg_module/_04847_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12148_  (.A(\reg_module/_04847_ ),
    .B(net382),
    .Y(\reg_module/_04848_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_12149_  (.A(\reg_module/_04812_ ),
    .B(\reg_module/_04848_ ),
    .Y(\wRs2Data[29] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12150_  (.A(\reg_module/_02566_ ),
    .B(\reg_module/gprf[830] ),
    .Y(\reg_module/_04849_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12151_  (.A(\reg_module/gprf[798] ),
    .B(net526),
    .Y(\reg_module/_04850_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12152_  (.A(\reg_module/_04849_ ),
    .B(net450),
    .C(\reg_module/_04850_ ),
    .Y(\reg_module/_04851_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12153_  (.A(\reg_module/_02509_ ),
    .B(\reg_module/gprf[894] ),
    .Y(\reg_module/_04852_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12154_  (.A(\reg_module/gprf[862] ),
    .B(net524),
    .Y(\reg_module/_04853_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12155_  (.A(\reg_module/_04852_ ),
    .B(\reg_module/_02574_ ),
    .C(\reg_module/_04853_ ),
    .Y(\reg_module/_04854_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12156_  (.A(\reg_module/_04851_ ),
    .B(\reg_module/_04854_ ),
    .Y(\reg_module/_04855_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12157_  (.A(\reg_module/_04855_ ),
    .B(net407),
    .Y(\reg_module/_04856_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12158_  (.A(\reg_module/_02571_ ),
    .B(\reg_module/gprf[958] ),
    .Y(\reg_module/_04857_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12159_  (.A(\reg_module/gprf[926] ),
    .B(net516),
    .Y(\reg_module/_04858_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12160_  (.A(\reg_module/_04857_ ),
    .B(net446),
    .C(\reg_module/_04858_ ),
    .Y(\reg_module/_04859_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12161_  (.A(\reg_module/_02602_ ),
    .B(\reg_module/gprf[1022] ),
    .Y(\reg_module/_04860_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12162_  (.A(\reg_module/gprf[990] ),
    .B(net516),
    .Y(\reg_module/_04861_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12163_  (.A(\reg_module/_04860_ ),
    .B(\reg_module/_02605_ ),
    .C(\reg_module/_04861_ ),
    .Y(\reg_module/_04862_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12164_  (.A(\reg_module/_04859_ ),
    .B(\reg_module/_04862_ ),
    .Y(\reg_module/_04863_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12165_  (.A(\reg_module/_04863_ ),
    .B(\reg_module/_04567_ ),
    .Y(\reg_module/_04864_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12166_  (.A(\reg_module/_04856_ ),
    .B(\reg_module/_04864_ ),
    .C(\reg_module/_02596_ ),
    .Y(\reg_module/_04865_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12167_  (.A(\reg_module/_04570_ ),
    .B(\reg_module/gprf[702] ),
    .Y(\reg_module/_04866_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12168_  (.A(\reg_module/gprf[670] ),
    .B(net516),
    .Y(\reg_module/_04867_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12169_  (.A(\reg_module/_04866_ ),
    .B(net446),
    .C(\reg_module/_04867_ ),
    .Y(\reg_module/_04868_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12170_  (.A(\reg_module/_02580_ ),
    .B(\reg_module/gprf[766] ),
    .Y(\reg_module/_04869_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12171_  (.A(\reg_module/gprf[734] ),
    .B(net516),
    .Y(\reg_module/_04870_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12172_  (.A(\reg_module/_04869_ ),
    .B(\reg_module/_04575_ ),
    .C(\reg_module/_04870_ ),
    .Y(\reg_module/_04871_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12173_  (.A(\reg_module/_04868_ ),
    .B(\reg_module/_04871_ ),
    .Y(\reg_module/_04872_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12174_  (.A(\reg_module/_04872_ ),
    .B(\reg_module/_02524_ ),
    .Y(\reg_module/_04873_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12175_  (.A(\reg_module/_02514_ ),
    .B(\reg_module/gprf[574] ),
    .Y(\reg_module/_04874_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12176_  (.A(\reg_module/gprf[542] ),
    .B(net516),
    .Y(\reg_module/_04875_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12177_  (.A(\reg_module/_04874_ ),
    .B(net446),
    .C(\reg_module/_04875_ ),
    .Y(\reg_module/_04876_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12178_  (.A(\reg_module/_04583_ ),
    .B(\reg_module/gprf[638] ),
    .Y(\reg_module/_04877_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12179_  (.A(\reg_module/gprf[606] ),
    .B(net518),
    .Y(\reg_module/_04878_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12180_  (.A(\reg_module/_04877_ ),
    .B(\reg_module/_02617_ ),
    .C(\reg_module/_04878_ ),
    .Y(\reg_module/_04879_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12181_  (.A(\reg_module/_04876_ ),
    .B(\reg_module/_04879_ ),
    .Y(\reg_module/_04880_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12182_  (.A(\reg_module/_04880_ ),
    .B(net407),
    .Y(\reg_module/_04881_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12183_  (.A(\reg_module/_04873_ ),
    .B(\reg_module/_04881_ ),
    .C(net388),
    .Y(\reg_module/_04882_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12184_  (.A(\reg_module/_04865_ ),
    .B(\reg_module/_04882_ ),
    .Y(\reg_module/_04883_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12185_  (.A(\reg_module/_04883_ ),
    .B(\reg_module/_02562_ ),
    .Y(\reg_module/_04884_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12186_  (.A(\reg_module/_02531_ ),
    .B(\reg_module/gprf[318] ),
    .Y(\reg_module/_04885_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12187_  (.A(\reg_module/gprf[286] ),
    .B(net505),
    .Y(\reg_module/_04886_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12188_  (.A(\reg_module/_04885_ ),
    .B(net441),
    .C(\reg_module/_04886_ ),
    .Y(\reg_module/_04887_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12189_  (.A(\reg_module/_04743_ ),
    .B(\reg_module/gprf[382] ),
    .Y(\reg_module/_04888_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12190_  (.A(\reg_module/gprf[350] ),
    .B(net505),
    .Y(\reg_module/_04889_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12191_  (.A(\reg_module/_04888_ ),
    .B(\reg_module/_02539_ ),
    .C(\reg_module/_04889_ ),
    .Y(\reg_module/_04890_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12192_  (.A(\reg_module/_04887_ ),
    .B(\reg_module/_04890_ ),
    .Y(\reg_module/_04891_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12193_  (.A(\reg_module/_04891_ ),
    .B(net405),
    .Y(\reg_module/_04892_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12194_  (.A(\reg_module/_04600_ ),
    .B(\reg_module/gprf[446] ),
    .Y(\reg_module/_04893_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12195_  (.A(\reg_module/gprf[414] ),
    .B(net507),
    .Y(\reg_module/_04894_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12196_  (.A(\reg_module/_04893_ ),
    .B(net441),
    .C(\reg_module/_04894_ ),
    .Y(\reg_module/_04895_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12197_  (.A(\reg_module/_02551_ ),
    .B(\reg_module/gprf[510] ),
    .Y(\reg_module/_04896_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12198_  (.A(\reg_module/gprf[478] ),
    .B(net507),
    .Y(\reg_module/_04897_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12199_  (.A(\reg_module/_04896_ ),
    .B(\reg_module/_04605_ ),
    .C(\reg_module/_04897_ ),
    .Y(\reg_module/_04898_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12200_  (.A(\reg_module/_04895_ ),
    .B(\reg_module/_04898_ ),
    .Y(\reg_module/_04899_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12201_  (.A(\reg_module/_04899_ ),
    .B(\reg_module/_02736_ ),
    .Y(\reg_module/_04900_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12202_  (.A(\reg_module/_04892_ ),
    .B(\reg_module/_04900_ ),
    .C(\reg_module/_04610_ ),
    .Y(\reg_module/_04901_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12203_  (.A(\reg_module/_04743_ ),
    .B(\reg_module/gprf[62] ),
    .Y(\reg_module/_04902_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12204_  (.A(\reg_module/gprf[30] ),
    .B(net505),
    .Y(\reg_module/_04903_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12205_  (.A(\reg_module/_04902_ ),
    .B(net440),
    .C(\reg_module/_04903_ ),
    .Y(\reg_module/_04904_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12206_  (.A(\reg_module/_04615_ ),
    .B(\reg_module/gprf[126] ),
    .Y(\reg_module/_04905_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12207_  (.A(\reg_module/gprf[94] ),
    .B(net507),
    .Y(\reg_module/_04906_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12208_  (.A(\reg_module/_04905_ ),
    .B(\reg_module/_02588_ ),
    .C(\reg_module/_04906_ ),
    .Y(\reg_module/_04907_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12209_  (.A(\reg_module/_04904_ ),
    .B(\reg_module/_04907_ ),
    .Y(\reg_module/_04908_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12210_  (.A(\reg_module/_04908_ ),
    .B(net405),
    .Y(\reg_module/_04909_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12211_  (.A(\reg_module/_02585_ ),
    .B(\reg_module/gprf[190] ),
    .Y(\reg_module/_04910_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12212_  (.A(\reg_module/gprf[158] ),
    .B(net506),
    .Y(\reg_module/_04911_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12213_  (.A(\reg_module/_04910_ ),
    .B(net440),
    .C(\reg_module/_04911_ ),
    .Y(\reg_module/_04912_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12214_  (.A(\reg_module/_02492_ ),
    .B(\reg_module/gprf[254] ),
    .Y(\reg_module/_04913_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12215_  (.A(\reg_module/gprf[222] ),
    .B(net506),
    .Y(\reg_module/_04914_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12216_  (.A(\reg_module/_04913_ ),
    .B(\reg_module/_02503_ ),
    .C(\reg_module/_04914_ ),
    .Y(\reg_module/_04915_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12217_  (.A(\reg_module/_04912_ ),
    .B(\reg_module/_04915_ ),
    .Y(\reg_module/_04916_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12218_  (.A(\reg_module/_04916_ ),
    .B(\reg_module/_02523_ ),
    .Y(\reg_module/_04917_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12219_  (.A(\reg_module/_04909_ ),
    .B(\reg_module/_04917_ ),
    .C(net390),
    .Y(\reg_module/_04918_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12220_  (.A(\reg_module/_04901_ ),
    .B(\reg_module/_04918_ ),
    .Y(\reg_module/_04919_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12221_  (.A(\reg_module/_04919_ ),
    .B(net382),
    .Y(\reg_module/_04920_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_12222_  (.A(\reg_module/_04884_ ),
    .B(\reg_module/_04920_ ),
    .Y(\wRs2Data[30] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12223_  (.A(\reg_module/_02566_ ),
    .B(\reg_module/gprf[831] ),
    .Y(\reg_module/_04921_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12224_  (.A(\reg_module/gprf[799] ),
    .B(net518),
    .Y(\reg_module/_04922_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12225_  (.A(\reg_module/_04921_ ),
    .B(net449),
    .C(\reg_module/_04922_ ),
    .Y(\reg_module/_04923_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12226_  (.A(\reg_module/_02509_ ),
    .B(\reg_module/gprf[895] ),
    .Y(\reg_module/_04924_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12227_  (.A(\reg_module/gprf[863] ),
    .B(net518),
    .Y(\reg_module/_04925_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12228_  (.A(\reg_module/_04924_ ),
    .B(\reg_module/_02574_ ),
    .C(\reg_module/_04925_ ),
    .Y(\reg_module/_04926_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12229_  (.A(\reg_module/_04923_ ),
    .B(\reg_module/_04926_ ),
    .Y(\reg_module/_04927_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12230_  (.A(\reg_module/_04927_ ),
    .B(net407),
    .Y(\reg_module/_04928_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12231_  (.A(\reg_module/_02571_ ),
    .B(\reg_module/gprf[959] ),
    .Y(\reg_module/_04929_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12232_  (.A(\reg_module/gprf[927] ),
    .B(net517),
    .Y(\reg_module/_04930_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12233_  (.A(\reg_module/_04929_ ),
    .B(net446),
    .C(\reg_module/_04930_ ),
    .Y(\reg_module/_04931_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12234_  (.A(\reg_module/_02602_ ),
    .B(\reg_module/gprf[1023] ),
    .Y(\reg_module/_04932_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12235_  (.A(\reg_module/gprf[991] ),
    .B(net517),
    .Y(\reg_module/_04933_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12236_  (.A(\reg_module/_04932_ ),
    .B(\reg_module/_02605_ ),
    .C(\reg_module/_04933_ ),
    .Y(\reg_module/_04934_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12237_  (.A(\reg_module/_04931_ ),
    .B(\reg_module/_04934_ ),
    .Y(\reg_module/_04935_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12238_  (.A(\reg_module/_04935_ ),
    .B(\reg_module/_04567_ ),
    .Y(\reg_module/_04936_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12239_  (.A(\reg_module/_04928_ ),
    .B(\reg_module/_04936_ ),
    .C(\reg_module/_02596_ ),
    .Y(\reg_module/_04937_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12240_  (.A(\reg_module/_04570_ ),
    .B(\reg_module/gprf[703] ),
    .Y(\reg_module/_04938_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12241_  (.A(\reg_module/gprf[671] ),
    .B(net516),
    .Y(\reg_module/_04939_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12242_  (.A(\reg_module/_04938_ ),
    .B(net446),
    .C(\reg_module/_04939_ ),
    .Y(\reg_module/_04940_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12243_  (.A(\reg_module/_02580_ ),
    .B(\reg_module/gprf[767] ),
    .Y(\reg_module/_04941_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12244_  (.A(\reg_module/gprf[735] ),
    .B(net517),
    .Y(\reg_module/_04942_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12245_  (.A(\reg_module/_04941_ ),
    .B(\reg_module/_04575_ ),
    .C(\reg_module/_04942_ ),
    .Y(\reg_module/_04943_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12246_  (.A(\reg_module/_04940_ ),
    .B(\reg_module/_04943_ ),
    .Y(\reg_module/_04944_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12247_  (.A(\reg_module/_04944_ ),
    .B(\reg_module/_02524_ ),
    .Y(\reg_module/_04945_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12248_  (.A(\reg_module/_02514_ ),
    .B(\reg_module/gprf[575] ),
    .Y(\reg_module/_04946_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12249_  (.A(\reg_module/gprf[543] ),
    .B(net524),
    .Y(\reg_module/_04947_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12250_  (.A(\reg_module/_04946_ ),
    .B(net446),
    .C(\reg_module/_04947_ ),
    .Y(\reg_module/_04948_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12251_  (.A(\reg_module/_04583_ ),
    .B(\reg_module/gprf[639] ),
    .Y(\reg_module/_04949_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12252_  (.A(\reg_module/gprf[607] ),
    .B(net518),
    .Y(\reg_module/_04950_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12253_  (.A(\reg_module/_04949_ ),
    .B(\reg_module/_02617_ ),
    .C(\reg_module/_04950_ ),
    .Y(\reg_module/_04951_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12254_  (.A(\reg_module/_04948_ ),
    .B(\reg_module/_04951_ ),
    .Y(\reg_module/_04952_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12255_  (.A(\reg_module/_04952_ ),
    .B(net407),
    .Y(\reg_module/_04953_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12256_  (.A(\reg_module/_04945_ ),
    .B(\reg_module/_04953_ ),
    .C(net388),
    .Y(\reg_module/_04954_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12257_  (.A(\reg_module/_04937_ ),
    .B(\reg_module/_04954_ ),
    .Y(\reg_module/_04955_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12258_  (.A(\reg_module/_04955_ ),
    .B(\reg_module/_02562_ ),
    .Y(\reg_module/_04956_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12259_  (.A(\reg_module/_02531_ ),
    .B(\reg_module/gprf[319] ),
    .Y(\reg_module/_04957_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12260_  (.A(\reg_module/gprf[287] ),
    .B(net505),
    .Y(\reg_module/_04958_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12261_  (.A(\reg_module/_04957_ ),
    .B(net440),
    .C(\reg_module/_04958_ ),
    .Y(\reg_module/_04959_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12262_  (.A(\reg_module/_02536_ ),
    .B(\reg_module/gprf[383] ),
    .Y(\reg_module/_04960_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12263_  (.A(\reg_module/gprf[351] ),
    .B(net515),
    .Y(\reg_module/_04961_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12264_  (.A(\reg_module/_04960_ ),
    .B(\reg_module/_02539_ ),
    .C(\reg_module/_04961_ ),
    .Y(\reg_module/_04962_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12265_  (.A(\reg_module/_04959_ ),
    .B(\reg_module/_04962_ ),
    .Y(\reg_module/_04963_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12266_  (.A(\reg_module/_04963_ ),
    .B(net405),
    .Y(\reg_module/_04964_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12267_  (.A(\reg_module/_04600_ ),
    .B(\reg_module/gprf[447] ),
    .Y(\reg_module/_04965_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12268_  (.A(\reg_module/gprf[415] ),
    .B(net505),
    .Y(\reg_module/_04966_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12269_  (.A(\reg_module/_04965_ ),
    .B(net440),
    .C(\reg_module/_04966_ ),
    .Y(\reg_module/_04967_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12270_  (.A(\reg_module/_02551_ ),
    .B(\reg_module/gprf[511] ),
    .Y(\reg_module/_04968_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12271_  (.A(\reg_module/gprf[479] ),
    .B(net505),
    .Y(\reg_module/_04969_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12272_  (.A(\reg_module/_04968_ ),
    .B(\reg_module/_04605_ ),
    .C(\reg_module/_04969_ ),
    .Y(\reg_module/_04970_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12273_  (.A(\reg_module/_04967_ ),
    .B(\reg_module/_04970_ ),
    .Y(\reg_module/_04971_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12274_  (.A(\reg_module/_04971_ ),
    .B(\reg_module/_02736_ ),
    .Y(\reg_module/_04972_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12275_  (.A(\reg_module/_04964_ ),
    .B(\reg_module/_04972_ ),
    .C(\reg_module/_04610_ ),
    .Y(\reg_module/_04973_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12276_  (.A(\reg_module/_02536_ ),
    .B(\reg_module/gprf[63] ),
    .Y(\reg_module/_04974_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12277_  (.A(\reg_module/gprf[31] ),
    .B(net506),
    .Y(\reg_module/_04975_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12278_  (.A(\reg_module/_04974_ ),
    .B(net440),
    .C(\reg_module/_04975_ ),
    .Y(\reg_module/_04976_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12279_  (.A(\reg_module/_04615_ ),
    .B(\reg_module/gprf[127] ),
    .Y(\reg_module/_04977_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12280_  (.A(\reg_module/gprf[95] ),
    .B(net507),
    .Y(\reg_module/_04978_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12281_  (.A(\reg_module/_04977_ ),
    .B(\reg_module/_02588_ ),
    .C(\reg_module/_04978_ ),
    .Y(\reg_module/_04979_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12282_  (.A(\reg_module/_04976_ ),
    .B(\reg_module/_04979_ ),
    .Y(\reg_module/_04980_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12283_  (.A(\reg_module/_04980_ ),
    .B(net405),
    .Y(\reg_module/_04981_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12284_  (.A(\reg_module/_02585_ ),
    .B(\reg_module/gprf[191] ),
    .Y(\reg_module/_04982_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12285_  (.A(\reg_module/gprf[159] ),
    .B(net506),
    .Y(\reg_module/_04983_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12286_  (.A(\reg_module/_04982_ ),
    .B(net440),
    .C(\reg_module/_04983_ ),
    .Y(\reg_module/_04984_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12287_  (.A(\reg_module/_02492_ ),
    .B(\reg_module/gprf[255] ),
    .Y(\reg_module/_04985_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12288_  (.A(\reg_module/gprf[223] ),
    .B(net506),
    .Y(\reg_module/_04986_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12289_  (.A(\reg_module/_04985_ ),
    .B(\reg_module/_02503_ ),
    .C(\reg_module/_04986_ ),
    .Y(\reg_module/_04987_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12290_  (.A(\reg_module/_04984_ ),
    .B(\reg_module/_04987_ ),
    .Y(\reg_module/_04988_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12291_  (.A(\reg_module/_04988_ ),
    .B(\reg_module/_02523_ ),
    .Y(\reg_module/_04989_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12292_  (.A(\reg_module/_04981_ ),
    .B(\reg_module/_04989_ ),
    .C(net390),
    .Y(\reg_module/_04990_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12293_  (.A(\reg_module/_04973_ ),
    .B(\reg_module/_04990_ ),
    .Y(\reg_module/_04991_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12294_  (.A(\reg_module/_04991_ ),
    .B(net382),
    .Y(\reg_module/_04992_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_12295_  (.A(\reg_module/_04956_ ),
    .B(\reg_module/_04992_ ),
    .Y(\wRs2Data[31] ));
 sky130_fd_sc_hd__inv_2 \reg_module/_12296_  (.A(net2192),
    .Y(\reg_module/_04993_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_12297_  (.A(net770),
    .B(\reg_module/_04993_ ),
    .Y(\reg_module/_04994_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12298_  (.A(\reg_module/gprf[192] ),
    .B(net770),
    .Y(\reg_module/_04995_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_12299_  (.A(net723),
    .Y(\reg_module/_04996_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_12300_  (.A(\reg_module/_04996_ ),
    .X(\reg_module/_04997_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12301_  (.A(\reg_module/_04997_ ),
    .X(\reg_module/_04998_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12302_  (.A(\reg_module/_04995_ ),
    .B(\reg_module/_04998_ ),
    .Y(\reg_module/_04999_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_12303_  (.A(net822),
    .Y(\reg_module/_05000_ ));
 sky130_fd_sc_hd__buf_1 \reg_module/_12304_  (.A(\reg_module/_05000_ ),
    .X(\reg_module/_05001_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12305_  (.A(\reg_module/_05001_ ),
    .X(\reg_module/_05002_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12306_  (.A(\reg_module/_05002_ ),
    .X(\reg_module/_05003_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12307_  (.A(\reg_module/_05003_ ),
    .B(\reg_module/gprf[160] ),
    .Y(\reg_module/_05004_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12308_  (.A(\reg_module/gprf[128] ),
    .B(net768),
    .Y(\reg_module/_05005_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12309_  (.A(\reg_module/_05004_ ),
    .B(net695),
    .C(\reg_module/_05005_ ),
    .Y(\reg_module/_05006_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_12310_  (.A1(\reg_module/_04994_ ),
    .A2(\reg_module/_04999_ ),
    .B1(\reg_module/_05006_ ),
    .Y(\reg_module/_05007_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_12311_  (.A(net660),
    .Y(\reg_module/_05008_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12312_  (.A(\reg_module/_05008_ ),
    .X(\reg_module/_05009_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12313_  (.A(\reg_module/_05009_ ),
    .X(\reg_module/_05010_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12314_  (.A(\reg_module/_05010_ ),
    .X(\reg_module/_05011_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12315_  (.A(\reg_module/_05007_ ),
    .B(\reg_module/_05011_ ),
    .Y(\reg_module/_05012_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12316_  (.A(\reg_module/_05001_ ),
    .X(\reg_module/_05013_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12317_  (.A(\reg_module/_05013_ ),
    .X(\reg_module/_05014_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12318_  (.A(\reg_module/_05014_ ),
    .B(\reg_module/gprf[32] ),
    .Y(\reg_module/_05015_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12319_  (.A(\reg_module/gprf[0] ),
    .B(net770),
    .Y(\reg_module/_05016_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12320_  (.A(\reg_module/_05015_ ),
    .B(net695),
    .C(\reg_module/_05016_ ),
    .Y(\reg_module/_05017_ ));
 sky130_fd_sc_hd__buf_1 \reg_module/_12321_  (.A(\reg_module/_05000_ ),
    .X(\reg_module/_05018_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12322_  (.A(\reg_module/_05018_ ),
    .X(\reg_module/_05019_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12323_  (.A(\reg_module/_05019_ ),
    .X(\reg_module/_05020_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12324_  (.A(\reg_module/_05020_ ),
    .B(\reg_module/gprf[96] ),
    .Y(\reg_module/_05021_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12325_  (.A(\reg_module/_04996_ ),
    .X(\reg_module/_05022_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12326_  (.A(\reg_module/_05022_ ),
    .X(\reg_module/_05023_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12327_  (.A(\reg_module/gprf[64] ),
    .B(net770),
    .Y(\reg_module/_05024_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12328_  (.A(\reg_module/_05021_ ),
    .B(\reg_module/_05023_ ),
    .C(\reg_module/_05024_ ),
    .Y(\reg_module/_05025_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12329_  (.A(\reg_module/_05017_ ),
    .B(\reg_module/_05025_ ),
    .Y(\reg_module/_05026_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12330_  (.A(\reg_module/_05026_ ),
    .B(net658),
    .Y(\reg_module/_05027_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12331_  (.A(\reg_module/_05012_ ),
    .B(\reg_module/_05027_ ),
    .C(net640),
    .Y(\reg_module/_05028_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12332_  (.A(\reg_module/_05001_ ),
    .X(\reg_module/_05029_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12333_  (.A(\reg_module/_05029_ ),
    .X(\reg_module/_05030_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12334_  (.A(\reg_module/_05030_ ),
    .B(\reg_module/gprf[288] ),
    .Y(\reg_module/_05031_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12335_  (.A(\reg_module/gprf[256] ),
    .B(net779),
    .Y(\reg_module/_05032_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12336_  (.A(\reg_module/_05031_ ),
    .B(net699),
    .C(\reg_module/_05032_ ),
    .Y(\reg_module/_05033_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_12337_  (.A(\reg_module/_05001_ ),
    .X(\reg_module/_05034_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12338_  (.A(\reg_module/_05034_ ),
    .X(\reg_module/_05035_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12339_  (.A(\reg_module/_05035_ ),
    .B(\reg_module/gprf[352] ),
    .Y(\reg_module/_05036_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12340_  (.A(\reg_module/_04996_ ),
    .X(\reg_module/_05037_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12341_  (.A(\reg_module/_05037_ ),
    .X(\reg_module/_05038_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12342_  (.A(\reg_module/gprf[320] ),
    .B(net779),
    .Y(\reg_module/_05039_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12343_  (.A(\reg_module/_05036_ ),
    .B(\reg_module/_05038_ ),
    .C(\reg_module/_05039_ ),
    .Y(\reg_module/_05040_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12344_  (.A(\reg_module/_05033_ ),
    .B(\reg_module/_05040_ ),
    .Y(\reg_module/_05041_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12345_  (.A(\reg_module/_05041_ ),
    .B(net661),
    .Y(\reg_module/_05042_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12346_  (.A(\reg_module/_05018_ ),
    .X(\reg_module/_05043_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12347_  (.A(\reg_module/_05043_ ),
    .X(\reg_module/_05044_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12348_  (.A(\reg_module/_05044_ ),
    .B(\reg_module/gprf[416] ),
    .Y(\reg_module/_05045_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12349_  (.A(\reg_module/gprf[384] ),
    .B(net771),
    .Y(\reg_module/_05046_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12350_  (.A(\reg_module/_05045_ ),
    .B(net696),
    .C(\reg_module/_05046_ ),
    .Y(\reg_module/_05047_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_12351_  (.A(\reg_module/_05000_ ),
    .X(\reg_module/_05048_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12352_  (.A(\reg_module/_05048_ ),
    .X(\reg_module/_05049_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12353_  (.A(\reg_module/_05049_ ),
    .B(\reg_module/gprf[480] ),
    .Y(\reg_module/_05050_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_12354_  (.A(\reg_module/_04996_ ),
    .X(\reg_module/_05051_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12355_  (.A(\reg_module/_05051_ ),
    .X(\reg_module/_05052_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12356_  (.A(\reg_module/gprf[448] ),
    .B(net771),
    .Y(\reg_module/_05053_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12357_  (.A(\reg_module/_05050_ ),
    .B(\reg_module/_05052_ ),
    .C(\reg_module/_05053_ ),
    .Y(\reg_module/_05054_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12358_  (.A(\reg_module/_05047_ ),
    .B(\reg_module/_05054_ ),
    .Y(\reg_module/_05055_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12359_  (.A(\reg_module/_05008_ ),
    .X(\reg_module/_05056_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12360_  (.A(\reg_module/_05056_ ),
    .X(\reg_module/_05057_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12361_  (.A(\reg_module/_05055_ ),
    .B(\reg_module/_05057_ ),
    .Y(\reg_module/_05058_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_12362_  (.A(net647),
    .Y(\reg_module/_05059_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12363_  (.A(\reg_module/_05059_ ),
    .X(\reg_module/_05060_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12364_  (.A(\reg_module/_05042_ ),
    .B(\reg_module/_05058_ ),
    .C(\reg_module/_05060_ ),
    .Y(\reg_module/_05061_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12365_  (.A(\reg_module/_05028_ ),
    .B(\reg_module/_05061_ ),
    .Y(\reg_module/_05062_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12366_  (.A(\reg_module/_05062_ ),
    .B(net632),
    .Y(\reg_module/_05063_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12367_  (.A(\reg_module/_05002_ ),
    .X(\reg_module/_05064_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12368_  (.A(\reg_module/_05064_ ),
    .B(\reg_module/gprf[800] ),
    .Y(\reg_module/_05065_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12369_  (.A(\reg_module/gprf[768] ),
    .B(net780),
    .Y(\reg_module/_05066_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12370_  (.A(\reg_module/_05065_ ),
    .B(net699),
    .C(\reg_module/_05066_ ),
    .Y(\reg_module/_05067_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12371_  (.A(\reg_module/_05001_ ),
    .X(\reg_module/_05068_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12372_  (.A(\reg_module/_05068_ ),
    .X(\reg_module/_05069_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12373_  (.A(\reg_module/_05069_ ),
    .B(\reg_module/gprf[864] ),
    .Y(\reg_module/_05070_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12374_  (.A(\reg_module/_04996_ ),
    .X(\reg_module/_05071_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12375_  (.A(\reg_module/_05071_ ),
    .X(\reg_module/_05072_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12376_  (.A(\reg_module/_05072_ ),
    .X(\reg_module/_05073_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12377_  (.A(\reg_module/gprf[832] ),
    .B(net780),
    .Y(\reg_module/_05074_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12378_  (.A(\reg_module/_05070_ ),
    .B(\reg_module/_05073_ ),
    .C(\reg_module/_05074_ ),
    .Y(\reg_module/_05075_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12379_  (.A(\reg_module/_05067_ ),
    .B(\reg_module/_05075_ ),
    .Y(\reg_module/_05076_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12380_  (.A(\reg_module/_05076_ ),
    .B(net658),
    .Y(\reg_module/_05077_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12381_  (.A(\reg_module/_05018_ ),
    .X(\reg_module/_05078_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12382_  (.A(\reg_module/_05078_ ),
    .X(\reg_module/_05079_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12383_  (.A(\reg_module/_05079_ ),
    .B(\reg_module/gprf[928] ),
    .Y(\reg_module/_05080_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12384_  (.A(\reg_module/gprf[896] ),
    .B(net772),
    .Y(\reg_module/_05081_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12385_  (.A(\reg_module/_05080_ ),
    .B(net696),
    .C(\reg_module/_05081_ ),
    .Y(\reg_module/_05082_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12386_  (.A(\reg_module/_05018_ ),
    .X(\reg_module/_05083_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_12387_  (.A(\reg_module/_05083_ ),
    .X(\reg_module/_05084_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12388_  (.A(\reg_module/_05084_ ),
    .B(\reg_module/gprf[992] ),
    .Y(\reg_module/_05085_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_12389_  (.A(\reg_module/_04996_ ),
    .X(\reg_module/_05086_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12390_  (.A(\reg_module/_05086_ ),
    .X(\reg_module/_05087_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12391_  (.A(\reg_module/gprf[960] ),
    .B(net772),
    .Y(\reg_module/_05088_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12392_  (.A(\reg_module/_05085_ ),
    .B(\reg_module/_05087_ ),
    .C(\reg_module/_05088_ ),
    .Y(\reg_module/_05089_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12393_  (.A(\reg_module/_05082_ ),
    .B(\reg_module/_05089_ ),
    .Y(\reg_module/_05090_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12394_  (.A(\reg_module/_05008_ ),
    .X(\reg_module/_05091_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12395_  (.A(\reg_module/_05091_ ),
    .X(\reg_module/_05092_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12396_  (.A(\reg_module/_05090_ ),
    .B(\reg_module/_05092_ ),
    .Y(\reg_module/_05093_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_12397_  (.A(\reg_module/_05059_ ),
    .X(\reg_module/_05094_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12398_  (.A(\reg_module/_05094_ ),
    .X(\reg_module/_05095_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12399_  (.A(\reg_module/_05077_ ),
    .B(\reg_module/_05093_ ),
    .C(\reg_module/_05095_ ),
    .Y(\reg_module/_05096_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12400_  (.A(\reg_module/_05069_ ),
    .B(\reg_module/gprf[672] ),
    .Y(\reg_module/_05097_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12401_  (.A(\reg_module/gprf[640] ),
    .B(net770),
    .Y(\reg_module/_05098_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12402_  (.A(\reg_module/_05097_ ),
    .B(net695),
    .C(\reg_module/_05098_ ),
    .Y(\reg_module/_05099_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_12403_  (.A(\reg_module/_05018_ ),
    .X(\reg_module/_05100_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12404_  (.A(\reg_module/_05100_ ),
    .X(\reg_module/_05101_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12405_  (.A(\reg_module/_05101_ ),
    .B(\reg_module/gprf[736] ),
    .Y(\reg_module/_05102_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12406_  (.A(\reg_module/_04997_ ),
    .X(\reg_module/_05103_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12407_  (.A(\reg_module/gprf[704] ),
    .B(net770),
    .Y(\reg_module/_05104_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12408_  (.A(\reg_module/_05102_ ),
    .B(\reg_module/_05103_ ),
    .C(\reg_module/_05104_ ),
    .Y(\reg_module/_05105_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12409_  (.A(\reg_module/_05099_ ),
    .B(\reg_module/_05105_ ),
    .Y(\reg_module/_05106_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12410_  (.A(\reg_module/_05106_ ),
    .B(\reg_module/_05092_ ),
    .Y(\reg_module/_05107_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12411_  (.A(\reg_module/_05018_ ),
    .X(\reg_module/_05108_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12412_  (.A(\reg_module/_05108_ ),
    .X(\reg_module/_05109_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12413_  (.A(\reg_module/_05109_ ),
    .B(\reg_module/gprf[544] ),
    .Y(\reg_module/_05110_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12414_  (.A(\reg_module/gprf[512] ),
    .B(net769),
    .Y(\reg_module/_05111_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12415_  (.A(\reg_module/_05110_ ),
    .B(net695),
    .C(\reg_module/_05111_ ),
    .Y(\reg_module/_05112_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12416_  (.A(\reg_module/_05000_ ),
    .X(\reg_module/_05113_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12417_  (.A(\reg_module/_05113_ ),
    .X(\reg_module/_05114_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12418_  (.A(\reg_module/_05114_ ),
    .B(\reg_module/gprf[608] ),
    .Y(\reg_module/_05115_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12419_  (.A(\reg_module/_05051_ ),
    .X(\reg_module/_05116_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12420_  (.A(\reg_module/gprf[576] ),
    .B(net769),
    .Y(\reg_module/_05117_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12421_  (.A(\reg_module/_05115_ ),
    .B(\reg_module/_05116_ ),
    .C(\reg_module/_05117_ ),
    .Y(\reg_module/_05118_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12422_  (.A(\reg_module/_05112_ ),
    .B(\reg_module/_05118_ ),
    .Y(\reg_module/_05119_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12423_  (.A(\reg_module/_05119_ ),
    .B(net658),
    .Y(\reg_module/_05120_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12424_  (.A(\reg_module/_05107_ ),
    .B(\reg_module/_05120_ ),
    .C(net640),
    .Y(\reg_module/_05121_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12425_  (.A(\reg_module/_05096_ ),
    .B(\reg_module/_05121_ ),
    .Y(\reg_module/_05122_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_12426_  (.A(net632),
    .Y(\reg_module/_05123_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12427_  (.A(\reg_module/_05123_ ),
    .X(\reg_module/_05124_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12428_  (.A(\reg_module/_05122_ ),
    .B(\reg_module/_05124_ ),
    .Y(\reg_module/_05125_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_12429_  (.A(\reg_module/_05063_ ),
    .B(\reg_module/_05125_ ),
    .Y(\wRs1Data[0] ));
 sky130_fd_sc_hd__inv_2 \reg_module/_12430_  (.A(net2170),
    .Y(\reg_module/_05126_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_12431_  (.A(net769),
    .B(\reg_module/_05126_ ),
    .Y(\reg_module/_05127_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12432_  (.A(\reg_module/gprf[193] ),
    .B(net768),
    .Y(\reg_module/_05128_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12433_  (.A(\reg_module/_05128_ ),
    .B(\reg_module/_05103_ ),
    .Y(\reg_module/_05129_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12434_  (.A(\reg_module/_05064_ ),
    .B(\reg_module/gprf[161] ),
    .Y(\reg_module/_05130_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12435_  (.A(\reg_module/gprf[129] ),
    .B(net768),
    .Y(\reg_module/_05131_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12436_  (.A(\reg_module/_05130_ ),
    .B(net695),
    .C(\reg_module/_05131_ ),
    .Y(\reg_module/_05132_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_12437_  (.A1(\reg_module/_05127_ ),
    .A2(\reg_module/_05129_ ),
    .B1(\reg_module/_05132_ ),
    .Y(\reg_module/_05133_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12438_  (.A(\reg_module/_05133_ ),
    .B(\reg_module/_05011_ ),
    .Y(\reg_module/_05134_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12439_  (.A(\reg_module/_05013_ ),
    .X(\reg_module/_05135_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12440_  (.A(\reg_module/_05135_ ),
    .B(\reg_module/gprf[33] ),
    .Y(\reg_module/_05136_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12441_  (.A(\reg_module/gprf[1] ),
    .B(net768),
    .Y(\reg_module/_05137_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12442_  (.A(\reg_module/_05136_ ),
    .B(net717),
    .C(\reg_module/_05137_ ),
    .Y(\reg_module/_05138_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12443_  (.A(\reg_module/_05019_ ),
    .X(\reg_module/_05139_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12444_  (.A(\reg_module/_05139_ ),
    .B(\reg_module/gprf[97] ),
    .Y(\reg_module/_05140_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12445_  (.A(\reg_module/gprf[65] ),
    .B(net768),
    .Y(\reg_module/_05141_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12446_  (.A(\reg_module/_05140_ ),
    .B(\reg_module/_05023_ ),
    .C(\reg_module/_05141_ ),
    .Y(\reg_module/_05142_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12447_  (.A(\reg_module/_05138_ ),
    .B(\reg_module/_05142_ ),
    .Y(\reg_module/_05143_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12448_  (.A(\reg_module/_05143_ ),
    .B(net658),
    .Y(\reg_module/_05144_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12449_  (.A(\reg_module/_05134_ ),
    .B(\reg_module/_05144_ ),
    .C(net640),
    .Y(\reg_module/_05145_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12450_  (.A(\reg_module/_05030_ ),
    .B(\reg_module/gprf[289] ),
    .Y(\reg_module/_05146_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12451_  (.A(\reg_module/gprf[257] ),
    .B(net779),
    .Y(\reg_module/_05147_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12452_  (.A(\reg_module/_05146_ ),
    .B(net699),
    .C(\reg_module/_05147_ ),
    .Y(\reg_module/_05148_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12453_  (.A(\reg_module/_05078_ ),
    .X(\reg_module/_05149_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12454_  (.A(\reg_module/_05149_ ),
    .B(\reg_module/gprf[353] ),
    .Y(\reg_module/_05150_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12455_  (.A(\reg_module/gprf[321] ),
    .B(net772),
    .Y(\reg_module/_05151_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12456_  (.A(\reg_module/_05150_ ),
    .B(\reg_module/_05038_ ),
    .C(\reg_module/_05151_ ),
    .Y(\reg_module/_05152_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12457_  (.A(\reg_module/_05148_ ),
    .B(\reg_module/_05152_ ),
    .Y(\reg_module/_05153_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12458_  (.A(\reg_module/_05153_ ),
    .B(net658),
    .Y(\reg_module/_05154_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12459_  (.A(\reg_module/_05044_ ),
    .B(\reg_module/gprf[417] ),
    .Y(\reg_module/_05155_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12460_  (.A(\reg_module/gprf[385] ),
    .B(net771),
    .Y(\reg_module/_05156_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12461_  (.A(\reg_module/_05155_ ),
    .B(net696),
    .C(\reg_module/_05156_ ),
    .Y(\reg_module/_05157_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12462_  (.A(\reg_module/_05049_ ),
    .B(\reg_module/gprf[481] ),
    .Y(\reg_module/_05158_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12463_  (.A(\reg_module/gprf[449] ),
    .B(net771),
    .Y(\reg_module/_05159_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12464_  (.A(\reg_module/_05158_ ),
    .B(\reg_module/_05052_ ),
    .C(\reg_module/_05159_ ),
    .Y(\reg_module/_05160_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12465_  (.A(\reg_module/_05157_ ),
    .B(\reg_module/_05160_ ),
    .Y(\reg_module/_05161_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12466_  (.A(\reg_module/_05161_ ),
    .B(\reg_module/_05057_ ),
    .Y(\reg_module/_05162_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12467_  (.A(\reg_module/_05154_ ),
    .B(\reg_module/_05162_ ),
    .C(\reg_module/_05060_ ),
    .Y(\reg_module/_05163_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12468_  (.A(\reg_module/_05145_ ),
    .B(\reg_module/_05163_ ),
    .Y(\reg_module/_05164_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12469_  (.A(\reg_module/_05164_ ),
    .B(net633),
    .Y(\reg_module/_05165_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12470_  (.A(\reg_module/_05064_ ),
    .B(\reg_module/gprf[801] ),
    .Y(\reg_module/_05166_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12471_  (.A(\reg_module/gprf[769] ),
    .B(net821),
    .Y(\reg_module/_05167_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12472_  (.A(\reg_module/_05166_ ),
    .B(net722),
    .C(\reg_module/_05167_ ),
    .Y(\reg_module/_05168_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12473_  (.A(\reg_module/_05069_ ),
    .B(\reg_module/gprf[865] ),
    .Y(\reg_module/_05169_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12474_  (.A(\reg_module/_05072_ ),
    .X(\reg_module/_05170_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12475_  (.A(\reg_module/gprf[833] ),
    .B(net821),
    .Y(\reg_module/_05171_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12476_  (.A(\reg_module/_05169_ ),
    .B(\reg_module/_05170_ ),
    .C(\reg_module/_05171_ ),
    .Y(\reg_module/_05172_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12477_  (.A(\reg_module/_05168_ ),
    .B(\reg_module/_05172_ ),
    .Y(\reg_module/_05173_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12478_  (.A(\reg_module/_05173_ ),
    .B(net661),
    .Y(\reg_module/_05174_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12479_  (.A(\reg_module/_05079_ ),
    .B(\reg_module/gprf[929] ),
    .Y(\reg_module/_05175_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12480_  (.A(\reg_module/gprf[897] ),
    .B(net772),
    .Y(\reg_module/_05176_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12481_  (.A(\reg_module/_05175_ ),
    .B(net696),
    .C(\reg_module/_05176_ ),
    .Y(\reg_module/_05177_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12482_  (.A(\reg_module/_05083_ ),
    .X(\reg_module/_05178_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12483_  (.A(\reg_module/_05178_ ),
    .B(\reg_module/gprf[993] ),
    .Y(\reg_module/_05179_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12484_  (.A(\reg_module/gprf[961] ),
    .B(net771),
    .Y(\reg_module/_05180_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12485_  (.A(\reg_module/_05179_ ),
    .B(\reg_module/_05087_ ),
    .C(\reg_module/_05180_ ),
    .Y(\reg_module/_05181_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12486_  (.A(\reg_module/_05177_ ),
    .B(\reg_module/_05181_ ),
    .Y(\reg_module/_05182_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12487_  (.A(\reg_module/_05091_ ),
    .X(\reg_module/_05183_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12488_  (.A(\reg_module/_05182_ ),
    .B(\reg_module/_05183_ ),
    .Y(\reg_module/_05184_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12489_  (.A(\reg_module/_05174_ ),
    .B(\reg_module/_05184_ ),
    .C(\reg_module/_05095_ ),
    .Y(\reg_module/_05185_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12490_  (.A(\reg_module/_05069_ ),
    .B(\reg_module/gprf[673] ),
    .Y(\reg_module/_05186_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12491_  (.A(\reg_module/gprf[641] ),
    .B(net769),
    .Y(\reg_module/_05187_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12492_  (.A(\reg_module/_05186_ ),
    .B(net695),
    .C(\reg_module/_05187_ ),
    .Y(\reg_module/_05188_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12493_  (.A(\reg_module/_05101_ ),
    .B(\reg_module/gprf[737] ),
    .Y(\reg_module/_05189_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12494_  (.A(\reg_module/gprf[705] ),
    .B(net768),
    .Y(\reg_module/_05190_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12495_  (.A(\reg_module/_05189_ ),
    .B(\reg_module/_05103_ ),
    .C(\reg_module/_05190_ ),
    .Y(\reg_module/_05191_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12496_  (.A(\reg_module/_05188_ ),
    .B(\reg_module/_05191_ ),
    .Y(\reg_module/_05192_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12497_  (.A(\reg_module/_05192_ ),
    .B(\reg_module/_05092_ ),
    .Y(\reg_module/_05193_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12498_  (.A(\reg_module/_05109_ ),
    .B(\reg_module/gprf[545] ),
    .Y(\reg_module/_05194_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12499_  (.A(\reg_module/gprf[513] ),
    .B(net811),
    .Y(\reg_module/_05195_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12500_  (.A(\reg_module/_05194_ ),
    .B(net717),
    .C(\reg_module/_05195_ ),
    .Y(\reg_module/_05196_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12501_  (.A(\reg_module/_05114_ ),
    .B(\reg_module/gprf[609] ),
    .Y(\reg_module/_05197_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12502_  (.A(\reg_module/gprf[577] ),
    .B(net769),
    .Y(\reg_module/_05198_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12503_  (.A(\reg_module/_05197_ ),
    .B(\reg_module/_05116_ ),
    .C(\reg_module/_05198_ ),
    .Y(\reg_module/_05199_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12504_  (.A(\reg_module/_05196_ ),
    .B(\reg_module/_05199_ ),
    .Y(\reg_module/_05200_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12505_  (.A(\reg_module/_05200_ ),
    .B(net658),
    .Y(\reg_module/_05201_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12506_  (.A(\reg_module/_05193_ ),
    .B(\reg_module/_05201_ ),
    .C(net641),
    .Y(\reg_module/_05202_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12507_  (.A(\reg_module/_05185_ ),
    .B(\reg_module/_05202_ ),
    .Y(\reg_module/_05203_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_12508_  (.A(\reg_module/_05123_ ),
    .X(\reg_module/_05204_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12509_  (.A(\reg_module/_05203_ ),
    .B(\reg_module/_05204_ ),
    .Y(\reg_module/_05205_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_12510_  (.A(\reg_module/_05165_ ),
    .B(\reg_module/_05205_ ),
    .Y(\wRs1Data[1] ));
 sky130_fd_sc_hd__inv_2 \reg_module/_12511_  (.A(net2218),
    .Y(\reg_module/_05206_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_12512_  (.A(net810),
    .B(\reg_module/_05206_ ),
    .Y(\reg_module/_05207_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12513_  (.A(\reg_module/gprf[194] ),
    .B(net810),
    .Y(\reg_module/_05208_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12514_  (.A(\reg_module/_05208_ ),
    .B(\reg_module/_05103_ ),
    .Y(\reg_module/_05209_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12515_  (.A(\reg_module/_05064_ ),
    .B(\reg_module/gprf[162] ),
    .Y(\reg_module/_05210_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12516_  (.A(\reg_module/gprf[130] ),
    .B(net810),
    .Y(\reg_module/_05211_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12517_  (.A(\reg_module/_05210_ ),
    .B(net717),
    .C(\reg_module/_05211_ ),
    .Y(\reg_module/_05212_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_12518_  (.A1(\reg_module/_05207_ ),
    .A2(\reg_module/_05209_ ),
    .B1(\reg_module/_05212_ ),
    .Y(\reg_module/_05213_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12519_  (.A(\reg_module/_05213_ ),
    .B(\reg_module/_05011_ ),
    .Y(\reg_module/_05214_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12520_  (.A(\reg_module/_05135_ ),
    .B(\reg_module/gprf[34] ),
    .Y(\reg_module/_05215_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12521_  (.A(\reg_module/gprf[2] ),
    .B(net810),
    .Y(\reg_module/_05216_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12522_  (.A(\reg_module/_05215_ ),
    .B(net717),
    .C(\reg_module/_05216_ ),
    .Y(\reg_module/_05217_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12523_  (.A(\reg_module/_05139_ ),
    .B(\reg_module/gprf[98] ),
    .Y(\reg_module/_05218_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12524_  (.A(\reg_module/gprf[66] ),
    .B(net811),
    .Y(\reg_module/_05219_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12525_  (.A(\reg_module/_05218_ ),
    .B(\reg_module/_05023_ ),
    .C(\reg_module/_05219_ ),
    .Y(\reg_module/_05220_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12526_  (.A(\reg_module/_05217_ ),
    .B(\reg_module/_05220_ ),
    .Y(\reg_module/_05221_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12527_  (.A(\reg_module/_05221_ ),
    .B(net672),
    .Y(\reg_module/_05222_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12528_  (.A(\reg_module/_05214_ ),
    .B(\reg_module/_05222_ ),
    .C(net647),
    .Y(\reg_module/_05223_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12529_  (.A(\reg_module/_05029_ ),
    .X(\reg_module/_05224_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12530_  (.A(\reg_module/_05224_ ),
    .B(\reg_module/gprf[290] ),
    .Y(\reg_module/_05225_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12531_  (.A(\reg_module/gprf[258] ),
    .B(net820),
    .Y(\reg_module/_05226_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12532_  (.A(\reg_module/_05225_ ),
    .B(net722),
    .C(\reg_module/_05226_ ),
    .Y(\reg_module/_05227_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12533_  (.A(\reg_module/_05149_ ),
    .B(\reg_module/gprf[354] ),
    .Y(\reg_module/_05228_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12534_  (.A(\reg_module/gprf[322] ),
    .B(net820),
    .Y(\reg_module/_05229_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12535_  (.A(\reg_module/_05228_ ),
    .B(\reg_module/_05038_ ),
    .C(\reg_module/_05229_ ),
    .Y(\reg_module/_05230_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12536_  (.A(\reg_module/_05227_ ),
    .B(\reg_module/_05230_ ),
    .Y(\reg_module/_05231_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12537_  (.A(\reg_module/_05231_ ),
    .B(net673),
    .Y(\reg_module/_05232_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12538_  (.A(\reg_module/_05044_ ),
    .B(\reg_module/gprf[418] ),
    .Y(\reg_module/_05233_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12539_  (.A(\reg_module/gprf[386] ),
    .B(net812),
    .Y(\reg_module/_05234_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12540_  (.A(\reg_module/_05233_ ),
    .B(net717),
    .C(\reg_module/_05234_ ),
    .Y(\reg_module/_05235_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12541_  (.A(\reg_module/_05049_ ),
    .B(\reg_module/gprf[482] ),
    .Y(\reg_module/_05236_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12542_  (.A(\reg_module/gprf[450] ),
    .B(net812),
    .Y(\reg_module/_05237_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12543_  (.A(\reg_module/_05236_ ),
    .B(\reg_module/_05052_ ),
    .C(\reg_module/_05237_ ),
    .Y(\reg_module/_05238_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12544_  (.A(\reg_module/_05235_ ),
    .B(\reg_module/_05238_ ),
    .Y(\reg_module/_05239_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12545_  (.A(\reg_module/_05239_ ),
    .B(\reg_module/_05057_ ),
    .Y(\reg_module/_05240_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12546_  (.A(\reg_module/_05232_ ),
    .B(\reg_module/_05240_ ),
    .C(\reg_module/_05060_ ),
    .Y(\reg_module/_05241_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12547_  (.A(\reg_module/_05223_ ),
    .B(\reg_module/_05241_ ),
    .Y(\reg_module/_05242_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12548_  (.A(\reg_module/_05242_ ),
    .B(net633),
    .Y(\reg_module/_05243_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12549_  (.A(\reg_module/_05064_ ),
    .B(\reg_module/gprf[802] ),
    .Y(\reg_module/_05244_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12550_  (.A(\reg_module/gprf[770] ),
    .B(net820),
    .Y(\reg_module/_05245_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12551_  (.A(\reg_module/_05244_ ),
    .B(net722),
    .C(\reg_module/_05245_ ),
    .Y(\reg_module/_05246_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12552_  (.A(\reg_module/_05069_ ),
    .B(\reg_module/gprf[866] ),
    .Y(\reg_module/_05247_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12553_  (.A(\reg_module/gprf[834] ),
    .B(net820),
    .Y(\reg_module/_05248_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12554_  (.A(\reg_module/_05247_ ),
    .B(\reg_module/_05170_ ),
    .C(\reg_module/_05248_ ),
    .Y(\reg_module/_05249_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12555_  (.A(\reg_module/_05246_ ),
    .B(\reg_module/_05249_ ),
    .Y(\reg_module/_05250_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12556_  (.A(\reg_module/_05250_ ),
    .B(net672),
    .Y(\reg_module/_05251_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12557_  (.A(\reg_module/_05079_ ),
    .B(\reg_module/gprf[930] ),
    .Y(\reg_module/_05252_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12558_  (.A(\reg_module/gprf[898] ),
    .B(net812),
    .Y(\reg_module/_05253_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12559_  (.A(\reg_module/_05252_ ),
    .B(net718),
    .C(\reg_module/_05253_ ),
    .Y(\reg_module/_05254_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12560_  (.A(\reg_module/_05178_ ),
    .B(\reg_module/gprf[994] ),
    .Y(\reg_module/_05255_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12561_  (.A(\reg_module/_05086_ ),
    .X(\reg_module/_05256_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12562_  (.A(\reg_module/gprf[962] ),
    .B(net813),
    .Y(\reg_module/_05257_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12563_  (.A(\reg_module/_05255_ ),
    .B(\reg_module/_05256_ ),
    .C(\reg_module/_05257_ ),
    .Y(\reg_module/_05258_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12564_  (.A(\reg_module/_05254_ ),
    .B(\reg_module/_05258_ ),
    .Y(\reg_module/_05259_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12565_  (.A(\reg_module/_05259_ ),
    .B(\reg_module/_05183_ ),
    .Y(\reg_module/_05260_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12566_  (.A(\reg_module/_05251_ ),
    .B(\reg_module/_05260_ ),
    .C(\reg_module/_05095_ ),
    .Y(\reg_module/_05261_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12567_  (.A(\reg_module/_05068_ ),
    .X(\reg_module/_05262_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12568_  (.A(\reg_module/_05262_ ),
    .B(\reg_module/gprf[674] ),
    .Y(\reg_module/_05263_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12569_  (.A(\reg_module/gprf[642] ),
    .B(net811),
    .Y(\reg_module/_05264_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12570_  (.A(\reg_module/_05263_ ),
    .B(net719),
    .C(\reg_module/_05264_ ),
    .Y(\reg_module/_05265_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12571_  (.A(\reg_module/_05101_ ),
    .B(\reg_module/gprf[738] ),
    .Y(\reg_module/_05266_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12572_  (.A(\reg_module/gprf[706] ),
    .B(net815),
    .Y(\reg_module/_05267_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12573_  (.A(\reg_module/_05266_ ),
    .B(\reg_module/_05103_ ),
    .C(\reg_module/_05267_ ),
    .Y(\reg_module/_05268_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12574_  (.A(\reg_module/_05265_ ),
    .B(\reg_module/_05268_ ),
    .Y(\reg_module/_05269_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12575_  (.A(\reg_module/_05269_ ),
    .B(\reg_module/_05092_ ),
    .Y(\reg_module/_05270_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12576_  (.A(\reg_module/_05109_ ),
    .B(\reg_module/gprf[546] ),
    .Y(\reg_module/_05271_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12577_  (.A(\reg_module/gprf[514] ),
    .B(net815),
    .Y(\reg_module/_05272_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12578_  (.A(\reg_module/_05271_ ),
    .B(net717),
    .C(\reg_module/_05272_ ),
    .Y(\reg_module/_05273_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12579_  (.A(\reg_module/_05114_ ),
    .B(\reg_module/gprf[610] ),
    .Y(\reg_module/_05274_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12580_  (.A(\reg_module/gprf[578] ),
    .B(net810),
    .Y(\reg_module/_05275_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12581_  (.A(\reg_module/_05274_ ),
    .B(\reg_module/_05116_ ),
    .C(\reg_module/_05275_ ),
    .Y(\reg_module/_05276_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12582_  (.A(\reg_module/_05273_ ),
    .B(\reg_module/_05276_ ),
    .Y(\reg_module/_05277_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12583_  (.A(\reg_module/_05277_ ),
    .B(net672),
    .Y(\reg_module/_05278_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12584_  (.A(\reg_module/_05270_ ),
    .B(\reg_module/_05278_ ),
    .C(net647),
    .Y(\reg_module/_05279_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12585_  (.A(\reg_module/_05261_ ),
    .B(\reg_module/_05279_ ),
    .Y(\reg_module/_05280_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12586_  (.A(\reg_module/_05280_ ),
    .B(\reg_module/_05204_ ),
    .Y(\reg_module/_05281_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_12587_  (.A(\reg_module/_05243_ ),
    .B(\reg_module/_05281_ ),
    .Y(\wRs1Data[2] ));
 sky130_fd_sc_hd__buf_4 \reg_module/_12588_  (.A(\reg_module/_05113_ ),
    .X(\reg_module/_05282_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12589_  (.A(\reg_module/_05282_ ),
    .X(\reg_module/_05283_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12590_  (.A(\reg_module/_05283_ ),
    .B(\reg_module/gprf[547] ),
    .Y(\reg_module/_05284_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12591_  (.A(\reg_module/gprf[515] ),
    .B(net830),
    .Y(\reg_module/_05285_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12592_  (.A(\reg_module/_05284_ ),
    .B(net727),
    .C(\reg_module/_05285_ ),
    .Y(\reg_module/_05286_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12593_  (.A(\reg_module/_05001_ ),
    .X(\reg_module/_05287_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12594_  (.A(\reg_module/_05287_ ),
    .X(\reg_module/_05288_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12595_  (.A(\reg_module/_05288_ ),
    .B(\reg_module/gprf[611] ),
    .Y(\reg_module/_05289_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_12596_  (.A(\reg_module/_05071_ ),
    .X(\reg_module/_05290_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12597_  (.A(\reg_module/_05290_ ),
    .X(\reg_module/_05291_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12598_  (.A(\reg_module/gprf[579] ),
    .B(net831),
    .Y(\reg_module/_05292_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12599_  (.A(\reg_module/_05289_ ),
    .B(\reg_module/_05291_ ),
    .C(\reg_module/_05292_ ),
    .Y(\reg_module/_05293_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12600_  (.A(\reg_module/_05286_ ),
    .B(\reg_module/_05293_ ),
    .Y(\reg_module/_05294_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12601_  (.A(\reg_module/_05294_ ),
    .B(net676),
    .Y(\reg_module/_05295_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12602_  (.A(\reg_module/_05135_ ),
    .B(\reg_module/gprf[675] ),
    .Y(\reg_module/_05296_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12603_  (.A(\reg_module/gprf[643] ),
    .B(net816),
    .Y(\reg_module/_05297_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12604_  (.A(\reg_module/_05296_ ),
    .B(net719),
    .C(\reg_module/_05297_ ),
    .Y(\reg_module/_05298_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12605_  (.A(\reg_module/_05139_ ),
    .B(\reg_module/gprf[739] ),
    .Y(\reg_module/_05299_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12606_  (.A(\reg_module/_05022_ ),
    .X(\reg_module/_05300_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12607_  (.A(\reg_module/gprf[707] ),
    .B(net816),
    .Y(\reg_module/_05301_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12608_  (.A(\reg_module/_05299_ ),
    .B(\reg_module/_05300_ ),
    .C(\reg_module/_05301_ ),
    .Y(\reg_module/_05302_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12609_  (.A(\reg_module/_05298_ ),
    .B(\reg_module/_05302_ ),
    .Y(\reg_module/_05303_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12610_  (.A(\reg_module/_05010_ ),
    .X(\reg_module/_05304_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12611_  (.A(\reg_module/_05303_ ),
    .B(\reg_module/_05304_ ),
    .Y(\reg_module/_05305_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12612_  (.A(\reg_module/_05295_ ),
    .B(\reg_module/_05305_ ),
    .C(net647),
    .Y(\reg_module/_05306_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12613_  (.A(\reg_module/_05224_ ),
    .B(\reg_module/gprf[803] ),
    .Y(\reg_module/_05307_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12614_  (.A(\reg_module/gprf[771] ),
    .B(net825),
    .Y(\reg_module/_05308_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12615_  (.A(\reg_module/_05307_ ),
    .B(net724),
    .C(\reg_module/_05308_ ),
    .Y(\reg_module/_05309_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12616_  (.A(\reg_module/_05149_ ),
    .B(\reg_module/gprf[867] ),
    .Y(\reg_module/_05310_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12617_  (.A(\reg_module/gprf[835] ),
    .B(net817),
    .Y(\reg_module/_05311_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12618_  (.A(\reg_module/_05310_ ),
    .B(\reg_module/_05038_ ),
    .C(\reg_module/_05311_ ),
    .Y(\reg_module/_05312_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12619_  (.A(\reg_module/_05309_ ),
    .B(\reg_module/_05312_ ),
    .Y(\reg_module/_05313_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12620_  (.A(\reg_module/_05313_ ),
    .B(net671),
    .Y(\reg_module/_05314_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12621_  (.A(\reg_module/_05043_ ),
    .X(\reg_module/_05315_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12622_  (.A(\reg_module/_05315_ ),
    .B(\reg_module/gprf[931] ),
    .Y(\reg_module/_05316_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12623_  (.A(\reg_module/gprf[899] ),
    .B(net817),
    .Y(\reg_module/_05317_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12624_  (.A(\reg_module/_05316_ ),
    .B(net720),
    .C(\reg_module/_05317_ ),
    .Y(\reg_module/_05318_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12625_  (.A(\reg_module/_05049_ ),
    .B(\reg_module/gprf[995] ),
    .Y(\reg_module/_05319_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12626_  (.A(\reg_module/gprf[963] ),
    .B(net817),
    .Y(\reg_module/_05320_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12627_  (.A(\reg_module/_05319_ ),
    .B(\reg_module/_05052_ ),
    .C(\reg_module/_05320_ ),
    .Y(\reg_module/_05321_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12628_  (.A(\reg_module/_05318_ ),
    .B(\reg_module/_05321_ ),
    .Y(\reg_module/_05322_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12629_  (.A(\reg_module/_05322_ ),
    .B(\reg_module/_05057_ ),
    .Y(\reg_module/_05323_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12630_  (.A(\reg_module/_05314_ ),
    .B(\reg_module/_05323_ ),
    .C(\reg_module/_05060_ ),
    .Y(\reg_module/_05324_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12631_  (.A(\reg_module/_05306_ ),
    .B(\reg_module/_05324_ ),
    .Y(\reg_module/_05325_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12632_  (.A(\reg_module/_05204_ ),
    .X(\reg_module/_05326_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12633_  (.A(\reg_module/_05325_ ),
    .B(\reg_module/_05326_ ),
    .Y(\reg_module/_05327_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12634_  (.A(\reg_module/_05064_ ),
    .B(\reg_module/gprf[291] ),
    .Y(\reg_module/_05328_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12635_  (.A(\reg_module/gprf[259] ),
    .B(net825),
    .Y(\reg_module/_05329_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12636_  (.A(\reg_module/_05328_ ),
    .B(net724),
    .C(\reg_module/_05329_ ),
    .Y(\reg_module/_05330_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12637_  (.A(\reg_module/_05262_ ),
    .B(\reg_module/gprf[355] ),
    .Y(\reg_module/_05331_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12638_  (.A(\reg_module/gprf[323] ),
    .B(net817),
    .Y(\reg_module/_05332_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12639_  (.A(\reg_module/_05331_ ),
    .B(\reg_module/_05170_ ),
    .C(\reg_module/_05332_ ),
    .Y(\reg_module/_05333_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12640_  (.A(\reg_module/_05330_ ),
    .B(\reg_module/_05333_ ),
    .Y(\reg_module/_05334_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12641_  (.A(\reg_module/_05334_ ),
    .B(net672),
    .Y(\reg_module/_05335_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12642_  (.A(\reg_module/_05079_ ),
    .B(\reg_module/gprf[419] ),
    .Y(\reg_module/_05336_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12643_  (.A(\reg_module/gprf[387] ),
    .B(net813),
    .Y(\reg_module/_05337_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12644_  (.A(\reg_module/_05336_ ),
    .B(net718),
    .C(\reg_module/_05337_ ),
    .Y(\reg_module/_05338_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12645_  (.A(\reg_module/_05178_ ),
    .B(\reg_module/gprf[483] ),
    .Y(\reg_module/_05339_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12646_  (.A(\reg_module/gprf[451] ),
    .B(net812),
    .Y(\reg_module/_05340_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12647_  (.A(\reg_module/_05339_ ),
    .B(\reg_module/_05256_ ),
    .C(\reg_module/_05340_ ),
    .Y(\reg_module/_05341_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12648_  (.A(\reg_module/_05338_ ),
    .B(\reg_module/_05341_ ),
    .Y(\reg_module/_05342_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12649_  (.A(\reg_module/_05342_ ),
    .B(\reg_module/_05183_ ),
    .Y(\reg_module/_05343_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12650_  (.A(\reg_module/_05335_ ),
    .B(\reg_module/_05343_ ),
    .C(\reg_module/_05095_ ),
    .Y(\reg_module/_05344_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12651_  (.A(\reg_module/_05262_ ),
    .B(\reg_module/gprf[35] ),
    .Y(\reg_module/_05345_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12652_  (.A(\reg_module/gprf[3] ),
    .B(net815),
    .Y(\reg_module/_05346_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12653_  (.A(\reg_module/_05345_ ),
    .B(net719),
    .C(\reg_module/_05346_ ),
    .Y(\reg_module/_05347_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12654_  (.A(\reg_module/_05101_ ),
    .B(\reg_module/gprf[99] ),
    .Y(\reg_module/_05348_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12655_  (.A(\reg_module/gprf[67] ),
    .B(net810),
    .Y(\reg_module/_05349_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12656_  (.A(\reg_module/_05348_ ),
    .B(\reg_module/_05103_ ),
    .C(\reg_module/_05349_ ),
    .Y(\reg_module/_05350_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12657_  (.A(\reg_module/_05347_ ),
    .B(\reg_module/_05350_ ),
    .Y(\reg_module/_05351_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12658_  (.A(\reg_module/_05351_ ),
    .B(net671),
    .Y(\reg_module/_05352_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12659_  (.A(\reg_module/_05108_ ),
    .X(\reg_module/_05353_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12660_  (.A(\reg_module/_05353_ ),
    .B(\reg_module/gprf[163] ),
    .Y(\reg_module/_05354_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12661_  (.A(\reg_module/gprf[131] ),
    .B(net815),
    .Y(\reg_module/_05355_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12662_  (.A(\reg_module/_05354_ ),
    .B(net719),
    .C(\reg_module/_05355_ ),
    .Y(\reg_module/_05356_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12663_  (.A(\reg_module/_05113_ ),
    .X(\reg_module/_05357_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12664_  (.A(\reg_module/_05357_ ),
    .B(\reg_module/gprf[227] ),
    .Y(\reg_module/_05358_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12665_  (.A(\reg_module/gprf[195] ),
    .B(net815),
    .Y(\reg_module/_05359_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12666_  (.A(\reg_module/_05358_ ),
    .B(\reg_module/_05116_ ),
    .C(\reg_module/_05359_ ),
    .Y(\reg_module/_05360_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12667_  (.A(\reg_module/_05356_ ),
    .B(\reg_module/_05360_ ),
    .Y(\reg_module/_05361_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_12668_  (.A(\reg_module/_05009_ ),
    .X(\reg_module/_05362_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12669_  (.A(\reg_module/_05361_ ),
    .B(\reg_module/_05362_ ),
    .Y(\reg_module/_05363_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12670_  (.A(\reg_module/_05352_ ),
    .B(\reg_module/_05363_ ),
    .C(net647),
    .Y(\reg_module/_05364_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12671_  (.A(\reg_module/_05344_ ),
    .B(\reg_module/_05364_ ),
    .Y(\reg_module/_05365_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12672_  (.A(\reg_module/_05365_ ),
    .B(net633),
    .Y(\reg_module/_05366_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_12673_  (.A(\reg_module/_05327_ ),
    .B(\reg_module/_05366_ ),
    .Y(\wRs1Data[3] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12674_  (.A(\reg_module/_05283_ ),
    .B(\reg_module/gprf[548] ),
    .Y(\reg_module/_05367_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12675_  (.A(\reg_module/gprf[516] ),
    .B(net830),
    .Y(\reg_module/_05368_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12676_  (.A(\reg_module/_05367_ ),
    .B(net727),
    .C(\reg_module/_05368_ ),
    .Y(\reg_module/_05369_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12677_  (.A(\reg_module/_05288_ ),
    .B(\reg_module/gprf[612] ),
    .Y(\reg_module/_05370_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12678_  (.A(\reg_module/gprf[580] ),
    .B(net830),
    .Y(\reg_module/_05371_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12679_  (.A(\reg_module/_05370_ ),
    .B(\reg_module/_05291_ ),
    .C(\reg_module/_05371_ ),
    .Y(\reg_module/_05372_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12680_  (.A(\reg_module/_05369_ ),
    .B(\reg_module/_05372_ ),
    .Y(\reg_module/_05373_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12681_  (.A(\reg_module/_05373_ ),
    .B(net671),
    .Y(\reg_module/_05374_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12682_  (.A(\reg_module/_05135_ ),
    .B(\reg_module/gprf[676] ),
    .Y(\reg_module/_05375_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12683_  (.A(\reg_module/gprf[644] ),
    .B(net815),
    .Y(\reg_module/_05376_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12684_  (.A(\reg_module/_05375_ ),
    .B(net719),
    .C(\reg_module/_05376_ ),
    .Y(\reg_module/_05377_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12685_  (.A(\reg_module/_05139_ ),
    .B(\reg_module/gprf[740] ),
    .Y(\reg_module/_05378_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12686_  (.A(\reg_module/gprf[708] ),
    .B(net816),
    .Y(\reg_module/_05379_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12687_  (.A(\reg_module/_05378_ ),
    .B(\reg_module/_05300_ ),
    .C(\reg_module/_05379_ ),
    .Y(\reg_module/_05380_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12688_  (.A(\reg_module/_05377_ ),
    .B(\reg_module/_05380_ ),
    .Y(\reg_module/_05381_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12689_  (.A(\reg_module/_05381_ ),
    .B(\reg_module/_05304_ ),
    .Y(\reg_module/_05382_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12690_  (.A(\reg_module/_05374_ ),
    .B(\reg_module/_05382_ ),
    .C(net647),
    .Y(\reg_module/_05383_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12691_  (.A(\reg_module/_05224_ ),
    .B(\reg_module/gprf[804] ),
    .Y(\reg_module/_05384_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12692_  (.A(\reg_module/gprf[772] ),
    .B(net824),
    .Y(\reg_module/_05385_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12693_  (.A(\reg_module/_05384_ ),
    .B(net724),
    .C(\reg_module/_05385_ ),
    .Y(\reg_module/_05386_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12694_  (.A(\reg_module/_05149_ ),
    .B(\reg_module/gprf[868] ),
    .Y(\reg_module/_05387_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12695_  (.A(\reg_module/gprf[836] ),
    .B(net818),
    .Y(\reg_module/_05388_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12696_  (.A(\reg_module/_05387_ ),
    .B(\reg_module/_05038_ ),
    .C(\reg_module/_05388_ ),
    .Y(\reg_module/_05389_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12697_  (.A(\reg_module/_05386_ ),
    .B(\reg_module/_05389_ ),
    .Y(\reg_module/_05390_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12698_  (.A(\reg_module/_05390_ ),
    .B(net671),
    .Y(\reg_module/_05391_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12699_  (.A(\reg_module/_05315_ ),
    .B(\reg_module/gprf[932] ),
    .Y(\reg_module/_05392_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12700_  (.A(\reg_module/gprf[900] ),
    .B(net818),
    .Y(\reg_module/_05393_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12701_  (.A(\reg_module/_05392_ ),
    .B(net720),
    .C(\reg_module/_05393_ ),
    .Y(\reg_module/_05394_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12702_  (.A(\reg_module/_05049_ ),
    .B(\reg_module/gprf[996] ),
    .Y(\reg_module/_05395_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12703_  (.A(\reg_module/gprf[964] ),
    .B(net818),
    .Y(\reg_module/_05396_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12704_  (.A(\reg_module/_05395_ ),
    .B(\reg_module/_05052_ ),
    .C(\reg_module/_05396_ ),
    .Y(\reg_module/_05397_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12705_  (.A(\reg_module/_05394_ ),
    .B(\reg_module/_05397_ ),
    .Y(\reg_module/_05398_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12706_  (.A(\reg_module/_05398_ ),
    .B(\reg_module/_05057_ ),
    .Y(\reg_module/_05399_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_12707_  (.A(\reg_module/_05059_ ),
    .X(\reg_module/_05400_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12708_  (.A(\reg_module/_05391_ ),
    .B(\reg_module/_05399_ ),
    .C(\reg_module/_05400_ ),
    .Y(\reg_module/_05401_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12709_  (.A(\reg_module/_05383_ ),
    .B(\reg_module/_05401_ ),
    .Y(\reg_module/_05402_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12710_  (.A(\reg_module/_05402_ ),
    .B(\reg_module/_05326_ ),
    .Y(\reg_module/_05403_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12711_  (.A(\reg_module/_05002_ ),
    .X(\reg_module/_05404_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12712_  (.A(\reg_module/_05404_ ),
    .B(\reg_module/gprf[292] ),
    .Y(\reg_module/_05405_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12713_  (.A(\reg_module/gprf[260] ),
    .B(net836),
    .Y(\reg_module/_05406_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12714_  (.A(\reg_module/_05405_ ),
    .B(net729),
    .C(\reg_module/_05406_ ),
    .Y(\reg_module/_05407_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12715_  (.A(\reg_module/_05262_ ),
    .B(\reg_module/gprf[356] ),
    .Y(\reg_module/_05408_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12716_  (.A(\reg_module/gprf[324] ),
    .B(net832),
    .Y(\reg_module/_05409_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12717_  (.A(\reg_module/_05408_ ),
    .B(\reg_module/_05170_ ),
    .C(\reg_module/_05409_ ),
    .Y(\reg_module/_05410_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12718_  (.A(\reg_module/_05407_ ),
    .B(\reg_module/_05410_ ),
    .Y(\reg_module/_05411_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12719_  (.A(\reg_module/_05411_ ),
    .B(net676),
    .Y(\reg_module/_05412_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12720_  (.A(\reg_module/_05079_ ),
    .B(\reg_module/gprf[420] ),
    .Y(\reg_module/_05413_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12721_  (.A(\reg_module/gprf[388] ),
    .B(net813),
    .Y(\reg_module/_05414_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12722_  (.A(\reg_module/_05413_ ),
    .B(net718),
    .C(\reg_module/_05414_ ),
    .Y(\reg_module/_05415_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12723_  (.A(\reg_module/_05178_ ),
    .B(\reg_module/gprf[484] ),
    .Y(\reg_module/_05416_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12724_  (.A(\reg_module/gprf[452] ),
    .B(net812),
    .Y(\reg_module/_05417_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12725_  (.A(\reg_module/_05416_ ),
    .B(\reg_module/_05256_ ),
    .C(\reg_module/_05417_ ),
    .Y(\reg_module/_05418_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12726_  (.A(\reg_module/_05415_ ),
    .B(\reg_module/_05418_ ),
    .Y(\reg_module/_05419_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12727_  (.A(\reg_module/_05419_ ),
    .B(\reg_module/_05183_ ),
    .Y(\reg_module/_05420_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12728_  (.A(\reg_module/_05412_ ),
    .B(\reg_module/_05420_ ),
    .C(\reg_module/_05095_ ),
    .Y(\reg_module/_05421_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12729_  (.A(\reg_module/_05262_ ),
    .B(\reg_module/gprf[36] ),
    .Y(\reg_module/_05422_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12730_  (.A(\reg_module/gprf[4] ),
    .B(net831),
    .Y(\reg_module/_05423_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12731_  (.A(\reg_module/_05422_ ),
    .B(net727),
    .C(\reg_module/_05423_ ),
    .Y(\reg_module/_05424_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12732_  (.A(\reg_module/_05101_ ),
    .B(\reg_module/gprf[100] ),
    .Y(\reg_module/_05425_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12733_  (.A(\reg_module/_04997_ ),
    .X(\reg_module/_05426_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12734_  (.A(\reg_module/gprf[68] ),
    .B(net832),
    .Y(\reg_module/_05427_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12735_  (.A(\reg_module/_05425_ ),
    .B(\reg_module/_05426_ ),
    .C(\reg_module/_05427_ ),
    .Y(\reg_module/_05428_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12736_  (.A(\reg_module/_05424_ ),
    .B(\reg_module/_05428_ ),
    .Y(\reg_module/_05429_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12737_  (.A(\reg_module/_05429_ ),
    .B(net676),
    .Y(\reg_module/_05430_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12738_  (.A(\reg_module/_05353_ ),
    .B(\reg_module/gprf[164] ),
    .Y(\reg_module/_05431_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12739_  (.A(\reg_module/gprf[132] ),
    .B(net830),
    .Y(\reg_module/_05432_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12740_  (.A(\reg_module/_05431_ ),
    .B(net727),
    .C(\reg_module/_05432_ ),
    .Y(\reg_module/_05433_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12741_  (.A(\reg_module/_05357_ ),
    .B(\reg_module/gprf[228] ),
    .Y(\reg_module/_05434_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12742_  (.A(\reg_module/_05071_ ),
    .X(\reg_module/_05435_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12743_  (.A(\reg_module/gprf[196] ),
    .B(net830),
    .Y(\reg_module/_05436_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12744_  (.A(\reg_module/_05434_ ),
    .B(\reg_module/_05435_ ),
    .C(\reg_module/_05436_ ),
    .Y(\reg_module/_05437_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12745_  (.A(\reg_module/_05433_ ),
    .B(\reg_module/_05437_ ),
    .Y(\reg_module/_05438_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12746_  (.A(\reg_module/_05438_ ),
    .B(\reg_module/_05362_ ),
    .Y(\reg_module/_05439_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12747_  (.A(\reg_module/_05430_ ),
    .B(\reg_module/_05439_ ),
    .C(net649),
    .Y(\reg_module/_05440_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12748_  (.A(\reg_module/_05421_ ),
    .B(\reg_module/_05440_ ),
    .Y(\reg_module/_05441_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12749_  (.A(\reg_module/_05441_ ),
    .B(net633),
    .Y(\reg_module/_05442_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_12750_  (.A(\reg_module/_05403_ ),
    .B(\reg_module/_05442_ ),
    .Y(\wRs1Data[4] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12751_  (.A(\reg_module/_05283_ ),
    .B(\reg_module/gprf[549] ),
    .Y(\reg_module/_05443_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12752_  (.A(\reg_module/gprf[517] ),
    .B(net830),
    .Y(\reg_module/_05444_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12753_  (.A(\reg_module/_05443_ ),
    .B(net727),
    .C(\reg_module/_05444_ ),
    .Y(\reg_module/_05445_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12754_  (.A(\reg_module/_05288_ ),
    .B(\reg_module/gprf[613] ),
    .Y(\reg_module/_05446_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12755_  (.A(\reg_module/gprf[581] ),
    .B(net832),
    .Y(\reg_module/_05447_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12756_  (.A(\reg_module/_05446_ ),
    .B(\reg_module/_05291_ ),
    .C(\reg_module/_05447_ ),
    .Y(\reg_module/_05448_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12757_  (.A(\reg_module/_05445_ ),
    .B(\reg_module/_05448_ ),
    .Y(\reg_module/_05449_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12758_  (.A(\reg_module/_05449_ ),
    .B(net671),
    .Y(\reg_module/_05450_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12759_  (.A(\reg_module/_05135_ ),
    .B(\reg_module/gprf[677] ),
    .Y(\reg_module/_05451_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12760_  (.A(\reg_module/gprf[645] ),
    .B(net816),
    .Y(\reg_module/_05452_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12761_  (.A(\reg_module/_05451_ ),
    .B(net719),
    .C(\reg_module/_05452_ ),
    .Y(\reg_module/_05453_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12762_  (.A(\reg_module/_05139_ ),
    .B(\reg_module/gprf[741] ),
    .Y(\reg_module/_05454_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12763_  (.A(\reg_module/gprf[709] ),
    .B(net816),
    .Y(\reg_module/_05455_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12764_  (.A(\reg_module/_05454_ ),
    .B(\reg_module/_05300_ ),
    .C(\reg_module/_05455_ ),
    .Y(\reg_module/_05456_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12765_  (.A(\reg_module/_05453_ ),
    .B(\reg_module/_05456_ ),
    .Y(\reg_module/_05457_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12766_  (.A(\reg_module/_05457_ ),
    .B(\reg_module/_05304_ ),
    .Y(\reg_module/_05458_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12767_  (.A(\reg_module/_05450_ ),
    .B(\reg_module/_05458_ ),
    .C(net648),
    .Y(\reg_module/_05459_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12768_  (.A(\reg_module/_05224_ ),
    .B(\reg_module/gprf[805] ),
    .Y(\reg_module/_05460_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12769_  (.A(\reg_module/gprf[773] ),
    .B(net824),
    .Y(\reg_module/_05461_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12770_  (.A(\reg_module/_05460_ ),
    .B(net725),
    .C(\reg_module/_05461_ ),
    .Y(\reg_module/_05462_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12771_  (.A(\reg_module/_05149_ ),
    .B(\reg_module/gprf[869] ),
    .Y(\reg_module/_05463_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12772_  (.A(\reg_module/_05037_ ),
    .X(\reg_module/_05464_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12773_  (.A(\reg_module/gprf[837] ),
    .B(net817),
    .Y(\reg_module/_05465_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12774_  (.A(\reg_module/_05463_ ),
    .B(\reg_module/_05464_ ),
    .C(\reg_module/_05465_ ),
    .Y(\reg_module/_05466_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12775_  (.A(\reg_module/_05462_ ),
    .B(\reg_module/_05466_ ),
    .Y(\reg_module/_05467_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12776_  (.A(\reg_module/_05467_ ),
    .B(net671),
    .Y(\reg_module/_05468_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12777_  (.A(\reg_module/_05315_ ),
    .B(\reg_module/gprf[933] ),
    .Y(\reg_module/_05469_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12778_  (.A(\reg_module/gprf[901] ),
    .B(net817),
    .Y(\reg_module/_05470_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12779_  (.A(\reg_module/_05469_ ),
    .B(net720),
    .C(\reg_module/_05470_ ),
    .Y(\reg_module/_05471_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12780_  (.A(\reg_module/_05048_ ),
    .X(\reg_module/_05472_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12781_  (.A(\reg_module/_05472_ ),
    .B(\reg_module/gprf[997] ),
    .Y(\reg_module/_05473_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12782_  (.A(\reg_module/gprf[965] ),
    .B(net818),
    .Y(\reg_module/_05474_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12783_  (.A(\reg_module/_05473_ ),
    .B(\reg_module/_05052_ ),
    .C(\reg_module/_05474_ ),
    .Y(\reg_module/_05475_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12784_  (.A(\reg_module/_05471_ ),
    .B(\reg_module/_05475_ ),
    .Y(\reg_module/_05476_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_12785_  (.A(\reg_module/_05056_ ),
    .X(\reg_module/_05477_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12786_  (.A(\reg_module/_05476_ ),
    .B(\reg_module/_05477_ ),
    .Y(\reg_module/_05478_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12787_  (.A(\reg_module/_05468_ ),
    .B(\reg_module/_05478_ ),
    .C(\reg_module/_05400_ ),
    .Y(\reg_module/_05479_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12788_  (.A(\reg_module/_05459_ ),
    .B(\reg_module/_05479_ ),
    .Y(\reg_module/_05480_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12789_  (.A(\reg_module/_05480_ ),
    .B(\reg_module/_05326_ ),
    .Y(\reg_module/_05481_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12790_  (.A(\reg_module/_05404_ ),
    .B(\reg_module/gprf[293] ),
    .Y(\reg_module/_05482_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12791_  (.A(\reg_module/gprf[261] ),
    .B(net832),
    .Y(\reg_module/_05483_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12792_  (.A(\reg_module/_05482_ ),
    .B(net728),
    .C(\reg_module/_05483_ ),
    .Y(\reg_module/_05484_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12793_  (.A(\reg_module/_05262_ ),
    .B(\reg_module/gprf[357] ),
    .Y(\reg_module/_05485_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12794_  (.A(\reg_module/gprf[325] ),
    .B(net832),
    .Y(\reg_module/_05486_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12795_  (.A(\reg_module/_05485_ ),
    .B(\reg_module/_05170_ ),
    .C(\reg_module/_05486_ ),
    .Y(\reg_module/_05487_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12796_  (.A(\reg_module/_05484_ ),
    .B(\reg_module/_05487_ ),
    .Y(\reg_module/_05488_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12797_  (.A(\reg_module/_05488_ ),
    .B(net676),
    .Y(\reg_module/_05489_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12798_  (.A(\reg_module/_05043_ ),
    .X(\reg_module/_05490_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12799_  (.A(\reg_module/_05490_ ),
    .B(\reg_module/gprf[421] ),
    .Y(\reg_module/_05491_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12800_  (.A(\reg_module/gprf[389] ),
    .B(net820),
    .Y(\reg_module/_05492_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12801_  (.A(\reg_module/_05491_ ),
    .B(net722),
    .C(\reg_module/_05492_ ),
    .Y(\reg_module/_05493_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12802_  (.A(\reg_module/_05178_ ),
    .B(\reg_module/gprf[485] ),
    .Y(\reg_module/_05494_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12803_  (.A(\reg_module/gprf[453] ),
    .B(net812),
    .Y(\reg_module/_05495_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12804_  (.A(\reg_module/_05494_ ),
    .B(\reg_module/_05256_ ),
    .C(\reg_module/_05495_ ),
    .Y(\reg_module/_05496_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12805_  (.A(\reg_module/_05493_ ),
    .B(\reg_module/_05496_ ),
    .Y(\reg_module/_05497_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12806_  (.A(\reg_module/_05497_ ),
    .B(\reg_module/_05183_ ),
    .Y(\reg_module/_05498_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12807_  (.A(\reg_module/_05489_ ),
    .B(\reg_module/_05498_ ),
    .C(\reg_module/_05095_ ),
    .Y(\reg_module/_05499_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12808_  (.A(\reg_module/_05068_ ),
    .X(\reg_module/_05500_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12809_  (.A(\reg_module/_05500_ ),
    .B(\reg_module/gprf[37] ),
    .Y(\reg_module/_05501_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12810_  (.A(\reg_module/gprf[5] ),
    .B(net834),
    .Y(\reg_module/_05502_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12811_  (.A(\reg_module/_05501_ ),
    .B(net728),
    .C(\reg_module/_05502_ ),
    .Y(\reg_module/_05503_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12812_  (.A(\reg_module/_05100_ ),
    .X(\reg_module/_05504_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12813_  (.A(\reg_module/_05504_ ),
    .B(\reg_module/gprf[101] ),
    .Y(\reg_module/_05505_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12814_  (.A(\reg_module/gprf[69] ),
    .B(net833),
    .Y(\reg_module/_05506_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12815_  (.A(\reg_module/_05505_ ),
    .B(\reg_module/_05426_ ),
    .C(\reg_module/_05506_ ),
    .Y(\reg_module/_05507_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12816_  (.A(\reg_module/_05503_ ),
    .B(\reg_module/_05507_ ),
    .Y(\reg_module/_05508_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12817_  (.A(\reg_module/_05508_ ),
    .B(net676),
    .Y(\reg_module/_05509_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12818_  (.A(\reg_module/_05353_ ),
    .B(\reg_module/gprf[165] ),
    .Y(\reg_module/_05510_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12819_  (.A(\reg_module/gprf[133] ),
    .B(net831),
    .Y(\reg_module/_05511_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12820_  (.A(\reg_module/_05510_ ),
    .B(net727),
    .C(\reg_module/_05511_ ),
    .Y(\reg_module/_05512_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12821_  (.A(\reg_module/_05357_ ),
    .B(\reg_module/gprf[229] ),
    .Y(\reg_module/_05513_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12822_  (.A(\reg_module/gprf[197] ),
    .B(net831),
    .Y(\reg_module/_05514_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12823_  (.A(\reg_module/_05513_ ),
    .B(\reg_module/_05435_ ),
    .C(\reg_module/_05514_ ),
    .Y(\reg_module/_05515_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12824_  (.A(\reg_module/_05512_ ),
    .B(\reg_module/_05515_ ),
    .Y(\reg_module/_05516_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12825_  (.A(\reg_module/_05516_ ),
    .B(\reg_module/_05362_ ),
    .Y(\reg_module/_05517_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12826_  (.A(\reg_module/_05509_ ),
    .B(\reg_module/_05517_ ),
    .C(net649),
    .Y(\reg_module/_05518_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12827_  (.A(\reg_module/_05499_ ),
    .B(\reg_module/_05518_ ),
    .Y(\reg_module/_05519_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12828_  (.A(\reg_module/_05519_ ),
    .B(net633),
    .Y(\reg_module/_05520_ ));
 sky130_fd_sc_hd__nand2_4 \reg_module/_12829_  (.A(\reg_module/_05481_ ),
    .B(\reg_module/_05520_ ),
    .Y(\wRs1Data[5] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12830_  (.A(\reg_module/_05283_ ),
    .B(\reg_module/gprf[806] ),
    .Y(\reg_module/_05521_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12831_  (.A(\reg_module/gprf[774] ),
    .B(net835),
    .Y(\reg_module/_05522_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12832_  (.A(\reg_module/_05521_ ),
    .B(net729),
    .C(\reg_module/_05522_ ),
    .Y(\reg_module/_05523_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12833_  (.A(\reg_module/_05288_ ),
    .B(\reg_module/gprf[870] ),
    .Y(\reg_module/_05524_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12834_  (.A(\reg_module/gprf[838] ),
    .B(net835),
    .Y(\reg_module/_05525_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12835_  (.A(\reg_module/_05524_ ),
    .B(\reg_module/_05291_ ),
    .C(\reg_module/_05525_ ),
    .Y(\reg_module/_05526_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12836_  (.A(\reg_module/_05523_ ),
    .B(\reg_module/_05526_ ),
    .Y(\reg_module/_05527_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12837_  (.A(\reg_module/_05527_ ),
    .B(net674),
    .Y(\reg_module/_05528_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12838_  (.A(\reg_module/_05135_ ),
    .B(\reg_module/gprf[934] ),
    .Y(\reg_module/_05529_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12839_  (.A(\reg_module/gprf[902] ),
    .B(net824),
    .Y(\reg_module/_05530_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12840_  (.A(\reg_module/_05529_ ),
    .B(net724),
    .C(\reg_module/_05530_ ),
    .Y(\reg_module/_05531_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12841_  (.A(\reg_module/_05139_ ),
    .B(\reg_module/gprf[998] ),
    .Y(\reg_module/_05532_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12842_  (.A(\reg_module/gprf[966] ),
    .B(net825),
    .Y(\reg_module/_05533_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12843_  (.A(\reg_module/_05532_ ),
    .B(\reg_module/_05300_ ),
    .C(\reg_module/_05533_ ),
    .Y(\reg_module/_05534_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12844_  (.A(\reg_module/_05531_ ),
    .B(\reg_module/_05534_ ),
    .Y(\reg_module/_05535_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12845_  (.A(\reg_module/_05091_ ),
    .X(\reg_module/_05536_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12846_  (.A(\reg_module/_05535_ ),
    .B(\reg_module/_05536_ ),
    .Y(\reg_module/_05537_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_12847_  (.A(\reg_module/_05059_ ),
    .X(\reg_module/_05538_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12848_  (.A(\reg_module/_05538_ ),
    .X(\reg_module/_05539_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12849_  (.A(\reg_module/_05528_ ),
    .B(\reg_module/_05537_ ),
    .C(\reg_module/_05539_ ),
    .Y(\reg_module/_05540_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12850_  (.A(\reg_module/_05224_ ),
    .B(\reg_module/gprf[678] ),
    .Y(\reg_module/_05541_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12851_  (.A(\reg_module/gprf[646] ),
    .B(net824),
    .Y(\reg_module/_05542_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12852_  (.A(\reg_module/_05541_ ),
    .B(net724),
    .C(\reg_module/_05542_ ),
    .Y(\reg_module/_05543_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12853_  (.A(\reg_module/_05149_ ),
    .B(\reg_module/gprf[742] ),
    .Y(\reg_module/_05544_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12854_  (.A(\reg_module/gprf[710] ),
    .B(net824),
    .Y(\reg_module/_05545_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12855_  (.A(\reg_module/_05544_ ),
    .B(\reg_module/_05464_ ),
    .C(\reg_module/_05545_ ),
    .Y(\reg_module/_05546_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12856_  (.A(\reg_module/_05543_ ),
    .B(\reg_module/_05546_ ),
    .Y(\reg_module/_05547_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12857_  (.A(\reg_module/_05547_ ),
    .B(\reg_module/_05011_ ),
    .Y(\reg_module/_05548_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12858_  (.A(\reg_module/_05315_ ),
    .B(\reg_module/gprf[550] ),
    .Y(\reg_module/_05549_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12859_  (.A(\reg_module/gprf[518] ),
    .B(net840),
    .Y(\reg_module/_05550_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12860_  (.A(\reg_module/_05549_ ),
    .B(net731),
    .C(\reg_module/_05550_ ),
    .Y(\reg_module/_05551_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12861_  (.A(\reg_module/_05472_ ),
    .B(\reg_module/gprf[614] ),
    .Y(\reg_module/_05552_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12862_  (.A(\reg_module/_05051_ ),
    .X(\reg_module/_05553_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12863_  (.A(\reg_module/gprf[582] ),
    .B(net841),
    .Y(\reg_module/_05554_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12864_  (.A(\reg_module/_05552_ ),
    .B(\reg_module/_05553_ ),
    .C(\reg_module/_05554_ ),
    .Y(\reg_module/_05555_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12865_  (.A(\reg_module/_05551_ ),
    .B(\reg_module/_05555_ ),
    .Y(\reg_module/_05556_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12866_  (.A(\reg_module/_05556_ ),
    .B(net675),
    .Y(\reg_module/_05557_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12867_  (.A(\reg_module/_05548_ ),
    .B(\reg_module/_05557_ ),
    .C(net650),
    .Y(\reg_module/_05558_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12868_  (.A(\reg_module/_05540_ ),
    .B(\reg_module/_05558_ ),
    .Y(\reg_module/_05559_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12869_  (.A(\reg_module/_05559_ ),
    .B(\reg_module/_05326_ ),
    .Y(\reg_module/_05560_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12870_  (.A(\reg_module/_05404_ ),
    .B(\reg_module/gprf[294] ),
    .Y(\reg_module/_05561_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12871_  (.A(\reg_module/gprf[262] ),
    .B(net835),
    .Y(\reg_module/_05562_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12872_  (.A(\reg_module/_05561_ ),
    .B(net729),
    .C(\reg_module/_05562_ ),
    .Y(\reg_module/_05563_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12873_  (.A(\reg_module/_05500_ ),
    .B(\reg_module/gprf[358] ),
    .Y(\reg_module/_05564_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12874_  (.A(\reg_module/gprf[326] ),
    .B(net836),
    .Y(\reg_module/_05565_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12875_  (.A(\reg_module/_05564_ ),
    .B(\reg_module/_05170_ ),
    .C(\reg_module/_05565_ ),
    .Y(\reg_module/_05566_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12876_  (.A(\reg_module/_05563_ ),
    .B(\reg_module/_05566_ ),
    .Y(\reg_module/_05567_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12877_  (.A(\reg_module/_05567_ ),
    .B(net674),
    .Y(\reg_module/_05568_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12878_  (.A(\reg_module/_05490_ ),
    .B(\reg_module/gprf[422] ),
    .Y(\reg_module/_05569_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12879_  (.A(\reg_module/gprf[390] ),
    .B(net821),
    .Y(\reg_module/_05570_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12880_  (.A(\reg_module/_05569_ ),
    .B(net722),
    .C(\reg_module/_05570_ ),
    .Y(\reg_module/_05571_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12881_  (.A(\reg_module/_05178_ ),
    .B(\reg_module/gprf[486] ),
    .Y(\reg_module/_05572_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12882_  (.A(\reg_module/gprf[454] ),
    .B(net820),
    .Y(\reg_module/_05573_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12883_  (.A(\reg_module/_05572_ ),
    .B(\reg_module/_05256_ ),
    .C(\reg_module/_05573_ ),
    .Y(\reg_module/_05574_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12884_  (.A(\reg_module/_05571_ ),
    .B(\reg_module/_05574_ ),
    .Y(\reg_module/_05575_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12885_  (.A(\reg_module/_05575_ ),
    .B(\reg_module/_05183_ ),
    .Y(\reg_module/_05576_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12886_  (.A(\reg_module/_05094_ ),
    .X(\reg_module/_05577_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12887_  (.A(\reg_module/_05568_ ),
    .B(\reg_module/_05576_ ),
    .C(\reg_module/_05577_ ),
    .Y(\reg_module/_05578_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12888_  (.A(\reg_module/_05500_ ),
    .B(\reg_module/gprf[38] ),
    .Y(\reg_module/_05579_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12889_  (.A(\reg_module/gprf[6] ),
    .B(net838),
    .Y(\reg_module/_05580_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12890_  (.A(\reg_module/_05579_ ),
    .B(net731),
    .C(\reg_module/_05580_ ),
    .Y(\reg_module/_05581_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12891_  (.A(\reg_module/_05504_ ),
    .B(\reg_module/gprf[102] ),
    .Y(\reg_module/_05582_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12892_  (.A(\reg_module/gprf[70] ),
    .B(net839),
    .Y(\reg_module/_05583_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12893_  (.A(\reg_module/_05582_ ),
    .B(\reg_module/_05426_ ),
    .C(\reg_module/_05583_ ),
    .Y(\reg_module/_05584_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12894_  (.A(\reg_module/_05581_ ),
    .B(\reg_module/_05584_ ),
    .Y(\reg_module/_05585_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12895_  (.A(\reg_module/_05585_ ),
    .B(net675),
    .Y(\reg_module/_05586_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12896_  (.A(\reg_module/_05353_ ),
    .B(\reg_module/gprf[166] ),
    .Y(\reg_module/_05587_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12897_  (.A(\reg_module/gprf[134] ),
    .B(net834),
    .Y(\reg_module/_05588_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12898_  (.A(\reg_module/_05587_ ),
    .B(net728),
    .C(\reg_module/_05588_ ),
    .Y(\reg_module/_05589_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12899_  (.A(\reg_module/_05357_ ),
    .B(\reg_module/gprf[230] ),
    .Y(\reg_module/_05590_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12900_  (.A(\reg_module/gprf[198] ),
    .B(net833),
    .Y(\reg_module/_05591_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12901_  (.A(\reg_module/_05590_ ),
    .B(\reg_module/_05435_ ),
    .C(\reg_module/_05591_ ),
    .Y(\reg_module/_05592_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12902_  (.A(\reg_module/_05589_ ),
    .B(\reg_module/_05592_ ),
    .Y(\reg_module/_05593_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12903_  (.A(\reg_module/_05009_ ),
    .X(\reg_module/_05594_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12904_  (.A(\reg_module/_05593_ ),
    .B(\reg_module/_05594_ ),
    .Y(\reg_module/_05595_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12905_  (.A(\reg_module/_05586_ ),
    .B(\reg_module/_05595_ ),
    .C(net649),
    .Y(\reg_module/_05596_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12906_  (.A(\reg_module/_05578_ ),
    .B(\reg_module/_05596_ ),
    .Y(\reg_module/_05597_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12907_  (.A(\reg_module/_05597_ ),
    .B(net633),
    .Y(\reg_module/_05598_ ));
 sky130_fd_sc_hd__nand2_4 \reg_module/_12908_  (.A(\reg_module/_05560_ ),
    .B(\reg_module/_05598_ ),
    .Y(\wRs1Data[6] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12909_  (.A(\reg_module/_05283_ ),
    .B(\reg_module/gprf[807] ),
    .Y(\reg_module/_05599_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12910_  (.A(\reg_module/gprf[775] ),
    .B(net836),
    .Y(\reg_module/_05600_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12911_  (.A(\reg_module/_05599_ ),
    .B(net729),
    .C(\reg_module/_05600_ ),
    .Y(\reg_module/_05601_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12912_  (.A(\reg_module/_05288_ ),
    .B(\reg_module/gprf[871] ),
    .Y(\reg_module/_05602_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12913_  (.A(\reg_module/gprf[839] ),
    .B(net835),
    .Y(\reg_module/_05603_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12914_  (.A(\reg_module/_05602_ ),
    .B(\reg_module/_05291_ ),
    .C(\reg_module/_05603_ ),
    .Y(\reg_module/_05604_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12915_  (.A(\reg_module/_05601_ ),
    .B(\reg_module/_05604_ ),
    .Y(\reg_module/_05605_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12916_  (.A(\reg_module/_05605_ ),
    .B(net674),
    .Y(\reg_module/_05606_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12917_  (.A(\reg_module/_05013_ ),
    .X(\reg_module/_05607_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12918_  (.A(\reg_module/_05607_ ),
    .B(\reg_module/gprf[935] ),
    .Y(\reg_module/_05608_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12919_  (.A(\reg_module/gprf[903] ),
    .B(net826),
    .Y(\reg_module/_05609_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12920_  (.A(\reg_module/_05608_ ),
    .B(net725),
    .C(\reg_module/_05609_ ),
    .Y(\reg_module/_05610_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12921_  (.A(\reg_module/_05019_ ),
    .X(\reg_module/_05611_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12922_  (.A(\reg_module/_05611_ ),
    .B(\reg_module/gprf[999] ),
    .Y(\reg_module/_05612_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12923_  (.A(\reg_module/gprf[967] ),
    .B(net826),
    .Y(\reg_module/_05613_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12924_  (.A(\reg_module/_05612_ ),
    .B(\reg_module/_05300_ ),
    .C(\reg_module/_05613_ ),
    .Y(\reg_module/_05614_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12925_  (.A(\reg_module/_05610_ ),
    .B(\reg_module/_05614_ ),
    .Y(\reg_module/_05615_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12926_  (.A(\reg_module/_05615_ ),
    .B(\reg_module/_05536_ ),
    .Y(\reg_module/_05616_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12927_  (.A(\reg_module/_05606_ ),
    .B(\reg_module/_05616_ ),
    .C(\reg_module/_05539_ ),
    .Y(\reg_module/_05617_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12928_  (.A(\reg_module/_05224_ ),
    .B(\reg_module/gprf[679] ),
    .Y(\reg_module/_05618_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12929_  (.A(\reg_module/gprf[647] ),
    .B(net824),
    .Y(\reg_module/_05619_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12930_  (.A(\reg_module/_05618_ ),
    .B(net724),
    .C(\reg_module/_05619_ ),
    .Y(\reg_module/_05620_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12931_  (.A(\reg_module/_05078_ ),
    .X(\reg_module/_05621_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12932_  (.A(\reg_module/_05621_ ),
    .B(\reg_module/gprf[743] ),
    .Y(\reg_module/_05622_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12933_  (.A(\reg_module/gprf[711] ),
    .B(net825),
    .Y(\reg_module/_05623_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12934_  (.A(\reg_module/_05622_ ),
    .B(\reg_module/_05464_ ),
    .C(\reg_module/_05623_ ),
    .Y(\reg_module/_05624_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12935_  (.A(\reg_module/_05620_ ),
    .B(\reg_module/_05624_ ),
    .Y(\reg_module/_05625_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12936_  (.A(\reg_module/_05625_ ),
    .B(\reg_module/_05011_ ),
    .Y(\reg_module/_05626_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12937_  (.A(\reg_module/_05315_ ),
    .B(\reg_module/gprf[551] ),
    .Y(\reg_module/_05627_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12938_  (.A(\reg_module/gprf[519] ),
    .B(net841),
    .Y(\reg_module/_05628_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12939_  (.A(\reg_module/_05627_ ),
    .B(net731),
    .C(\reg_module/_05628_ ),
    .Y(\reg_module/_05629_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12940_  (.A(\reg_module/_05472_ ),
    .B(\reg_module/gprf[615] ),
    .Y(\reg_module/_05630_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12941_  (.A(\reg_module/gprf[583] ),
    .B(net840),
    .Y(\reg_module/_05631_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12942_  (.A(\reg_module/_05630_ ),
    .B(\reg_module/_05553_ ),
    .C(\reg_module/_05631_ ),
    .Y(\reg_module/_05632_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12943_  (.A(\reg_module/_05629_ ),
    .B(\reg_module/_05632_ ),
    .Y(\reg_module/_05633_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12944_  (.A(\reg_module/_05633_ ),
    .B(net677),
    .Y(\reg_module/_05634_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12945_  (.A(\reg_module/_05626_ ),
    .B(\reg_module/_05634_ ),
    .C(net648),
    .Y(\reg_module/_05635_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12946_  (.A(\reg_module/_05617_ ),
    .B(\reg_module/_05635_ ),
    .Y(\reg_module/_05636_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12947_  (.A(\reg_module/_05636_ ),
    .B(\reg_module/_05326_ ),
    .Y(\reg_module/_05637_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12948_  (.A(\reg_module/_05404_ ),
    .B(\reg_module/gprf[295] ),
    .Y(\reg_module/_05638_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12949_  (.A(\reg_module/gprf[263] ),
    .B(net835),
    .Y(\reg_module/_05639_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12950_  (.A(\reg_module/_05638_ ),
    .B(net729),
    .C(\reg_module/_05639_ ),
    .Y(\reg_module/_05640_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12951_  (.A(\reg_module/_05500_ ),
    .B(\reg_module/gprf[359] ),
    .Y(\reg_module/_05641_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12952_  (.A(\reg_module/_05072_ ),
    .X(\reg_module/_05642_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12953_  (.A(\reg_module/gprf[327] ),
    .B(net835),
    .Y(\reg_module/_05643_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12954_  (.A(\reg_module/_05641_ ),
    .B(\reg_module/_05642_ ),
    .C(\reg_module/_05643_ ),
    .Y(\reg_module/_05644_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12955_  (.A(\reg_module/_05640_ ),
    .B(\reg_module/_05644_ ),
    .Y(\reg_module/_05645_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12956_  (.A(\reg_module/_05645_ ),
    .B(net675),
    .Y(\reg_module/_05646_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12957_  (.A(\reg_module/_05490_ ),
    .B(\reg_module/gprf[423] ),
    .Y(\reg_module/_05647_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12958_  (.A(\reg_module/gprf[391] ),
    .B(net822),
    .Y(\reg_module/_05648_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12959_  (.A(\reg_module/_05647_ ),
    .B(net723),
    .C(\reg_module/_05648_ ),
    .Y(\reg_module/_05649_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_12960_  (.A(\reg_module/_05083_ ),
    .X(\reg_module/_05650_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12961_  (.A(\reg_module/_05650_ ),
    .B(\reg_module/gprf[487] ),
    .Y(\reg_module/_05651_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12962_  (.A(\reg_module/gprf[455] ),
    .B(net823),
    .Y(\reg_module/_05652_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12963_  (.A(\reg_module/_05651_ ),
    .B(\reg_module/_05256_ ),
    .C(\reg_module/_05652_ ),
    .Y(\reg_module/_05653_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12964_  (.A(\reg_module/_05649_ ),
    .B(\reg_module/_05653_ ),
    .Y(\reg_module/_05654_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_12965_  (.A(\reg_module/_05056_ ),
    .X(\reg_module/_05655_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12966_  (.A(\reg_module/_05654_ ),
    .B(\reg_module/_05655_ ),
    .Y(\reg_module/_05656_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12967_  (.A(\reg_module/_05646_ ),
    .B(\reg_module/_05656_ ),
    .C(\reg_module/_05577_ ),
    .Y(\reg_module/_05657_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12968_  (.A(\reg_module/_05500_ ),
    .B(\reg_module/gprf[39] ),
    .Y(\reg_module/_05658_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12969_  (.A(\reg_module/gprf[7] ),
    .B(net840),
    .Y(\reg_module/_05659_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12970_  (.A(\reg_module/_05658_ ),
    .B(net732),
    .C(\reg_module/_05659_ ),
    .Y(\reg_module/_05660_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12971_  (.A(\reg_module/_05504_ ),
    .B(\reg_module/gprf[103] ),
    .Y(\reg_module/_05661_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12972_  (.A(\reg_module/gprf[71] ),
    .B(net840),
    .Y(\reg_module/_05662_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12973_  (.A(\reg_module/_05661_ ),
    .B(\reg_module/_05426_ ),
    .C(\reg_module/_05662_ ),
    .Y(\reg_module/_05663_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12974_  (.A(\reg_module/_05660_ ),
    .B(\reg_module/_05663_ ),
    .Y(\reg_module/_05664_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12975_  (.A(\reg_module/_05664_ ),
    .B(net675),
    .Y(\reg_module/_05665_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12976_  (.A(\reg_module/_05353_ ),
    .B(\reg_module/gprf[167] ),
    .Y(\reg_module/_05666_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12977_  (.A(\reg_module/gprf[135] ),
    .B(net833),
    .Y(\reg_module/_05667_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12978_  (.A(\reg_module/_05666_ ),
    .B(net728),
    .C(\reg_module/_05667_ ),
    .Y(\reg_module/_05668_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12979_  (.A(\reg_module/_05357_ ),
    .B(\reg_module/gprf[231] ),
    .Y(\reg_module/_05669_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12980_  (.A(\reg_module/gprf[199] ),
    .B(net833),
    .Y(\reg_module/_05670_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12981_  (.A(\reg_module/_05669_ ),
    .B(\reg_module/_05435_ ),
    .C(\reg_module/_05670_ ),
    .Y(\reg_module/_05671_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12982_  (.A(\reg_module/_05668_ ),
    .B(\reg_module/_05671_ ),
    .Y(\reg_module/_05672_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12983_  (.A(\reg_module/_05672_ ),
    .B(\reg_module/_05594_ ),
    .Y(\reg_module/_05673_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12984_  (.A(\reg_module/_05665_ ),
    .B(\reg_module/_05673_ ),
    .C(net649),
    .Y(\reg_module/_05674_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12985_  (.A(\reg_module/_05657_ ),
    .B(\reg_module/_05674_ ),
    .Y(\reg_module/_05675_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12986_  (.A(\reg_module/_05675_ ),
    .B(net634),
    .Y(\reg_module/_05676_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_12987_  (.A(\reg_module/_05637_ ),
    .B(\reg_module/_05676_ ),
    .Y(\wRs1Data[7] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12988_  (.A(\reg_module/_05283_ ),
    .B(\reg_module/gprf[552] ),
    .Y(\reg_module/_05677_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12989_  (.A(\reg_module/gprf[520] ),
    .B(net837),
    .Y(\reg_module/_05678_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12990_  (.A(\reg_module/_05677_ ),
    .B(net729),
    .C(\reg_module/_05678_ ),
    .Y(\reg_module/_05679_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12991_  (.A(\reg_module/_05288_ ),
    .B(\reg_module/gprf[616] ),
    .Y(\reg_module/_05680_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12992_  (.A(\reg_module/gprf[584] ),
    .B(net837),
    .Y(\reg_module/_05681_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12993_  (.A(\reg_module/_05680_ ),
    .B(\reg_module/_05291_ ),
    .C(\reg_module/_05681_ ),
    .Y(\reg_module/_05682_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12994_  (.A(\reg_module/_05679_ ),
    .B(\reg_module/_05682_ ),
    .Y(\reg_module/_05683_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12995_  (.A(\reg_module/_05683_ ),
    .B(net674),
    .Y(\reg_module/_05684_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12996_  (.A(\reg_module/_05607_ ),
    .B(\reg_module/gprf[680] ),
    .Y(\reg_module/_05685_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12997_  (.A(\reg_module/gprf[648] ),
    .B(net826),
    .Y(\reg_module/_05686_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_12998_  (.A(\reg_module/_05685_ ),
    .B(net725),
    .C(\reg_module/_05686_ ),
    .Y(\reg_module/_05687_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_12999_  (.A(\reg_module/_05611_ ),
    .B(\reg_module/gprf[744] ),
    .Y(\reg_module/_05688_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13000_  (.A(\reg_module/gprf[712] ),
    .B(net826),
    .Y(\reg_module/_05689_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13001_  (.A(\reg_module/_05688_ ),
    .B(\reg_module/_05300_ ),
    .C(\reg_module/_05689_ ),
    .Y(\reg_module/_05690_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13002_  (.A(\reg_module/_05687_ ),
    .B(\reg_module/_05690_ ),
    .Y(\reg_module/_05691_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13003_  (.A(\reg_module/_05691_ ),
    .B(\reg_module/_05536_ ),
    .Y(\reg_module/_05692_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13004_  (.A(\reg_module/_05684_ ),
    .B(\reg_module/_05692_ ),
    .C(net648),
    .Y(\reg_module/_05693_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13005_  (.A(\reg_module/_05029_ ),
    .X(\reg_module/_05694_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13006_  (.A(\reg_module/_05694_ ),
    .B(\reg_module/gprf[808] ),
    .Y(\reg_module/_05695_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13007_  (.A(\reg_module/gprf[776] ),
    .B(net837),
    .Y(\reg_module/_05696_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13008_  (.A(\reg_module/_05695_ ),
    .B(net730),
    .C(\reg_module/_05696_ ),
    .Y(\reg_module/_05697_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13009_  (.A(\reg_module/_05621_ ),
    .B(\reg_module/gprf[872] ),
    .Y(\reg_module/_05698_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13010_  (.A(\reg_module/gprf[840] ),
    .B(net826),
    .Y(\reg_module/_05699_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13011_  (.A(\reg_module/_05698_ ),
    .B(\reg_module/_05464_ ),
    .C(\reg_module/_05699_ ),
    .Y(\reg_module/_05700_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13012_  (.A(\reg_module/_05697_ ),
    .B(\reg_module/_05700_ ),
    .Y(\reg_module/_05701_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13013_  (.A(\reg_module/_05701_ ),
    .B(net673),
    .Y(\reg_module/_05702_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13014_  (.A(\reg_module/_05315_ ),
    .B(\reg_module/gprf[936] ),
    .Y(\reg_module/_05703_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13015_  (.A(\reg_module/gprf[904] ),
    .B(net827),
    .Y(\reg_module/_05704_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13016_  (.A(\reg_module/_05703_ ),
    .B(net725),
    .C(\reg_module/_05704_ ),
    .Y(\reg_module/_05705_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13017_  (.A(\reg_module/_05472_ ),
    .B(\reg_module/gprf[1000] ),
    .Y(\reg_module/_05706_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13018_  (.A(\reg_module/gprf[968] ),
    .B(net827),
    .Y(\reg_module/_05707_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13019_  (.A(\reg_module/_05706_ ),
    .B(\reg_module/_05553_ ),
    .C(\reg_module/_05707_ ),
    .Y(\reg_module/_05708_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13020_  (.A(\reg_module/_05705_ ),
    .B(\reg_module/_05708_ ),
    .Y(\reg_module/_05709_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13021_  (.A(\reg_module/_05709_ ),
    .B(\reg_module/_05477_ ),
    .Y(\reg_module/_05710_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13022_  (.A(\reg_module/_05702_ ),
    .B(\reg_module/_05710_ ),
    .C(\reg_module/_05400_ ),
    .Y(\reg_module/_05711_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13023_  (.A(\reg_module/_05693_ ),
    .B(\reg_module/_05711_ ),
    .Y(\reg_module/_05712_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13024_  (.A(\reg_module/_05712_ ),
    .B(\reg_module/_05326_ ),
    .Y(\reg_module/_05713_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13025_  (.A(\reg_module/_05404_ ),
    .B(\reg_module/gprf[296] ),
    .Y(\reg_module/_05714_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13026_  (.A(\reg_module/gprf[264] ),
    .B(net841),
    .Y(\reg_module/_05715_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13027_  (.A(\reg_module/_05714_ ),
    .B(net730),
    .C(\reg_module/_05715_ ),
    .Y(\reg_module/_05716_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13028_  (.A(\reg_module/_05500_ ),
    .B(\reg_module/gprf[360] ),
    .Y(\reg_module/_05717_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13029_  (.A(\reg_module/gprf[328] ),
    .B(net836),
    .Y(\reg_module/_05718_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13030_  (.A(\reg_module/_05717_ ),
    .B(\reg_module/_05642_ ),
    .C(\reg_module/_05718_ ),
    .Y(\reg_module/_05719_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13031_  (.A(\reg_module/_05716_ ),
    .B(\reg_module/_05719_ ),
    .Y(\reg_module/_05720_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13032_  (.A(\reg_module/_05720_ ),
    .B(net674),
    .Y(\reg_module/_05721_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13033_  (.A(\reg_module/_05490_ ),
    .B(\reg_module/gprf[424] ),
    .Y(\reg_module/_05722_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13034_  (.A(\reg_module/gprf[392] ),
    .B(net822),
    .Y(\reg_module/_05723_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13035_  (.A(\reg_module/_05722_ ),
    .B(net722),
    .C(\reg_module/_05723_ ),
    .Y(\reg_module/_05724_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13036_  (.A(\reg_module/_05650_ ),
    .B(\reg_module/gprf[488] ),
    .Y(\reg_module/_05725_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13037_  (.A(\reg_module/_05086_ ),
    .X(\reg_module/_05726_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13038_  (.A(\reg_module/gprf[456] ),
    .B(net822),
    .Y(\reg_module/_05727_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13039_  (.A(\reg_module/_05725_ ),
    .B(\reg_module/_05726_ ),
    .C(\reg_module/_05727_ ),
    .Y(\reg_module/_05728_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13040_  (.A(\reg_module/_05724_ ),
    .B(\reg_module/_05728_ ),
    .Y(\reg_module/_05729_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13041_  (.A(\reg_module/_05729_ ),
    .B(\reg_module/_05655_ ),
    .Y(\reg_module/_05730_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13042_  (.A(\reg_module/_05721_ ),
    .B(\reg_module/_05730_ ),
    .C(\reg_module/_05577_ ),
    .Y(\reg_module/_05731_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13043_  (.A(\reg_module/_05068_ ),
    .X(\reg_module/_05732_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13044_  (.A(\reg_module/_05732_ ),
    .B(\reg_module/gprf[40] ),
    .Y(\reg_module/_05733_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13045_  (.A(\reg_module/gprf[8] ),
    .B(net841),
    .Y(\reg_module/_05734_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13046_  (.A(\reg_module/_05733_ ),
    .B(net732),
    .C(\reg_module/_05734_ ),
    .Y(\reg_module/_05735_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13047_  (.A(\reg_module/_05504_ ),
    .B(\reg_module/gprf[104] ),
    .Y(\reg_module/_05736_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13048_  (.A(\reg_module/gprf[72] ),
    .B(net840),
    .Y(\reg_module/_05737_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13049_  (.A(\reg_module/_05736_ ),
    .B(\reg_module/_05426_ ),
    .C(\reg_module/_05737_ ),
    .Y(\reg_module/_05738_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13050_  (.A(\reg_module/_05735_ ),
    .B(\reg_module/_05738_ ),
    .Y(\reg_module/_05739_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13051_  (.A(\reg_module/_05739_ ),
    .B(net675),
    .Y(\reg_module/_05740_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13052_  (.A(\reg_module/_05353_ ),
    .B(\reg_module/gprf[168] ),
    .Y(\reg_module/_05741_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13053_  (.A(\reg_module/gprf[136] ),
    .B(net833),
    .Y(\reg_module/_05742_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13054_  (.A(\reg_module/_05741_ ),
    .B(net728),
    .C(\reg_module/_05742_ ),
    .Y(\reg_module/_05743_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13055_  (.A(\reg_module/_05357_ ),
    .B(\reg_module/gprf[232] ),
    .Y(\reg_module/_05744_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13056_  (.A(\reg_module/gprf[200] ),
    .B(net833),
    .Y(\reg_module/_05745_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13057_  (.A(\reg_module/_05744_ ),
    .B(\reg_module/_05435_ ),
    .C(\reg_module/_05745_ ),
    .Y(\reg_module/_05746_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13058_  (.A(\reg_module/_05743_ ),
    .B(\reg_module/_05746_ ),
    .Y(\reg_module/_05747_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13059_  (.A(\reg_module/_05747_ ),
    .B(\reg_module/_05594_ ),
    .Y(\reg_module/_05748_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13060_  (.A(\reg_module/_05740_ ),
    .B(\reg_module/_05748_ ),
    .C(net649),
    .Y(\reg_module/_05749_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13061_  (.A(\reg_module/_05731_ ),
    .B(\reg_module/_05749_ ),
    .Y(\reg_module/_05750_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13062_  (.A(\reg_module/_05750_ ),
    .B(net634),
    .Y(\reg_module/_05751_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_13063_  (.A(\reg_module/_05713_ ),
    .B(\reg_module/_05751_ ),
    .Y(\wRs1Data[8] ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13064_  (.A(\reg_module/_05002_ ),
    .X(\reg_module/_05752_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13065_  (.A(\reg_module/_05752_ ),
    .B(\reg_module/gprf[809] ),
    .Y(\reg_module/_05753_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13066_  (.A(\reg_module/gprf[777] ),
    .B(net861),
    .Y(\reg_module/_05754_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13067_  (.A(\reg_module/_05753_ ),
    .B(net744),
    .C(\reg_module/_05754_ ),
    .Y(\reg_module/_05755_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13068_  (.A(\reg_module/_05287_ ),
    .X(\reg_module/_05756_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13069_  (.A(\reg_module/_05756_ ),
    .B(\reg_module/gprf[873] ),
    .Y(\reg_module/_05757_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13070_  (.A(\reg_module/_05290_ ),
    .X(\reg_module/_05758_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13071_  (.A(\reg_module/gprf[841] ),
    .B(net861),
    .Y(\reg_module/_05759_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13072_  (.A(\reg_module/_05757_ ),
    .B(\reg_module/_05758_ ),
    .C(\reg_module/_05759_ ),
    .Y(\reg_module/_05760_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13073_  (.A(\reg_module/_05755_ ),
    .B(\reg_module/_05760_ ),
    .Y(\reg_module/_05761_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13074_  (.A(\reg_module/_05761_ ),
    .B(net679),
    .Y(\reg_module/_05762_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13075_  (.A(\reg_module/_05607_ ),
    .B(\reg_module/gprf[937] ),
    .Y(\reg_module/_05763_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13076_  (.A(\reg_module/gprf[905] ),
    .B(net847),
    .Y(\reg_module/_05764_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13077_  (.A(\reg_module/_05763_ ),
    .B(net736),
    .C(\reg_module/_05764_ ),
    .Y(\reg_module/_05765_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13078_  (.A(\reg_module/_05611_ ),
    .B(\reg_module/gprf[1001] ),
    .Y(\reg_module/_05766_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13079_  (.A(\reg_module/_05022_ ),
    .X(\reg_module/_05767_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13080_  (.A(\reg_module/gprf[969] ),
    .B(net826),
    .Y(\reg_module/_05768_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13081_  (.A(\reg_module/_05766_ ),
    .B(\reg_module/_05767_ ),
    .C(\reg_module/_05768_ ),
    .Y(\reg_module/_05769_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13082_  (.A(\reg_module/_05765_ ),
    .B(\reg_module/_05769_ ),
    .Y(\reg_module/_05770_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13083_  (.A(\reg_module/_05770_ ),
    .B(\reg_module/_05536_ ),
    .Y(\reg_module/_05771_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13084_  (.A(\reg_module/_05762_ ),
    .B(\reg_module/_05771_ ),
    .C(\reg_module/_05539_ ),
    .Y(\reg_module/_05772_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13085_  (.A(\reg_module/_05694_ ),
    .B(\reg_module/gprf[681] ),
    .Y(\reg_module/_05773_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13086_  (.A(\reg_module/gprf[649] ),
    .B(net827),
    .Y(\reg_module/_05774_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13087_  (.A(\reg_module/_05773_ ),
    .B(net725),
    .C(\reg_module/_05774_ ),
    .Y(\reg_module/_05775_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13088_  (.A(\reg_module/_05621_ ),
    .B(\reg_module/gprf[745] ),
    .Y(\reg_module/_05776_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13089_  (.A(\reg_module/gprf[713] ),
    .B(net827),
    .Y(\reg_module/_05777_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13090_  (.A(\reg_module/_05776_ ),
    .B(\reg_module/_05464_ ),
    .C(\reg_module/_05777_ ),
    .Y(\reg_module/_05778_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13091_  (.A(\reg_module/_05775_ ),
    .B(\reg_module/_05778_ ),
    .Y(\reg_module/_05779_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13092_  (.A(\reg_module/_05779_ ),
    .B(\reg_module/_05011_ ),
    .Y(\reg_module/_05780_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13093_  (.A(\reg_module/_05019_ ),
    .X(\reg_module/_05781_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13094_  (.A(\reg_module/_05781_ ),
    .B(\reg_module/gprf[553] ),
    .Y(\reg_module/_05782_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13095_  (.A(\reg_module/gprf[521] ),
    .B(net865),
    .Y(\reg_module/_05783_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13096_  (.A(\reg_module/_05782_ ),
    .B(net745),
    .C(\reg_module/_05783_ ),
    .Y(\reg_module/_05784_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13097_  (.A(\reg_module/_05472_ ),
    .B(\reg_module/gprf[617] ),
    .Y(\reg_module/_05785_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13098_  (.A(\reg_module/gprf[585] ),
    .B(net865),
    .Y(\reg_module/_05786_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13099_  (.A(\reg_module/_05785_ ),
    .B(\reg_module/_05553_ ),
    .C(\reg_module/_05786_ ),
    .Y(\reg_module/_05787_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13100_  (.A(\reg_module/_05784_ ),
    .B(\reg_module/_05787_ ),
    .Y(\reg_module/_05788_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13101_  (.A(\reg_module/_05788_ ),
    .B(net680),
    .Y(\reg_module/_05789_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13102_  (.A(\reg_module/_05780_ ),
    .B(\reg_module/_05789_ ),
    .C(net652),
    .Y(\reg_module/_05790_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13103_  (.A(\reg_module/_05772_ ),
    .B(\reg_module/_05790_ ),
    .Y(\reg_module/_05791_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13104_  (.A(\reg_module/_05204_ ),
    .X(\reg_module/_05792_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13105_  (.A(\reg_module/_05791_ ),
    .B(\reg_module/_05792_ ),
    .Y(\reg_module/_05793_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13106_  (.A(\reg_module/_05404_ ),
    .B(\reg_module/gprf[297] ),
    .Y(\reg_module/_05794_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13107_  (.A(\reg_module/gprf[265] ),
    .B(net841),
    .Y(\reg_module/_05795_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13108_  (.A(\reg_module/_05794_ ),
    .B(net730),
    .C(\reg_module/_05795_ ),
    .Y(\reg_module/_05796_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13109_  (.A(\reg_module/_05732_ ),
    .B(\reg_module/gprf[361] ),
    .Y(\reg_module/_05797_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13110_  (.A(\reg_module/gprf[329] ),
    .B(net836),
    .Y(\reg_module/_05798_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13111_  (.A(\reg_module/_05797_ ),
    .B(\reg_module/_05642_ ),
    .C(\reg_module/_05798_ ),
    .Y(\reg_module/_05799_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13112_  (.A(\reg_module/_05796_ ),
    .B(\reg_module/_05799_ ),
    .Y(\reg_module/_05800_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13113_  (.A(\reg_module/_05800_ ),
    .B(net674),
    .Y(\reg_module/_05801_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13114_  (.A(\reg_module/_05490_ ),
    .B(\reg_module/gprf[425] ),
    .Y(\reg_module/_05802_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13115_  (.A(\reg_module/gprf[393] ),
    .B(net822),
    .Y(\reg_module/_05803_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13116_  (.A(\reg_module/_05802_ ),
    .B(net723),
    .C(\reg_module/_05803_ ),
    .Y(\reg_module/_05804_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13117_  (.A(\reg_module/_05650_ ),
    .B(\reg_module/gprf[489] ),
    .Y(\reg_module/_05805_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13118_  (.A(\reg_module/gprf[457] ),
    .B(net822),
    .Y(\reg_module/_05806_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13119_  (.A(\reg_module/_05805_ ),
    .B(\reg_module/_05726_ ),
    .C(\reg_module/_05806_ ),
    .Y(\reg_module/_05807_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13120_  (.A(\reg_module/_05804_ ),
    .B(\reg_module/_05807_ ),
    .Y(\reg_module/_05808_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13121_  (.A(\reg_module/_05808_ ),
    .B(\reg_module/_05655_ ),
    .Y(\reg_module/_05809_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13122_  (.A(\reg_module/_05801_ ),
    .B(\reg_module/_05809_ ),
    .C(\reg_module/_05577_ ),
    .Y(\reg_module/_05810_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13123_  (.A(\reg_module/_05732_ ),
    .B(\reg_module/gprf[41] ),
    .Y(\reg_module/_05811_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13124_  (.A(\reg_module/gprf[9] ),
    .B(net842),
    .Y(\reg_module/_05812_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13125_  (.A(\reg_module/_05811_ ),
    .B(net732),
    .C(\reg_module/_05812_ ),
    .Y(\reg_module/_05813_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13126_  (.A(\reg_module/_05504_ ),
    .B(\reg_module/gprf[105] ),
    .Y(\reg_module/_05814_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13127_  (.A(\reg_module/gprf[73] ),
    .B(net840),
    .Y(\reg_module/_05815_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13128_  (.A(\reg_module/_05814_ ),
    .B(\reg_module/_05426_ ),
    .C(\reg_module/_05815_ ),
    .Y(\reg_module/_05816_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13129_  (.A(\reg_module/_05813_ ),
    .B(\reg_module/_05816_ ),
    .Y(\reg_module/_05817_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13130_  (.A(\reg_module/_05817_ ),
    .B(net677),
    .Y(\reg_module/_05818_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13131_  (.A(\reg_module/_05108_ ),
    .X(\reg_module/_05819_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13132_  (.A(\reg_module/_05819_ ),
    .B(\reg_module/gprf[169] ),
    .Y(\reg_module/_05820_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13133_  (.A(\reg_module/gprf[137] ),
    .B(net838),
    .Y(\reg_module/_05821_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13134_  (.A(\reg_module/_05820_ ),
    .B(net731),
    .C(\reg_module/_05821_ ),
    .Y(\reg_module/_05822_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13135_  (.A(\reg_module/_05113_ ),
    .X(\reg_module/_05823_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13136_  (.A(\reg_module/_05823_ ),
    .B(\reg_module/gprf[233] ),
    .Y(\reg_module/_05824_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13137_  (.A(\reg_module/gprf[201] ),
    .B(net838),
    .Y(\reg_module/_05825_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13138_  (.A(\reg_module/_05824_ ),
    .B(\reg_module/_05435_ ),
    .C(\reg_module/_05825_ ),
    .Y(\reg_module/_05826_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13139_  (.A(\reg_module/_05822_ ),
    .B(\reg_module/_05826_ ),
    .Y(\reg_module/_05827_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13140_  (.A(\reg_module/_05827_ ),
    .B(\reg_module/_05594_ ),
    .Y(\reg_module/_05828_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13141_  (.A(\reg_module/_05818_ ),
    .B(\reg_module/_05828_ ),
    .C(net649),
    .Y(\reg_module/_05829_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13142_  (.A(\reg_module/_05810_ ),
    .B(\reg_module/_05829_ ),
    .Y(\reg_module/_05830_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13143_  (.A(\reg_module/_05830_ ),
    .B(net634),
    .Y(\reg_module/_05831_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_13144_  (.A(\reg_module/_05793_ ),
    .B(\reg_module/_05831_ ),
    .Y(\wRs1Data[9] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13145_  (.A(\reg_module/_05752_ ),
    .B(\reg_module/gprf[810] ),
    .Y(\reg_module/_05832_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13146_  (.A(\reg_module/gprf[778] ),
    .B(net861),
    .Y(\reg_module/_05833_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13147_  (.A(\reg_module/_05832_ ),
    .B(net744),
    .C(\reg_module/_05833_ ),
    .Y(\reg_module/_05834_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13148_  (.A(\reg_module/_05756_ ),
    .B(\reg_module/gprf[874] ),
    .Y(\reg_module/_05835_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13149_  (.A(\reg_module/gprf[842] ),
    .B(net861),
    .Y(\reg_module/_05836_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13150_  (.A(\reg_module/_05835_ ),
    .B(\reg_module/_05758_ ),
    .C(\reg_module/_05836_ ),
    .Y(\reg_module/_05837_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13151_  (.A(\reg_module/_05834_ ),
    .B(\reg_module/_05837_ ),
    .Y(\reg_module/_05838_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13152_  (.A(\reg_module/_05838_ ),
    .B(net679),
    .Y(\reg_module/_05839_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13153_  (.A(\reg_module/_05607_ ),
    .B(\reg_module/gprf[938] ),
    .Y(\reg_module/_05840_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13154_  (.A(\reg_module/gprf[906] ),
    .B(net847),
    .Y(\reg_module/_05841_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13155_  (.A(\reg_module/_05840_ ),
    .B(net736),
    .C(\reg_module/_05841_ ),
    .Y(\reg_module/_05842_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13156_  (.A(\reg_module/_05611_ ),
    .B(\reg_module/gprf[1002] ),
    .Y(\reg_module/_05843_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13157_  (.A(\reg_module/gprf[970] ),
    .B(net847),
    .Y(\reg_module/_05844_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13158_  (.A(\reg_module/_05843_ ),
    .B(\reg_module/_05767_ ),
    .C(\reg_module/_05844_ ),
    .Y(\reg_module/_05845_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13159_  (.A(\reg_module/_05842_ ),
    .B(\reg_module/_05845_ ),
    .Y(\reg_module/_05846_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13160_  (.A(\reg_module/_05846_ ),
    .B(\reg_module/_05536_ ),
    .Y(\reg_module/_05847_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13161_  (.A(\reg_module/_05839_ ),
    .B(\reg_module/_05847_ ),
    .C(\reg_module/_05539_ ),
    .Y(\reg_module/_05848_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13162_  (.A(\reg_module/_05694_ ),
    .B(\reg_module/gprf[682] ),
    .Y(\reg_module/_05849_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13163_  (.A(\reg_module/gprf[650] ),
    .B(net861),
    .Y(\reg_module/_05850_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13164_  (.A(\reg_module/_05849_ ),
    .B(net744),
    .C(\reg_module/_05850_ ),
    .Y(\reg_module/_05851_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13165_  (.A(\reg_module/_05621_ ),
    .B(\reg_module/gprf[746] ),
    .Y(\reg_module/_05852_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13166_  (.A(\reg_module/gprf[714] ),
    .B(net847),
    .Y(\reg_module/_05853_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13167_  (.A(\reg_module/_05852_ ),
    .B(\reg_module/_05464_ ),
    .C(\reg_module/_05853_ ),
    .Y(\reg_module/_05854_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13168_  (.A(\reg_module/_05851_ ),
    .B(\reg_module/_05854_ ),
    .Y(\reg_module/_05855_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13169_  (.A(\reg_module/_05010_ ),
    .X(\reg_module/_05856_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13170_  (.A(\reg_module/_05855_ ),
    .B(\reg_module/_05856_ ),
    .Y(\reg_module/_05857_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13171_  (.A(\reg_module/_05781_ ),
    .B(\reg_module/gprf[554] ),
    .Y(\reg_module/_05858_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13172_  (.A(\reg_module/gprf[522] ),
    .B(net865),
    .Y(\reg_module/_05859_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13173_  (.A(\reg_module/_05858_ ),
    .B(net745),
    .C(\reg_module/_05859_ ),
    .Y(\reg_module/_05860_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13174_  (.A(\reg_module/_05472_ ),
    .B(\reg_module/gprf[618] ),
    .Y(\reg_module/_05861_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13175_  (.A(\reg_module/gprf[586] ),
    .B(net866),
    .Y(\reg_module/_05862_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13176_  (.A(\reg_module/_05861_ ),
    .B(\reg_module/_05553_ ),
    .C(\reg_module/_05862_ ),
    .Y(\reg_module/_05863_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13177_  (.A(\reg_module/_05860_ ),
    .B(\reg_module/_05863_ ),
    .Y(\reg_module/_05864_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13178_  (.A(\reg_module/_05864_ ),
    .B(net680),
    .Y(\reg_module/_05865_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13179_  (.A(\reg_module/_05857_ ),
    .B(\reg_module/_05865_ ),
    .C(net652),
    .Y(\reg_module/_05866_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13180_  (.A(\reg_module/_05848_ ),
    .B(\reg_module/_05866_ ),
    .Y(\reg_module/_05867_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13181_  (.A(\reg_module/_05867_ ),
    .B(\reg_module/_05792_ ),
    .Y(\reg_module/_05868_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13182_  (.A(\reg_module/_05029_ ),
    .X(\reg_module/_05869_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13183_  (.A(\reg_module/_05869_ ),
    .B(\reg_module/gprf[298] ),
    .Y(\reg_module/_05870_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13184_  (.A(\reg_module/gprf[266] ),
    .B(net864),
    .Y(\reg_module/_05871_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13185_  (.A(\reg_module/_05870_ ),
    .B(net746),
    .C(\reg_module/_05871_ ),
    .Y(\reg_module/_05872_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13186_  (.A(\reg_module/_05732_ ),
    .B(\reg_module/gprf[362] ),
    .Y(\reg_module/_05873_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13187_  (.A(\reg_module/gprf[330] ),
    .B(net864),
    .Y(\reg_module/_05874_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13188_  (.A(\reg_module/_05873_ ),
    .B(\reg_module/_05642_ ),
    .C(\reg_module/_05874_ ),
    .Y(\reg_module/_05875_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13189_  (.A(\reg_module/_05872_ ),
    .B(\reg_module/_05875_ ),
    .Y(\reg_module/_05876_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13190_  (.A(\reg_module/_05876_ ),
    .B(net679),
    .Y(\reg_module/_05877_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13191_  (.A(\reg_module/_05490_ ),
    .B(\reg_module/gprf[426] ),
    .Y(\reg_module/_05878_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13192_  (.A(\reg_module/gprf[394] ),
    .B(net846),
    .Y(\reg_module/_05879_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13193_  (.A(\reg_module/_05878_ ),
    .B(net735),
    .C(\reg_module/_05879_ ),
    .Y(\reg_module/_05880_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13194_  (.A(\reg_module/_05650_ ),
    .B(\reg_module/gprf[490] ),
    .Y(\reg_module/_05881_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13195_  (.A(\reg_module/gprf[458] ),
    .B(net845),
    .Y(\reg_module/_05882_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13196_  (.A(\reg_module/_05881_ ),
    .B(\reg_module/_05726_ ),
    .C(\reg_module/_05882_ ),
    .Y(\reg_module/_05883_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13197_  (.A(\reg_module/_05880_ ),
    .B(\reg_module/_05883_ ),
    .Y(\reg_module/_05884_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13198_  (.A(\reg_module/_05884_ ),
    .B(\reg_module/_05655_ ),
    .Y(\reg_module/_05885_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13199_  (.A(\reg_module/_05877_ ),
    .B(\reg_module/_05885_ ),
    .C(\reg_module/_05577_ ),
    .Y(\reg_module/_05886_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13200_  (.A(\reg_module/_05732_ ),
    .B(\reg_module/gprf[42] ),
    .Y(\reg_module/_05887_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13201_  (.A(\reg_module/gprf[10] ),
    .B(net865),
    .Y(\reg_module/_05888_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13202_  (.A(\reg_module/_05887_ ),
    .B(net745),
    .C(\reg_module/_05888_ ),
    .Y(\reg_module/_05889_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13203_  (.A(\reg_module/_05504_ ),
    .B(\reg_module/gprf[106] ),
    .Y(\reg_module/_05890_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13204_  (.A(\reg_module/_04997_ ),
    .X(\reg_module/_05891_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13205_  (.A(\reg_module/gprf[74] ),
    .B(net866),
    .Y(\reg_module/_05892_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13206_  (.A(\reg_module/_05890_ ),
    .B(\reg_module/_05891_ ),
    .C(\reg_module/_05892_ ),
    .Y(\reg_module/_05893_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13207_  (.A(\reg_module/_05889_ ),
    .B(\reg_module/_05893_ ),
    .Y(\reg_module/_05894_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13208_  (.A(\reg_module/_05894_ ),
    .B(net680),
    .Y(\reg_module/_05895_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13209_  (.A(\reg_module/_05819_ ),
    .B(\reg_module/gprf[170] ),
    .Y(\reg_module/_05896_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13210_  (.A(\reg_module/gprf[138] ),
    .B(net838),
    .Y(\reg_module/_05897_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13211_  (.A(\reg_module/_05896_ ),
    .B(net731),
    .C(\reg_module/_05897_ ),
    .Y(\reg_module/_05898_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13212_  (.A(\reg_module/_05823_ ),
    .B(\reg_module/gprf[234] ),
    .Y(\reg_module/_05899_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13213_  (.A(\reg_module/_05071_ ),
    .X(\reg_module/_05900_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13214_  (.A(\reg_module/gprf[202] ),
    .B(net838),
    .Y(\reg_module/_05901_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13215_  (.A(\reg_module/_05899_ ),
    .B(\reg_module/_05900_ ),
    .C(\reg_module/_05901_ ),
    .Y(\reg_module/_05902_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13216_  (.A(\reg_module/_05898_ ),
    .B(\reg_module/_05902_ ),
    .Y(\reg_module/_05903_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13217_  (.A(\reg_module/_05903_ ),
    .B(\reg_module/_05594_ ),
    .Y(\reg_module/_05904_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13218_  (.A(\reg_module/_05895_ ),
    .B(\reg_module/_05904_ ),
    .C(net652),
    .Y(\reg_module/_05905_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13219_  (.A(\reg_module/_05886_ ),
    .B(\reg_module/_05905_ ),
    .Y(\reg_module/_05906_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13220_  (.A(\reg_module/_05906_ ),
    .B(net637),
    .Y(\reg_module/_05907_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_13221_  (.A(\reg_module/_05868_ ),
    .B(\reg_module/_05907_ ),
    .Y(\wRs1Data[10] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13222_  (.A(\reg_module/_05752_ ),
    .B(\reg_module/gprf[555] ),
    .Y(\reg_module/_05908_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13223_  (.A(\reg_module/gprf[523] ),
    .B(net862),
    .Y(\reg_module/_05909_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13224_  (.A(\reg_module/_05908_ ),
    .B(net744),
    .C(\reg_module/_05909_ ),
    .Y(\reg_module/_05910_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13225_  (.A(\reg_module/_05756_ ),
    .B(\reg_module/gprf[619] ),
    .Y(\reg_module/_05911_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13226_  (.A(\reg_module/gprf[587] ),
    .B(net862),
    .Y(\reg_module/_05912_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13227_  (.A(\reg_module/_05911_ ),
    .B(\reg_module/_05758_ ),
    .C(\reg_module/_05912_ ),
    .Y(\reg_module/_05913_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13228_  (.A(\reg_module/_05910_ ),
    .B(\reg_module/_05913_ ),
    .Y(\reg_module/_05914_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13229_  (.A(\reg_module/_05914_ ),
    .B(net679),
    .Y(\reg_module/_05915_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13230_  (.A(\reg_module/_05607_ ),
    .B(\reg_module/gprf[683] ),
    .Y(\reg_module/_05916_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13231_  (.A(\reg_module/gprf[651] ),
    .B(net847),
    .Y(\reg_module/_05917_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13232_  (.A(\reg_module/_05916_ ),
    .B(net736),
    .C(\reg_module/_05917_ ),
    .Y(\reg_module/_05918_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13233_  (.A(\reg_module/_05611_ ),
    .B(\reg_module/gprf[747] ),
    .Y(\reg_module/_05919_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13234_  (.A(\reg_module/gprf[715] ),
    .B(net847),
    .Y(\reg_module/_05920_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13235_  (.A(\reg_module/_05919_ ),
    .B(\reg_module/_05767_ ),
    .C(\reg_module/_05920_ ),
    .Y(\reg_module/_05921_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13236_  (.A(\reg_module/_05918_ ),
    .B(\reg_module/_05921_ ),
    .Y(\reg_module/_05922_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13237_  (.A(\reg_module/_05922_ ),
    .B(\reg_module/_05536_ ),
    .Y(\reg_module/_05923_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13238_  (.A(\reg_module/_05915_ ),
    .B(\reg_module/_05923_ ),
    .C(net653),
    .Y(\reg_module/_05924_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13239_  (.A(\reg_module/_05694_ ),
    .B(\reg_module/gprf[811] ),
    .Y(\reg_module/_05925_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13240_  (.A(\reg_module/gprf[779] ),
    .B(net861),
    .Y(\reg_module/_05926_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13241_  (.A(\reg_module/_05925_ ),
    .B(net744),
    .C(\reg_module/_05926_ ),
    .Y(\reg_module/_05927_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13242_  (.A(\reg_module/_05621_ ),
    .B(\reg_module/gprf[875] ),
    .Y(\reg_module/_05928_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13243_  (.A(\reg_module/_05037_ ),
    .X(\reg_module/_05929_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13244_  (.A(\reg_module/gprf[843] ),
    .B(net862),
    .Y(\reg_module/_05930_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13245_  (.A(\reg_module/_05928_ ),
    .B(\reg_module/_05929_ ),
    .C(\reg_module/_05930_ ),
    .Y(\reg_module/_05931_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13246_  (.A(\reg_module/_05927_ ),
    .B(\reg_module/_05931_ ),
    .Y(\reg_module/_05932_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13247_  (.A(\reg_module/_05932_ ),
    .B(net679),
    .Y(\reg_module/_05933_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13248_  (.A(\reg_module/_05781_ ),
    .B(\reg_module/gprf[939] ),
    .Y(\reg_module/_05934_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13249_  (.A(\reg_module/gprf[907] ),
    .B(net850),
    .Y(\reg_module/_05935_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13250_  (.A(\reg_module/_05934_ ),
    .B(net736),
    .C(\reg_module/_05935_ ),
    .Y(\reg_module/_05936_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13251_  (.A(\reg_module/_05048_ ),
    .X(\reg_module/_05937_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13252_  (.A(\reg_module/_05937_ ),
    .B(\reg_module/gprf[1003] ),
    .Y(\reg_module/_05938_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13253_  (.A(\reg_module/gprf[971] ),
    .B(net850),
    .Y(\reg_module/_05939_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13254_  (.A(\reg_module/_05938_ ),
    .B(\reg_module/_05553_ ),
    .C(\reg_module/_05939_ ),
    .Y(\reg_module/_05940_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13255_  (.A(\reg_module/_05936_ ),
    .B(\reg_module/_05940_ ),
    .Y(\reg_module/_05941_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13256_  (.A(\reg_module/_05941_ ),
    .B(\reg_module/_05477_ ),
    .Y(\reg_module/_05942_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13257_  (.A(\reg_module/_05933_ ),
    .B(\reg_module/_05942_ ),
    .C(\reg_module/_05400_ ),
    .Y(\reg_module/_05943_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13258_  (.A(\reg_module/_05924_ ),
    .B(\reg_module/_05943_ ),
    .Y(\reg_module/_05944_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13259_  (.A(\reg_module/_05944_ ),
    .B(\reg_module/_05792_ ),
    .Y(\reg_module/_05945_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13260_  (.A(\reg_module/_05869_ ),
    .B(\reg_module/gprf[299] ),
    .Y(\reg_module/_05946_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13261_  (.A(\reg_module/gprf[267] ),
    .B(net863),
    .Y(\reg_module/_05947_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13262_  (.A(\reg_module/_05946_ ),
    .B(net744),
    .C(\reg_module/_05947_ ),
    .Y(\reg_module/_05948_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13263_  (.A(\reg_module/_05732_ ),
    .B(\reg_module/gprf[363] ),
    .Y(\reg_module/_05949_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13264_  (.A(\reg_module/gprf[331] ),
    .B(net863),
    .Y(\reg_module/_05950_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13265_  (.A(\reg_module/_05949_ ),
    .B(\reg_module/_05642_ ),
    .C(\reg_module/_05950_ ),
    .Y(\reg_module/_05951_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13266_  (.A(\reg_module/_05948_ ),
    .B(\reg_module/_05951_ ),
    .Y(\reg_module/_05952_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13267_  (.A(\reg_module/_05952_ ),
    .B(net679),
    .Y(\reg_module/_05953_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13268_  (.A(\reg_module/_05043_ ),
    .X(\reg_module/_05954_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13269_  (.A(\reg_module/_05954_ ),
    .B(\reg_module/gprf[427] ),
    .Y(\reg_module/_05955_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13270_  (.A(\reg_module/gprf[395] ),
    .B(net845),
    .Y(\reg_module/_05956_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13271_  (.A(\reg_module/_05955_ ),
    .B(net735),
    .C(\reg_module/_05956_ ),
    .Y(\reg_module/_05957_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13272_  (.A(\reg_module/_05650_ ),
    .B(\reg_module/gprf[491] ),
    .Y(\reg_module/_05958_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13273_  (.A(\reg_module/gprf[459] ),
    .B(net845),
    .Y(\reg_module/_05959_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13274_  (.A(\reg_module/_05958_ ),
    .B(\reg_module/_05726_ ),
    .C(\reg_module/_05959_ ),
    .Y(\reg_module/_05960_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13275_  (.A(\reg_module/_05957_ ),
    .B(\reg_module/_05960_ ),
    .Y(\reg_module/_05961_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13276_  (.A(\reg_module/_05961_ ),
    .B(\reg_module/_05655_ ),
    .Y(\reg_module/_05962_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13277_  (.A(\reg_module/_05953_ ),
    .B(\reg_module/_05962_ ),
    .C(\reg_module/_05577_ ),
    .Y(\reg_module/_05963_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13278_  (.A(\reg_module/_05068_ ),
    .X(\reg_module/_05964_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13279_  (.A(\reg_module/_05964_ ),
    .B(\reg_module/gprf[43] ),
    .Y(\reg_module/_05965_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13280_  (.A(\reg_module/gprf[11] ),
    .B(net865),
    .Y(\reg_module/_05966_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13281_  (.A(\reg_module/_05965_ ),
    .B(net745),
    .C(\reg_module/_05966_ ),
    .Y(\reg_module/_05967_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13282_  (.A(\reg_module/_05100_ ),
    .X(\reg_module/_05968_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13283_  (.A(\reg_module/_05968_ ),
    .B(\reg_module/gprf[107] ),
    .Y(\reg_module/_05969_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13284_  (.A(\reg_module/gprf[75] ),
    .B(net866),
    .Y(\reg_module/_05970_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13285_  (.A(\reg_module/_05969_ ),
    .B(\reg_module/_05891_ ),
    .C(\reg_module/_05970_ ),
    .Y(\reg_module/_05971_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13286_  (.A(\reg_module/_05967_ ),
    .B(\reg_module/_05971_ ),
    .Y(\reg_module/_05972_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13287_  (.A(\reg_module/_05972_ ),
    .B(net680),
    .Y(\reg_module/_05973_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13288_  (.A(\reg_module/_05819_ ),
    .B(\reg_module/gprf[171] ),
    .Y(\reg_module/_05974_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13289_  (.A(\reg_module/gprf[139] ),
    .B(net838),
    .Y(\reg_module/_05975_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13290_  (.A(\reg_module/_05974_ ),
    .B(net731),
    .C(\reg_module/_05975_ ),
    .Y(\reg_module/_05976_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13291_  (.A(\reg_module/_05823_ ),
    .B(\reg_module/gprf[235] ),
    .Y(\reg_module/_05977_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13292_  (.A(\reg_module/gprf[203] ),
    .B(net839),
    .Y(\reg_module/_05978_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13293_  (.A(\reg_module/_05977_ ),
    .B(\reg_module/_05900_ ),
    .C(\reg_module/_05978_ ),
    .Y(\reg_module/_05979_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13294_  (.A(\reg_module/_05976_ ),
    .B(\reg_module/_05979_ ),
    .Y(\reg_module/_05980_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13295_  (.A(\reg_module/_05980_ ),
    .B(\reg_module/_05594_ ),
    .Y(\reg_module/_05981_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13296_  (.A(\reg_module/_05973_ ),
    .B(\reg_module/_05981_ ),
    .C(net652),
    .Y(\reg_module/_05982_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13297_  (.A(\reg_module/_05963_ ),
    .B(\reg_module/_05982_ ),
    .Y(\reg_module/_05983_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13298_  (.A(\reg_module/_05983_ ),
    .B(net637),
    .Y(\reg_module/_05984_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_13299_  (.A(\reg_module/_05945_ ),
    .B(\reg_module/_05984_ ),
    .Y(\wRs1Data[11] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13300_  (.A(\reg_module/_05752_ ),
    .B(\reg_module/gprf[812] ),
    .Y(\reg_module/_05985_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13301_  (.A(\reg_module/gprf[780] ),
    .B(net870),
    .Y(\reg_module/_05986_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13302_  (.A(\reg_module/_05985_ ),
    .B(net747),
    .C(\reg_module/_05986_ ),
    .Y(\reg_module/_05987_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13303_  (.A(\reg_module/_05756_ ),
    .B(\reg_module/gprf[876] ),
    .Y(\reg_module/_05988_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13304_  (.A(\reg_module/gprf[844] ),
    .B(net863),
    .Y(\reg_module/_05989_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13305_  (.A(\reg_module/_05988_ ),
    .B(\reg_module/_05758_ ),
    .C(\reg_module/_05989_ ),
    .Y(\reg_module/_05990_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13306_  (.A(\reg_module/_05987_ ),
    .B(\reg_module/_05990_ ),
    .Y(\reg_module/_05991_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13307_  (.A(\reg_module/_05991_ ),
    .B(net681),
    .Y(\reg_module/_05992_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13308_  (.A(\reg_module/_05607_ ),
    .B(\reg_module/gprf[940] ),
    .Y(\reg_module/_05993_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13309_  (.A(\reg_module/gprf[908] ),
    .B(net848),
    .Y(\reg_module/_05994_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13310_  (.A(\reg_module/_05993_ ),
    .B(net736),
    .C(\reg_module/_05994_ ),
    .Y(\reg_module/_05995_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13311_  (.A(\reg_module/_05611_ ),
    .B(\reg_module/gprf[1004] ),
    .Y(\reg_module/_05996_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13312_  (.A(\reg_module/gprf[972] ),
    .B(net848),
    .Y(\reg_module/_05997_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13313_  (.A(\reg_module/_05996_ ),
    .B(\reg_module/_05767_ ),
    .C(\reg_module/_05997_ ),
    .Y(\reg_module/_05998_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13314_  (.A(\reg_module/_05995_ ),
    .B(\reg_module/_05998_ ),
    .Y(\reg_module/_05999_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_13315_  (.A(\reg_module/_05091_ ),
    .X(\reg_module/_06000_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13316_  (.A(\reg_module/_05999_ ),
    .B(\reg_module/_06000_ ),
    .Y(\reg_module/_06001_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13317_  (.A(\reg_module/_05992_ ),
    .B(\reg_module/_06001_ ),
    .C(\reg_module/_05539_ ),
    .Y(\reg_module/_06002_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13318_  (.A(\reg_module/_05694_ ),
    .B(\reg_module/gprf[684] ),
    .Y(\reg_module/_06003_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13319_  (.A(\reg_module/gprf[652] ),
    .B(net849),
    .Y(\reg_module/_06004_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13320_  (.A(\reg_module/_06003_ ),
    .B(net737),
    .C(\reg_module/_06004_ ),
    .Y(\reg_module/_06005_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13321_  (.A(\reg_module/_05621_ ),
    .B(\reg_module/gprf[748] ),
    .Y(\reg_module/_06006_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13322_  (.A(\reg_module/gprf[716] ),
    .B(net849),
    .Y(\reg_module/_06007_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13323_  (.A(\reg_module/_06006_ ),
    .B(\reg_module/_05929_ ),
    .C(\reg_module/_06007_ ),
    .Y(\reg_module/_06008_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13324_  (.A(\reg_module/_06005_ ),
    .B(\reg_module/_06008_ ),
    .Y(\reg_module/_06009_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13325_  (.A(\reg_module/_06009_ ),
    .B(\reg_module/_05856_ ),
    .Y(\reg_module/_06010_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13326_  (.A(\reg_module/_05781_ ),
    .B(\reg_module/gprf[556] ),
    .Y(\reg_module/_06011_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13327_  (.A(\reg_module/gprf[524] ),
    .B(net874),
    .Y(\reg_module/_06012_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13328_  (.A(\reg_module/_06011_ ),
    .B(net749),
    .C(\reg_module/_06012_ ),
    .Y(\reg_module/_06013_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13329_  (.A(\reg_module/_05937_ ),
    .B(\reg_module/gprf[620] ),
    .Y(\reg_module/_06014_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13330_  (.A(\reg_module/_05051_ ),
    .X(\reg_module/_06015_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13331_  (.A(\reg_module/gprf[588] ),
    .B(net868),
    .Y(\reg_module/_06016_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13332_  (.A(\reg_module/_06014_ ),
    .B(\reg_module/_06015_ ),
    .C(\reg_module/_06016_ ),
    .Y(\reg_module/_06017_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13333_  (.A(\reg_module/_06013_ ),
    .B(\reg_module/_06017_ ),
    .Y(\reg_module/_06018_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13334_  (.A(\reg_module/_06018_ ),
    .B(net684),
    .Y(\reg_module/_06019_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13335_  (.A(\reg_module/_06010_ ),
    .B(\reg_module/_06019_ ),
    .C(net651),
    .Y(\reg_module/_06020_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13336_  (.A(\reg_module/_06002_ ),
    .B(\reg_module/_06020_ ),
    .Y(\reg_module/_06021_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13337_  (.A(\reg_module/_06021_ ),
    .B(\reg_module/_05792_ ),
    .Y(\reg_module/_06022_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13338_  (.A(\reg_module/_05869_ ),
    .B(\reg_module/gprf[300] ),
    .Y(\reg_module/_06023_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13339_  (.A(\reg_module/gprf[268] ),
    .B(net873),
    .Y(\reg_module/_06024_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13340_  (.A(\reg_module/_06023_ ),
    .B(net747),
    .C(\reg_module/_06024_ ),
    .Y(\reg_module/_06025_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13341_  (.A(\reg_module/_05964_ ),
    .B(\reg_module/gprf[364] ),
    .Y(\reg_module/_06026_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13342_  (.A(\reg_module/gprf[332] ),
    .B(net871),
    .Y(\reg_module/_06027_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13343_  (.A(\reg_module/_06026_ ),
    .B(\reg_module/_05642_ ),
    .C(\reg_module/_06027_ ),
    .Y(\reg_module/_06028_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13344_  (.A(\reg_module/_06025_ ),
    .B(\reg_module/_06028_ ),
    .Y(\reg_module/_06029_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13345_  (.A(\reg_module/_06029_ ),
    .B(net681),
    .Y(\reg_module/_06030_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13346_  (.A(\reg_module/_05954_ ),
    .B(\reg_module/gprf[428] ),
    .Y(\reg_module/_06031_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13347_  (.A(\reg_module/gprf[396] ),
    .B(net855),
    .Y(\reg_module/_06032_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13348_  (.A(\reg_module/_06031_ ),
    .B(net741),
    .C(\reg_module/_06032_ ),
    .Y(\reg_module/_06033_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13349_  (.A(\reg_module/_05650_ ),
    .B(\reg_module/gprf[492] ),
    .Y(\reg_module/_06034_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13350_  (.A(\reg_module/gprf[460] ),
    .B(net855),
    .Y(\reg_module/_06035_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13351_  (.A(\reg_module/_06034_ ),
    .B(\reg_module/_05726_ ),
    .C(\reg_module/_06035_ ),
    .Y(\reg_module/_06036_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13352_  (.A(\reg_module/_06033_ ),
    .B(\reg_module/_06036_ ),
    .Y(\reg_module/_06037_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13353_  (.A(\reg_module/_06037_ ),
    .B(\reg_module/_05655_ ),
    .Y(\reg_module/_06038_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13354_  (.A(\reg_module/_05094_ ),
    .X(\reg_module/_06039_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13355_  (.A(\reg_module/_06030_ ),
    .B(\reg_module/_06038_ ),
    .C(\reg_module/_06039_ ),
    .Y(\reg_module/_06040_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13356_  (.A(\reg_module/_05964_ ),
    .B(\reg_module/gprf[44] ),
    .Y(\reg_module/_06041_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13357_  (.A(\reg_module/gprf[12] ),
    .B(net875),
    .Y(\reg_module/_06042_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13358_  (.A(\reg_module/_06041_ ),
    .B(net749),
    .C(\reg_module/_06042_ ),
    .Y(\reg_module/_06043_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13359_  (.A(\reg_module/_05968_ ),
    .B(\reg_module/gprf[108] ),
    .Y(\reg_module/_06044_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13360_  (.A(\reg_module/gprf[76] ),
    .B(net875),
    .Y(\reg_module/_06045_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13361_  (.A(\reg_module/_06044_ ),
    .B(\reg_module/_05891_ ),
    .C(\reg_module/_06045_ ),
    .Y(\reg_module/_06046_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13362_  (.A(\reg_module/_06043_ ),
    .B(\reg_module/_06046_ ),
    .Y(\reg_module/_06047_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13363_  (.A(\reg_module/_06047_ ),
    .B(net684),
    .Y(\reg_module/_06048_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13364_  (.A(\reg_module/_05819_ ),
    .B(\reg_module/gprf[172] ),
    .Y(\reg_module/_06049_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13365_  (.A(\reg_module/gprf[140] ),
    .B(net867),
    .Y(\reg_module/_06050_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13366_  (.A(\reg_module/_06049_ ),
    .B(net746),
    .C(\reg_module/_06050_ ),
    .Y(\reg_module/_06051_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13367_  (.A(\reg_module/_05823_ ),
    .B(\reg_module/gprf[236] ),
    .Y(\reg_module/_06052_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13368_  (.A(\reg_module/gprf[204] ),
    .B(net867),
    .Y(\reg_module/_06053_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13369_  (.A(\reg_module/_06052_ ),
    .B(\reg_module/_05900_ ),
    .C(\reg_module/_06053_ ),
    .Y(\reg_module/_06054_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13370_  (.A(\reg_module/_06051_ ),
    .B(\reg_module/_06054_ ),
    .Y(\reg_module/_06055_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13371_  (.A(\reg_module/_05009_ ),
    .X(\reg_module/_06056_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13372_  (.A(\reg_module/_06055_ ),
    .B(\reg_module/_06056_ ),
    .Y(\reg_module/_06057_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13373_  (.A(\reg_module/_06048_ ),
    .B(\reg_module/_06057_ ),
    .C(net651),
    .Y(\reg_module/_06058_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13374_  (.A(\reg_module/_06040_ ),
    .B(\reg_module/_06058_ ),
    .Y(\reg_module/_06059_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13375_  (.A(\reg_module/_06059_ ),
    .B(net636),
    .Y(\reg_module/_06060_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_13376_  (.A(\reg_module/_06022_ ),
    .B(\reg_module/_06060_ ),
    .Y(\wRs1Data[12] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13377_  (.A(\reg_module/_05752_ ),
    .B(\reg_module/gprf[813] ),
    .Y(\reg_module/_06061_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13378_  (.A(\reg_module/gprf[781] ),
    .B(net870),
    .Y(\reg_module/_06062_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13379_  (.A(\reg_module/_06061_ ),
    .B(net747),
    .C(\reg_module/_06062_ ),
    .Y(\reg_module/_06063_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13380_  (.A(\reg_module/_05756_ ),
    .B(\reg_module/gprf[877] ),
    .Y(\reg_module/_06064_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13381_  (.A(\reg_module/gprf[845] ),
    .B(net863),
    .Y(\reg_module/_06065_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13382_  (.A(\reg_module/_06064_ ),
    .B(\reg_module/_05758_ ),
    .C(\reg_module/_06065_ ),
    .Y(\reg_module/_06066_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13383_  (.A(\reg_module/_06063_ ),
    .B(\reg_module/_06066_ ),
    .Y(\reg_module/_06067_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13384_  (.A(\reg_module/_06067_ ),
    .B(net681),
    .Y(\reg_module/_06068_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13385_  (.A(\reg_module/_05013_ ),
    .X(\reg_module/_06069_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13386_  (.A(\reg_module/_06069_ ),
    .B(\reg_module/gprf[941] ),
    .Y(\reg_module/_06070_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13387_  (.A(\reg_module/gprf[909] ),
    .B(net849),
    .Y(\reg_module/_06071_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13388_  (.A(\reg_module/_06070_ ),
    .B(net736),
    .C(\reg_module/_06071_ ),
    .Y(\reg_module/_06072_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13389_  (.A(\reg_module/_05100_ ),
    .X(\reg_module/_06073_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13390_  (.A(\reg_module/_06073_ ),
    .B(\reg_module/gprf[1005] ),
    .Y(\reg_module/_06074_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13391_  (.A(\reg_module/gprf[973] ),
    .B(net848),
    .Y(\reg_module/_06075_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13392_  (.A(\reg_module/_06074_ ),
    .B(\reg_module/_05767_ ),
    .C(\reg_module/_06075_ ),
    .Y(\reg_module/_06076_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13393_  (.A(\reg_module/_06072_ ),
    .B(\reg_module/_06076_ ),
    .Y(\reg_module/_06077_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13394_  (.A(\reg_module/_06077_ ),
    .B(\reg_module/_06000_ ),
    .Y(\reg_module/_06078_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13395_  (.A(\reg_module/_06068_ ),
    .B(\reg_module/_06078_ ),
    .C(\reg_module/_05539_ ),
    .Y(\reg_module/_06079_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13396_  (.A(\reg_module/_05694_ ),
    .B(\reg_module/gprf[685] ),
    .Y(\reg_module/_06080_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13397_  (.A(\reg_module/gprf[653] ),
    .B(net863),
    .Y(\reg_module/_06081_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13398_  (.A(\reg_module/_06080_ ),
    .B(net746),
    .C(\reg_module/_06081_ ),
    .Y(\reg_module/_06082_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13399_  (.A(\reg_module/_05078_ ),
    .X(\reg_module/_06083_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13400_  (.A(\reg_module/_06083_ ),
    .B(\reg_module/gprf[749] ),
    .Y(\reg_module/_06084_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13401_  (.A(\reg_module/gprf[717] ),
    .B(net863),
    .Y(\reg_module/_06085_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13402_  (.A(\reg_module/_06084_ ),
    .B(\reg_module/_05929_ ),
    .C(\reg_module/_06085_ ),
    .Y(\reg_module/_06086_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13403_  (.A(\reg_module/_06082_ ),
    .B(\reg_module/_06086_ ),
    .Y(\reg_module/_06087_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13404_  (.A(\reg_module/_06087_ ),
    .B(\reg_module/_05856_ ),
    .Y(\reg_module/_06088_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13405_  (.A(\reg_module/_05781_ ),
    .B(\reg_module/gprf[557] ),
    .Y(\reg_module/_06089_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13406_  (.A(\reg_module/gprf[525] ),
    .B(net874),
    .Y(\reg_module/_06090_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13407_  (.A(\reg_module/_06089_ ),
    .B(net749),
    .C(\reg_module/_06090_ ),
    .Y(\reg_module/_06091_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13408_  (.A(\reg_module/_05937_ ),
    .B(\reg_module/gprf[621] ),
    .Y(\reg_module/_06092_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13409_  (.A(\reg_module/gprf[589] ),
    .B(net868),
    .Y(\reg_module/_06093_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13410_  (.A(\reg_module/_06092_ ),
    .B(\reg_module/_06015_ ),
    .C(\reg_module/_06093_ ),
    .Y(\reg_module/_06094_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13411_  (.A(\reg_module/_06091_ ),
    .B(\reg_module/_06094_ ),
    .Y(\reg_module/_06095_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13412_  (.A(\reg_module/_06095_ ),
    .B(net684),
    .Y(\reg_module/_06096_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13413_  (.A(\reg_module/_06088_ ),
    .B(\reg_module/_06096_ ),
    .C(net651),
    .Y(\reg_module/_06097_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13414_  (.A(\reg_module/_06079_ ),
    .B(\reg_module/_06097_ ),
    .Y(\reg_module/_06098_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13415_  (.A(\reg_module/_06098_ ),
    .B(\reg_module/_05792_ ),
    .Y(\reg_module/_06099_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13416_  (.A(\reg_module/_05869_ ),
    .B(\reg_module/gprf[301] ),
    .Y(\reg_module/_06100_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13417_  (.A(\reg_module/gprf[269] ),
    .B(net872),
    .Y(\reg_module/_06101_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13418_  (.A(\reg_module/_06100_ ),
    .B(net747),
    .C(\reg_module/_06101_ ),
    .Y(\reg_module/_06102_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13419_  (.A(\reg_module/_05964_ ),
    .B(\reg_module/gprf[365] ),
    .Y(\reg_module/_06103_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13420_  (.A(\reg_module/_05072_ ),
    .X(\reg_module/_06104_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13421_  (.A(\reg_module/gprf[333] ),
    .B(net873),
    .Y(\reg_module/_06105_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13422_  (.A(\reg_module/_06103_ ),
    .B(\reg_module/_06104_ ),
    .C(\reg_module/_06105_ ),
    .Y(\reg_module/_06106_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13423_  (.A(\reg_module/_06102_ ),
    .B(\reg_module/_06106_ ),
    .Y(\reg_module/_06107_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13424_  (.A(\reg_module/_06107_ ),
    .B(net682),
    .Y(\reg_module/_06108_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13425_  (.A(\reg_module/_05954_ ),
    .B(\reg_module/gprf[429] ),
    .Y(\reg_module/_06109_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13426_  (.A(\reg_module/gprf[397] ),
    .B(net853),
    .Y(\reg_module/_06110_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13427_  (.A(\reg_module/_06109_ ),
    .B(net739),
    .C(\reg_module/_06110_ ),
    .Y(\reg_module/_06111_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13428_  (.A(\reg_module/_05083_ ),
    .X(\reg_module/_06112_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13429_  (.A(\reg_module/_06112_ ),
    .B(\reg_module/gprf[493] ),
    .Y(\reg_module/_06113_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13430_  (.A(\reg_module/gprf[461] ),
    .B(net855),
    .Y(\reg_module/_06114_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13431_  (.A(\reg_module/_06113_ ),
    .B(\reg_module/_05726_ ),
    .C(\reg_module/_06114_ ),
    .Y(\reg_module/_06115_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13432_  (.A(\reg_module/_06111_ ),
    .B(\reg_module/_06115_ ),
    .Y(\reg_module/_06116_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13433_  (.A(\reg_module/_05056_ ),
    .X(\reg_module/_06117_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13434_  (.A(\reg_module/_06116_ ),
    .B(\reg_module/_06117_ ),
    .Y(\reg_module/_06118_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13435_  (.A(\reg_module/_06108_ ),
    .B(\reg_module/_06118_ ),
    .C(\reg_module/_06039_ ),
    .Y(\reg_module/_06119_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13436_  (.A(\reg_module/_05964_ ),
    .B(\reg_module/gprf[45] ),
    .Y(\reg_module/_06120_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13437_  (.A(\reg_module/gprf[13] ),
    .B(net876),
    .Y(\reg_module/_06121_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13438_  (.A(\reg_module/_06120_ ),
    .B(net751),
    .C(\reg_module/_06121_ ),
    .Y(\reg_module/_06122_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13439_  (.A(\reg_module/_05968_ ),
    .B(\reg_module/gprf[109] ),
    .Y(\reg_module/_06123_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13440_  (.A(\reg_module/gprf[77] ),
    .B(net875),
    .Y(\reg_module/_06124_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13441_  (.A(\reg_module/_06123_ ),
    .B(\reg_module/_05891_ ),
    .C(\reg_module/_06124_ ),
    .Y(\reg_module/_06125_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13442_  (.A(\reg_module/_06122_ ),
    .B(\reg_module/_06125_ ),
    .Y(\reg_module/_06126_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13443_  (.A(\reg_module/_06126_ ),
    .B(net684),
    .Y(\reg_module/_06127_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13444_  (.A(\reg_module/_05819_ ),
    .B(\reg_module/gprf[173] ),
    .Y(\reg_module/_06128_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13445_  (.A(\reg_module/gprf[141] ),
    .B(net875),
    .Y(\reg_module/_06129_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13446_  (.A(\reg_module/_06128_ ),
    .B(net750),
    .C(\reg_module/_06129_ ),
    .Y(\reg_module/_06130_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13447_  (.A(\reg_module/_05823_ ),
    .B(\reg_module/gprf[237] ),
    .Y(\reg_module/_06131_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13448_  (.A(\reg_module/gprf[205] ),
    .B(net868),
    .Y(\reg_module/_06132_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13449_  (.A(\reg_module/_06131_ ),
    .B(\reg_module/_05900_ ),
    .C(\reg_module/_06132_ ),
    .Y(\reg_module/_06133_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13450_  (.A(\reg_module/_06130_ ),
    .B(\reg_module/_06133_ ),
    .Y(\reg_module/_06134_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13451_  (.A(\reg_module/_06134_ ),
    .B(\reg_module/_06056_ ),
    .Y(\reg_module/_06135_ ));
 sky130_fd_sc_hd__nand3_2 \reg_module/_13452_  (.A(\reg_module/_06127_ ),
    .B(\reg_module/_06135_ ),
    .C(net651),
    .Y(\reg_module/_06136_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13453_  (.A(\reg_module/_06119_ ),
    .B(\reg_module/_06136_ ),
    .Y(\reg_module/_06137_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13454_  (.A(\reg_module/_06137_ ),
    .B(net636),
    .Y(\reg_module/_06138_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13455_  (.A(\reg_module/_06099_ ),
    .B(\reg_module/_06138_ ),
    .Y(\wRs1Data[13] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13456_  (.A(\reg_module/_05752_ ),
    .B(\reg_module/gprf[558] ),
    .Y(\reg_module/_06139_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13457_  (.A(\reg_module/gprf[526] ),
    .B(net871),
    .Y(\reg_module/_06140_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13458_  (.A(\reg_module/_06139_ ),
    .B(net747),
    .C(\reg_module/_06140_ ),
    .Y(\reg_module/_06141_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13459_  (.A(\reg_module/_05756_ ),
    .B(\reg_module/gprf[622] ),
    .Y(\reg_module/_06142_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13460_  (.A(\reg_module/gprf[590] ),
    .B(net871),
    .Y(\reg_module/_06143_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13461_  (.A(\reg_module/_06142_ ),
    .B(\reg_module/_05758_ ),
    .C(\reg_module/_06143_ ),
    .Y(\reg_module/_06144_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13462_  (.A(\reg_module/_06141_ ),
    .B(\reg_module/_06144_ ),
    .Y(\reg_module/_06145_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13463_  (.A(\reg_module/_06145_ ),
    .B(net681),
    .Y(\reg_module/_06146_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13464_  (.A(\reg_module/_06069_ ),
    .B(\reg_module/gprf[686] ),
    .Y(\reg_module/_06147_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13465_  (.A(\reg_module/gprf[654] ),
    .B(net848),
    .Y(\reg_module/_06148_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13466_  (.A(\reg_module/_06147_ ),
    .B(net737),
    .C(\reg_module/_06148_ ),
    .Y(\reg_module/_06149_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13467_  (.A(\reg_module/_06073_ ),
    .B(\reg_module/gprf[750] ),
    .Y(\reg_module/_06150_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13468_  (.A(\reg_module/gprf[718] ),
    .B(net848),
    .Y(\reg_module/_06151_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13469_  (.A(\reg_module/_06150_ ),
    .B(\reg_module/_05767_ ),
    .C(\reg_module/_06151_ ),
    .Y(\reg_module/_06152_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13470_  (.A(\reg_module/_06149_ ),
    .B(\reg_module/_06152_ ),
    .Y(\reg_module/_06153_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13471_  (.A(\reg_module/_06153_ ),
    .B(\reg_module/_06000_ ),
    .Y(\reg_module/_06154_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13472_  (.A(\reg_module/_06146_ ),
    .B(\reg_module/_06154_ ),
    .C(net653),
    .Y(\reg_module/_06155_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13473_  (.A(\reg_module/_05287_ ),
    .X(\reg_module/_06156_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13474_  (.A(\reg_module/_06156_ ),
    .B(\reg_module/gprf[814] ),
    .Y(\reg_module/_06157_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13475_  (.A(\reg_module/gprf[782] ),
    .B(net859),
    .Y(\reg_module/_06158_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13476_  (.A(\reg_module/_06157_ ),
    .B(net748),
    .C(\reg_module/_06158_ ),
    .Y(\reg_module/_06159_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13477_  (.A(\reg_module/_06083_ ),
    .B(\reg_module/gprf[878] ),
    .Y(\reg_module/_06160_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13478_  (.A(\reg_module/gprf[846] ),
    .B(net857),
    .Y(\reg_module/_06161_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13479_  (.A(\reg_module/_06160_ ),
    .B(\reg_module/_05929_ ),
    .C(\reg_module/_06161_ ),
    .Y(\reg_module/_06162_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13480_  (.A(\reg_module/_06159_ ),
    .B(\reg_module/_06162_ ),
    .Y(\reg_module/_06163_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13481_  (.A(\reg_module/_06163_ ),
    .B(net687),
    .Y(\reg_module/_06164_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13482_  (.A(\reg_module/_05781_ ),
    .B(\reg_module/gprf[942] ),
    .Y(\reg_module/_06165_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13483_  (.A(\reg_module/gprf[910] ),
    .B(net857),
    .Y(\reg_module/_06166_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13484_  (.A(\reg_module/_06165_ ),
    .B(net742),
    .C(\reg_module/_06166_ ),
    .Y(\reg_module/_06167_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13485_  (.A(\reg_module/_05937_ ),
    .B(\reg_module/gprf[1006] ),
    .Y(\reg_module/_06168_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13486_  (.A(\reg_module/gprf[974] ),
    .B(net857),
    .Y(\reg_module/_06169_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13487_  (.A(\reg_module/_06168_ ),
    .B(\reg_module/_06015_ ),
    .C(\reg_module/_06169_ ),
    .Y(\reg_module/_06170_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13488_  (.A(\reg_module/_06167_ ),
    .B(\reg_module/_06170_ ),
    .Y(\reg_module/_06171_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13489_  (.A(\reg_module/_06171_ ),
    .B(\reg_module/_05477_ ),
    .Y(\reg_module/_06172_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13490_  (.A(\reg_module/_06164_ ),
    .B(\reg_module/_06172_ ),
    .C(\reg_module/_05400_ ),
    .Y(\reg_module/_06173_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13491_  (.A(\reg_module/_06155_ ),
    .B(\reg_module/_06173_ ),
    .Y(\reg_module/_06174_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13492_  (.A(\reg_module/_06174_ ),
    .B(\reg_module/_05792_ ),
    .Y(\reg_module/_06175_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13493_  (.A(\reg_module/_05869_ ),
    .B(\reg_module/gprf[302] ),
    .Y(\reg_module/_06176_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13494_  (.A(\reg_module/gprf[270] ),
    .B(net872),
    .Y(\reg_module/_06177_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13495_  (.A(\reg_module/_06176_ ),
    .B(net748),
    .C(\reg_module/_06177_ ),
    .Y(\reg_module/_06178_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13496_  (.A(\reg_module/_05964_ ),
    .B(\reg_module/gprf[366] ),
    .Y(\reg_module/_06179_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13497_  (.A(\reg_module/gprf[334] ),
    .B(net872),
    .Y(\reg_module/_06180_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13498_  (.A(\reg_module/_06179_ ),
    .B(\reg_module/_06104_ ),
    .C(\reg_module/_06180_ ),
    .Y(\reg_module/_06181_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13499_  (.A(\reg_module/_06178_ ),
    .B(\reg_module/_06181_ ),
    .Y(\reg_module/_06182_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13500_  (.A(\reg_module/_06182_ ),
    .B(net681),
    .Y(\reg_module/_06183_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13501_  (.A(\reg_module/_05954_ ),
    .B(\reg_module/gprf[430] ),
    .Y(\reg_module/_06184_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13502_  (.A(\reg_module/gprf[398] ),
    .B(net853),
    .Y(\reg_module/_06185_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13503_  (.A(\reg_module/_06184_ ),
    .B(net739),
    .C(\reg_module/_06185_ ),
    .Y(\reg_module/_06186_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13504_  (.A(\reg_module/_06112_ ),
    .B(\reg_module/gprf[494] ),
    .Y(\reg_module/_06187_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13505_  (.A(\reg_module/_05086_ ),
    .X(\reg_module/_06188_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13506_  (.A(\reg_module/gprf[462] ),
    .B(net853),
    .Y(\reg_module/_06189_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13507_  (.A(\reg_module/_06187_ ),
    .B(\reg_module/_06188_ ),
    .C(\reg_module/_06189_ ),
    .Y(\reg_module/_06190_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13508_  (.A(\reg_module/_06186_ ),
    .B(\reg_module/_06190_ ),
    .Y(\reg_module/_06191_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13509_  (.A(\reg_module/_06191_ ),
    .B(\reg_module/_06117_ ),
    .Y(\reg_module/_06192_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13510_  (.A(\reg_module/_06183_ ),
    .B(\reg_module/_06192_ ),
    .C(\reg_module/_06039_ ),
    .Y(\reg_module/_06193_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13511_  (.A(\reg_module/_05034_ ),
    .X(\reg_module/_06194_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13512_  (.A(\reg_module/_06194_ ),
    .B(\reg_module/gprf[46] ),
    .Y(\reg_module/_06195_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13513_  (.A(\reg_module/gprf[14] ),
    .B(net877),
    .Y(\reg_module/_06196_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13514_  (.A(\reg_module/_06195_ ),
    .B(net750),
    .C(\reg_module/_06196_ ),
    .Y(\reg_module/_06197_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13515_  (.A(\reg_module/_05968_ ),
    .B(\reg_module/gprf[110] ),
    .Y(\reg_module/_06198_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13516_  (.A(\reg_module/gprf[78] ),
    .B(net875),
    .Y(\reg_module/_06199_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13517_  (.A(\reg_module/_06198_ ),
    .B(\reg_module/_05891_ ),
    .C(\reg_module/_06199_ ),
    .Y(\reg_module/_06200_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13518_  (.A(\reg_module/_06197_ ),
    .B(\reg_module/_06200_ ),
    .Y(\reg_module/_06201_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13519_  (.A(\reg_module/_06201_ ),
    .B(net683),
    .Y(\reg_module/_06202_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13520_  (.A(\reg_module/_05819_ ),
    .B(\reg_module/gprf[174] ),
    .Y(\reg_module/_06203_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13521_  (.A(\reg_module/gprf[142] ),
    .B(net875),
    .Y(\reg_module/_06204_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13522_  (.A(\reg_module/_06203_ ),
    .B(net749),
    .C(\reg_module/_06204_ ),
    .Y(\reg_module/_06205_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13523_  (.A(\reg_module/_05823_ ),
    .B(\reg_module/gprf[238] ),
    .Y(\reg_module/_06206_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13524_  (.A(\reg_module/gprf[206] ),
    .B(net867),
    .Y(\reg_module/_06207_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13525_  (.A(\reg_module/_06206_ ),
    .B(\reg_module/_05900_ ),
    .C(\reg_module/_06207_ ),
    .Y(\reg_module/_06208_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13526_  (.A(\reg_module/_06205_ ),
    .B(\reg_module/_06208_ ),
    .Y(\reg_module/_06209_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13527_  (.A(\reg_module/_06209_ ),
    .B(\reg_module/_06056_ ),
    .Y(\reg_module/_06210_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13528_  (.A(\reg_module/_06202_ ),
    .B(\reg_module/_06210_ ),
    .C(net654),
    .Y(\reg_module/_06211_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13529_  (.A(\reg_module/_06193_ ),
    .B(\reg_module/_06211_ ),
    .Y(\reg_module/_06212_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13530_  (.A(\reg_module/_06212_ ),
    .B(net637),
    .Y(\reg_module/_06213_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13531_  (.A(\reg_module/_06175_ ),
    .B(\reg_module/_06213_ ),
    .Y(\wRs1Data[14] ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13532_  (.A(\reg_module/_05002_ ),
    .X(\reg_module/_06214_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13533_  (.A(\reg_module/_06214_ ),
    .B(\reg_module/gprf[815] ),
    .Y(\reg_module/_06215_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13534_  (.A(\reg_module/gprf[783] ),
    .B(net872),
    .Y(\reg_module/_06216_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13535_  (.A(\reg_module/_06215_ ),
    .B(net748),
    .C(\reg_module/_06216_ ),
    .Y(\reg_module/_06217_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13536_  (.A(\reg_module/_05287_ ),
    .X(\reg_module/_06218_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13537_  (.A(\reg_module/_06218_ ),
    .B(\reg_module/gprf[879] ),
    .Y(\reg_module/_06219_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13538_  (.A(\reg_module/_05072_ ),
    .X(\reg_module/_06220_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13539_  (.A(\reg_module/gprf[847] ),
    .B(net870),
    .Y(\reg_module/_06221_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13540_  (.A(\reg_module/_06219_ ),
    .B(\reg_module/_06220_ ),
    .C(\reg_module/_06221_ ),
    .Y(\reg_module/_06222_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13541_  (.A(\reg_module/_06217_ ),
    .B(\reg_module/_06222_ ),
    .Y(\reg_module/_06223_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13542_  (.A(\reg_module/_06223_ ),
    .B(net682),
    .Y(\reg_module/_06224_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13543_  (.A(\reg_module/_06069_ ),
    .B(\reg_module/gprf[943] ),
    .Y(\reg_module/_06225_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13544_  (.A(\reg_module/gprf[911] ),
    .B(net856),
    .Y(\reg_module/_06226_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13545_  (.A(\reg_module/_06225_ ),
    .B(net742),
    .C(\reg_module/_06226_ ),
    .Y(\reg_module/_06227_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13546_  (.A(\reg_module/_06073_ ),
    .B(\reg_module/gprf[1007] ),
    .Y(\reg_module/_06228_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13547_  (.A(\reg_module/_05022_ ),
    .X(\reg_module/_06229_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13548_  (.A(\reg_module/gprf[975] ),
    .B(net856),
    .Y(\reg_module/_06230_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13549_  (.A(\reg_module/_06228_ ),
    .B(\reg_module/_06229_ ),
    .C(\reg_module/_06230_ ),
    .Y(\reg_module/_06231_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13550_  (.A(\reg_module/_06227_ ),
    .B(\reg_module/_06231_ ),
    .Y(\reg_module/_06232_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13551_  (.A(\reg_module/_06232_ ),
    .B(\reg_module/_06000_ ),
    .Y(\reg_module/_06233_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13552_  (.A(\reg_module/_05538_ ),
    .X(\reg_module/_06234_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13553_  (.A(\reg_module/_06224_ ),
    .B(\reg_module/_06233_ ),
    .C(\reg_module/_06234_ ),
    .Y(\reg_module/_06235_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13554_  (.A(\reg_module/_06156_ ),
    .B(\reg_module/gprf[687] ),
    .Y(\reg_module/_06236_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13555_  (.A(\reg_module/gprf[655] ),
    .B(net849),
    .Y(\reg_module/_06237_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13556_  (.A(\reg_module/_06236_ ),
    .B(net737),
    .C(\reg_module/_06237_ ),
    .Y(\reg_module/_06238_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13557_  (.A(\reg_module/_06083_ ),
    .B(\reg_module/gprf[751] ),
    .Y(\reg_module/_06239_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13558_  (.A(\reg_module/gprf[719] ),
    .B(net849),
    .Y(\reg_module/_06240_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13559_  (.A(\reg_module/_06239_ ),
    .B(\reg_module/_05929_ ),
    .C(\reg_module/_06240_ ),
    .Y(\reg_module/_06241_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13560_  (.A(\reg_module/_06238_ ),
    .B(\reg_module/_06241_ ),
    .Y(\reg_module/_06242_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13561_  (.A(\reg_module/_06242_ ),
    .B(\reg_module/_05856_ ),
    .Y(\reg_module/_06243_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13562_  (.A(\reg_module/_05019_ ),
    .X(\reg_module/_06244_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13563_  (.A(\reg_module/_06244_ ),
    .B(\reg_module/gprf[559] ),
    .Y(\reg_module/_06245_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13564_  (.A(\reg_module/gprf[527] ),
    .B(net874),
    .Y(\reg_module/_06246_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13565_  (.A(\reg_module/_06245_ ),
    .B(net749),
    .C(\reg_module/_06246_ ),
    .Y(\reg_module/_06247_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13566_  (.A(\reg_module/_05937_ ),
    .B(\reg_module/gprf[623] ),
    .Y(\reg_module/_06248_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13567_  (.A(\reg_module/gprf[591] ),
    .B(net874),
    .Y(\reg_module/_06249_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13568_  (.A(\reg_module/_06248_ ),
    .B(\reg_module/_06015_ ),
    .C(\reg_module/_06249_ ),
    .Y(\reg_module/_06250_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13569_  (.A(\reg_module/_06247_ ),
    .B(\reg_module/_06250_ ),
    .Y(\reg_module/_06251_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13570_  (.A(\reg_module/_06251_ ),
    .B(net683),
    .Y(\reg_module/_06252_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13571_  (.A(\reg_module/_06243_ ),
    .B(\reg_module/_06252_ ),
    .C(net653),
    .Y(\reg_module/_06253_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13572_  (.A(\reg_module/_06235_ ),
    .B(\reg_module/_06253_ ),
    .Y(\reg_module/_06254_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13573_  (.A(\reg_module/_05204_ ),
    .X(\reg_module/_06255_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13574_  (.A(\reg_module/_06254_ ),
    .B(\reg_module/_06255_ ),
    .Y(\reg_module/_06256_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13575_  (.A(\reg_module/_05869_ ),
    .B(\reg_module/gprf[303] ),
    .Y(\reg_module/_06257_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13576_  (.A(\reg_module/gprf[271] ),
    .B(net872),
    .Y(\reg_module/_06258_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13577_  (.A(\reg_module/_06257_ ),
    .B(net748),
    .C(\reg_module/_06258_ ),
    .Y(\reg_module/_06259_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13578_  (.A(\reg_module/_06194_ ),
    .B(\reg_module/gprf[367] ),
    .Y(\reg_module/_06260_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13579_  (.A(\reg_module/gprf[335] ),
    .B(net872),
    .Y(\reg_module/_06261_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13580_  (.A(\reg_module/_06260_ ),
    .B(\reg_module/_06104_ ),
    .C(\reg_module/_06261_ ),
    .Y(\reg_module/_06262_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13581_  (.A(\reg_module/_06259_ ),
    .B(\reg_module/_06262_ ),
    .Y(\reg_module/_06263_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13582_  (.A(\reg_module/_06263_ ),
    .B(net681),
    .Y(\reg_module/_06264_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13583_  (.A(\reg_module/_05954_ ),
    .B(\reg_module/gprf[431] ),
    .Y(\reg_module/_06265_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13584_  (.A(\reg_module/gprf[399] ),
    .B(net853),
    .Y(\reg_module/_06266_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13585_  (.A(\reg_module/_06265_ ),
    .B(net740),
    .C(\reg_module/_06266_ ),
    .Y(\reg_module/_06267_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13586_  (.A(\reg_module/_06112_ ),
    .B(\reg_module/gprf[495] ),
    .Y(\reg_module/_06268_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13587_  (.A(\reg_module/gprf[463] ),
    .B(net853),
    .Y(\reg_module/_06269_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13588_  (.A(\reg_module/_06268_ ),
    .B(\reg_module/_06188_ ),
    .C(\reg_module/_06269_ ),
    .Y(\reg_module/_06270_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13589_  (.A(\reg_module/_06267_ ),
    .B(\reg_module/_06270_ ),
    .Y(\reg_module/_06271_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13590_  (.A(\reg_module/_06271_ ),
    .B(\reg_module/_06117_ ),
    .Y(\reg_module/_06272_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13591_  (.A(\reg_module/_06264_ ),
    .B(\reg_module/_06272_ ),
    .C(\reg_module/_06039_ ),
    .Y(\reg_module/_06273_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13592_  (.A(\reg_module/_06194_ ),
    .B(\reg_module/gprf[47] ),
    .Y(\reg_module/_06274_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13593_  (.A(\reg_module/gprf[15] ),
    .B(net876),
    .Y(\reg_module/_06275_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13594_  (.A(\reg_module/_06274_ ),
    .B(net750),
    .C(\reg_module/_06275_ ),
    .Y(\reg_module/_06276_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13595_  (.A(\reg_module/_05968_ ),
    .B(\reg_module/gprf[111] ),
    .Y(\reg_module/_06277_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13596_  (.A(\reg_module/gprf[79] ),
    .B(net876),
    .Y(\reg_module/_06278_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13597_  (.A(\reg_module/_06277_ ),
    .B(\reg_module/_05891_ ),
    .C(\reg_module/_06278_ ),
    .Y(\reg_module/_06279_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13598_  (.A(\reg_module/_06276_ ),
    .B(\reg_module/_06279_ ),
    .Y(\reg_module/_06280_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13599_  (.A(\reg_module/_06280_ ),
    .B(net683),
    .Y(\reg_module/_06281_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13600_  (.A(\reg_module/_05108_ ),
    .X(\reg_module/_06282_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13601_  (.A(\reg_module/_06282_ ),
    .B(\reg_module/gprf[175] ),
    .Y(\reg_module/_06283_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13602_  (.A(\reg_module/gprf[143] ),
    .B(net867),
    .Y(\reg_module/_06284_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13603_  (.A(\reg_module/_06283_ ),
    .B(net745),
    .C(\reg_module/_06284_ ),
    .Y(\reg_module/_06285_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13604_  (.A(\reg_module/_05113_ ),
    .X(\reg_module/_06286_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13605_  (.A(\reg_module/_06286_ ),
    .B(\reg_module/gprf[239] ),
    .Y(\reg_module/_06287_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13606_  (.A(\reg_module/gprf[207] ),
    .B(net868),
    .Y(\reg_module/_06288_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13607_  (.A(\reg_module/_06287_ ),
    .B(\reg_module/_05900_ ),
    .C(\reg_module/_06288_ ),
    .Y(\reg_module/_06289_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13608_  (.A(\reg_module/_06285_ ),
    .B(\reg_module/_06289_ ),
    .Y(\reg_module/_06290_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13609_  (.A(\reg_module/_06290_ ),
    .B(\reg_module/_06056_ ),
    .Y(\reg_module/_06291_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13610_  (.A(\reg_module/_06281_ ),
    .B(\reg_module/_06291_ ),
    .C(net651),
    .Y(\reg_module/_06292_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13611_  (.A(\reg_module/_06273_ ),
    .B(\reg_module/_06292_ ),
    .Y(\reg_module/_06293_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13612_  (.A(\reg_module/_06293_ ),
    .B(net637),
    .Y(\reg_module/_06294_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13613_  (.A(\reg_module/_06256_ ),
    .B(\reg_module/_06294_ ),
    .Y(\wRs1Data[15] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13614_  (.A(\reg_module/_06214_ ),
    .B(\reg_module/gprf[816] ),
    .Y(\reg_module/_06295_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13615_  (.A(\reg_module/gprf[784] ),
    .B(net858),
    .Y(\reg_module/_06296_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13616_  (.A(\reg_module/_06295_ ),
    .B(net742),
    .C(\reg_module/_06296_ ),
    .Y(\reg_module/_06297_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13617_  (.A(\reg_module/_06218_ ),
    .B(\reg_module/gprf[880] ),
    .Y(\reg_module/_06298_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13618_  (.A(\reg_module/gprf[848] ),
    .B(net870),
    .Y(\reg_module/_06299_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13619_  (.A(\reg_module/_06298_ ),
    .B(\reg_module/_06220_ ),
    .C(\reg_module/_06299_ ),
    .Y(\reg_module/_06300_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13620_  (.A(\reg_module/_06297_ ),
    .B(\reg_module/_06300_ ),
    .Y(\reg_module/_06301_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13621_  (.A(\reg_module/_06301_ ),
    .B(net678),
    .Y(\reg_module/_06302_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13622_  (.A(\reg_module/_06069_ ),
    .B(\reg_module/gprf[944] ),
    .Y(\reg_module/_06303_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13623_  (.A(\reg_module/gprf[912] ),
    .B(net856),
    .Y(\reg_module/_06304_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13624_  (.A(\reg_module/_06303_ ),
    .B(net742),
    .C(\reg_module/_06304_ ),
    .Y(\reg_module/_06305_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13625_  (.A(\reg_module/_06073_ ),
    .B(\reg_module/gprf[1008] ),
    .Y(\reg_module/_06306_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13626_  (.A(\reg_module/gprf[976] ),
    .B(net856),
    .Y(\reg_module/_06307_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13627_  (.A(\reg_module/_06306_ ),
    .B(\reg_module/_06229_ ),
    .C(\reg_module/_06307_ ),
    .Y(\reg_module/_06308_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13628_  (.A(\reg_module/_06305_ ),
    .B(\reg_module/_06308_ ),
    .Y(\reg_module/_06309_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13629_  (.A(\reg_module/_06309_ ),
    .B(\reg_module/_06000_ ),
    .Y(\reg_module/_06310_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13630_  (.A(\reg_module/_06302_ ),
    .B(\reg_module/_06310_ ),
    .C(\reg_module/_06234_ ),
    .Y(\reg_module/_06311_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13631_  (.A(\reg_module/_06156_ ),
    .B(\reg_module/gprf[688] ),
    .Y(\reg_module/_06312_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13632_  (.A(\reg_module/gprf[656] ),
    .B(net846),
    .Y(\reg_module/_06313_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13633_  (.A(\reg_module/_06312_ ),
    .B(net735),
    .C(\reg_module/_06313_ ),
    .Y(\reg_module/_06314_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13634_  (.A(\reg_module/_06083_ ),
    .B(\reg_module/gprf[752] ),
    .Y(\reg_module/_06315_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13635_  (.A(\reg_module/gprf[720] ),
    .B(net849),
    .Y(\reg_module/_06316_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13636_  (.A(\reg_module/_06315_ ),
    .B(\reg_module/_05929_ ),
    .C(\reg_module/_06316_ ),
    .Y(\reg_module/_06317_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13637_  (.A(\reg_module/_06314_ ),
    .B(\reg_module/_06317_ ),
    .Y(\reg_module/_06318_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13638_  (.A(\reg_module/_06318_ ),
    .B(\reg_module/_05856_ ),
    .Y(\reg_module/_06319_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13639_  (.A(\reg_module/_06244_ ),
    .B(\reg_module/gprf[560] ),
    .Y(\reg_module/_06320_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13640_  (.A(\reg_module/gprf[528] ),
    .B(net874),
    .Y(\reg_module/_06321_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13641_  (.A(\reg_module/_06320_ ),
    .B(net749),
    .C(\reg_module/_06321_ ),
    .Y(\reg_module/_06322_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13642_  (.A(\reg_module/_05937_ ),
    .B(\reg_module/gprf[624] ),
    .Y(\reg_module/_06323_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13643_  (.A(\reg_module/gprf[592] ),
    .B(net874),
    .Y(\reg_module/_06324_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13644_  (.A(\reg_module/_06323_ ),
    .B(\reg_module/_06015_ ),
    .C(\reg_module/_06324_ ),
    .Y(\reg_module/_06325_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13645_  (.A(\reg_module/_06322_ ),
    .B(\reg_module/_06325_ ),
    .Y(\reg_module/_06326_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13646_  (.A(\reg_module/_06326_ ),
    .B(net683),
    .Y(\reg_module/_06327_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13647_  (.A(\reg_module/_06319_ ),
    .B(\reg_module/_06327_ ),
    .C(net653),
    .Y(\reg_module/_06328_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13648_  (.A(\reg_module/_06311_ ),
    .B(\reg_module/_06328_ ),
    .Y(\reg_module/_06329_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13649_  (.A(\reg_module/_06329_ ),
    .B(\reg_module/_06255_ ),
    .Y(\reg_module/_06330_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13650_  (.A(\reg_module/_05029_ ),
    .X(\reg_module/_06331_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13651_  (.A(\reg_module/_06331_ ),
    .B(\reg_module/gprf[304] ),
    .Y(\reg_module/_06332_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13652_  (.A(\reg_module/gprf[272] ),
    .B(net858),
    .Y(\reg_module/_06333_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13653_  (.A(\reg_module/_06332_ ),
    .B(net743),
    .C(\reg_module/_06333_ ),
    .Y(\reg_module/_06334_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13654_  (.A(\reg_module/_06194_ ),
    .B(\reg_module/gprf[368] ),
    .Y(\reg_module/_06335_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13655_  (.A(\reg_module/gprf[336] ),
    .B(net858),
    .Y(\reg_module/_06336_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13656_  (.A(\reg_module/_06335_ ),
    .B(\reg_module/_06104_ ),
    .C(\reg_module/_06336_ ),
    .Y(\reg_module/_06337_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13657_  (.A(\reg_module/_06334_ ),
    .B(\reg_module/_06337_ ),
    .Y(\reg_module/_06338_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13658_  (.A(\reg_module/_06338_ ),
    .B(net678),
    .Y(\reg_module/_06339_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13659_  (.A(\reg_module/_05954_ ),
    .B(\reg_module/gprf[432] ),
    .Y(\reg_module/_06340_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13660_  (.A(\reg_module/gprf[400] ),
    .B(net854),
    .Y(\reg_module/_06341_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13661_  (.A(\reg_module/_06340_ ),
    .B(net740),
    .C(\reg_module/_06341_ ),
    .Y(\reg_module/_06342_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13662_  (.A(\reg_module/_06112_ ),
    .B(\reg_module/gprf[496] ),
    .Y(\reg_module/_06343_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13663_  (.A(\reg_module/gprf[464] ),
    .B(net855),
    .Y(\reg_module/_06344_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13664_  (.A(\reg_module/_06343_ ),
    .B(\reg_module/_06188_ ),
    .C(\reg_module/_06344_ ),
    .Y(\reg_module/_06345_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13665_  (.A(\reg_module/_06342_ ),
    .B(\reg_module/_06345_ ),
    .Y(\reg_module/_06346_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13666_  (.A(\reg_module/_06346_ ),
    .B(\reg_module/_06117_ ),
    .Y(\reg_module/_06347_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13667_  (.A(\reg_module/_06339_ ),
    .B(\reg_module/_06347_ ),
    .C(\reg_module/_06039_ ),
    .Y(\reg_module/_06348_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13668_  (.A(\reg_module/_06194_ ),
    .B(\reg_module/gprf[48] ),
    .Y(\reg_module/_06349_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13669_  (.A(\reg_module/gprf[16] ),
    .B(net877),
    .Y(\reg_module/_06350_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13670_  (.A(\reg_module/_06349_ ),
    .B(net750),
    .C(\reg_module/_06350_ ),
    .Y(\reg_module/_06351_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13671_  (.A(\reg_module/_05968_ ),
    .B(\reg_module/gprf[112] ),
    .Y(\reg_module/_06352_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13672_  (.A(\reg_module/_04997_ ),
    .X(\reg_module/_06353_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13673_  (.A(\reg_module/gprf[80] ),
    .B(net876),
    .Y(\reg_module/_06354_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13674_  (.A(\reg_module/_06352_ ),
    .B(\reg_module/_06353_ ),
    .C(\reg_module/_06354_ ),
    .Y(\reg_module/_06355_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13675_  (.A(\reg_module/_06351_ ),
    .B(\reg_module/_06355_ ),
    .Y(\reg_module/_06356_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13676_  (.A(\reg_module/_06356_ ),
    .B(net683),
    .Y(\reg_module/_06357_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13677_  (.A(\reg_module/_06282_ ),
    .B(\reg_module/gprf[176] ),
    .Y(\reg_module/_06358_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13678_  (.A(\reg_module/gprf[144] ),
    .B(net867),
    .Y(\reg_module/_06359_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13679_  (.A(\reg_module/_06358_ ),
    .B(net745),
    .C(\reg_module/_06359_ ),
    .Y(\reg_module/_06360_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13680_  (.A(\reg_module/_06286_ ),
    .B(\reg_module/gprf[240] ),
    .Y(\reg_module/_06361_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13681_  (.A(\reg_module/_05071_ ),
    .X(\reg_module/_06362_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13682_  (.A(\reg_module/gprf[208] ),
    .B(net865),
    .Y(\reg_module/_06363_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13683_  (.A(\reg_module/_06361_ ),
    .B(\reg_module/_06362_ ),
    .C(\reg_module/_06363_ ),
    .Y(\reg_module/_06364_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13684_  (.A(\reg_module/_06360_ ),
    .B(\reg_module/_06364_ ),
    .Y(\reg_module/_06365_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13685_  (.A(\reg_module/_06365_ ),
    .B(\reg_module/_06056_ ),
    .Y(\reg_module/_06366_ ));
 sky130_fd_sc_hd__nand3_2 \reg_module/_13686_  (.A(\reg_module/_06357_ ),
    .B(\reg_module/_06366_ ),
    .C(net652),
    .Y(\reg_module/_06367_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13687_  (.A(\reg_module/_06348_ ),
    .B(\reg_module/_06367_ ),
    .Y(\reg_module/_06368_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13688_  (.A(\reg_module/_06368_ ),
    .B(net636),
    .Y(\reg_module/_06369_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13689_  (.A(\reg_module/_06330_ ),
    .B(\reg_module/_06369_ ),
    .Y(\wRs1Data[16] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13690_  (.A(\reg_module/_06214_ ),
    .B(\reg_module/gprf[561] ),
    .Y(\reg_module/_06370_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13691_  (.A(\reg_module/gprf[529] ),
    .B(net870),
    .Y(\reg_module/_06371_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13692_  (.A(\reg_module/_06370_ ),
    .B(net747),
    .C(\reg_module/_06371_ ),
    .Y(\reg_module/_06372_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13693_  (.A(\reg_module/_06218_ ),
    .B(\reg_module/gprf[625] ),
    .Y(\reg_module/_06373_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13694_  (.A(\reg_module/gprf[593] ),
    .B(net870),
    .Y(\reg_module/_06374_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13695_  (.A(\reg_module/_06373_ ),
    .B(\reg_module/_06220_ ),
    .C(\reg_module/_06374_ ),
    .Y(\reg_module/_06375_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13696_  (.A(\reg_module/_06372_ ),
    .B(\reg_module/_06375_ ),
    .Y(\reg_module/_06376_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13697_  (.A(\reg_module/_06376_ ),
    .B(net682),
    .Y(\reg_module/_06377_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13698_  (.A(\reg_module/_06069_ ),
    .B(\reg_module/gprf[689] ),
    .Y(\reg_module/_06378_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13699_  (.A(\reg_module/gprf[657] ),
    .B(net846),
    .Y(\reg_module/_06379_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13700_  (.A(\reg_module/_06378_ ),
    .B(net738),
    .C(\reg_module/_06379_ ),
    .Y(\reg_module/_06380_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13701_  (.A(\reg_module/_06073_ ),
    .B(\reg_module/gprf[753] ),
    .Y(\reg_module/_06381_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13702_  (.A(\reg_module/gprf[721] ),
    .B(net848),
    .Y(\reg_module/_06382_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13703_  (.A(\reg_module/_06381_ ),
    .B(\reg_module/_06229_ ),
    .C(\reg_module/_06382_ ),
    .Y(\reg_module/_06383_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13704_  (.A(\reg_module/_06380_ ),
    .B(\reg_module/_06383_ ),
    .Y(\reg_module/_06384_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13705_  (.A(\reg_module/_06384_ ),
    .B(\reg_module/_06000_ ),
    .Y(\reg_module/_06385_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13706_  (.A(\reg_module/_06377_ ),
    .B(\reg_module/_06385_ ),
    .C(net653),
    .Y(\reg_module/_06386_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13707_  (.A(\reg_module/_06156_ ),
    .B(\reg_module/gprf[817] ),
    .Y(\reg_module/_06387_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13708_  (.A(\reg_module/gprf[785] ),
    .B(net858),
    .Y(\reg_module/_06388_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13709_  (.A(\reg_module/_06387_ ),
    .B(net743),
    .C(\reg_module/_06388_ ),
    .Y(\reg_module/_06389_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13710_  (.A(\reg_module/_06083_ ),
    .B(\reg_module/gprf[881] ),
    .Y(\reg_module/_06390_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13711_  (.A(\reg_module/_05037_ ),
    .X(\reg_module/_06391_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13712_  (.A(\reg_module/gprf[849] ),
    .B(net857),
    .Y(\reg_module/_06392_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13713_  (.A(\reg_module/_06390_ ),
    .B(\reg_module/_06391_ ),
    .C(\reg_module/_06392_ ),
    .Y(\reg_module/_06393_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13714_  (.A(\reg_module/_06389_ ),
    .B(\reg_module/_06393_ ),
    .Y(\reg_module/_06394_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13715_  (.A(\reg_module/_06394_ ),
    .B(net678),
    .Y(\reg_module/_06395_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13716_  (.A(\reg_module/_06244_ ),
    .B(\reg_module/gprf[945] ),
    .Y(\reg_module/_06396_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13717_  (.A(\reg_module/gprf[913] ),
    .B(net856),
    .Y(\reg_module/_06397_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13718_  (.A(\reg_module/_06396_ ),
    .B(net742),
    .C(\reg_module/_06397_ ),
    .Y(\reg_module/_06398_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13719_  (.A(\reg_module/_05048_ ),
    .X(\reg_module/_06399_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13720_  (.A(\reg_module/_06399_ ),
    .B(\reg_module/gprf[1009] ),
    .Y(\reg_module/_06400_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13721_  (.A(\reg_module/gprf[977] ),
    .B(net856),
    .Y(\reg_module/_06401_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13722_  (.A(\reg_module/_06400_ ),
    .B(\reg_module/_06015_ ),
    .C(\reg_module/_06401_ ),
    .Y(\reg_module/_06402_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13723_  (.A(\reg_module/_06398_ ),
    .B(\reg_module/_06402_ ),
    .Y(\reg_module/_06403_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13724_  (.A(\reg_module/_06403_ ),
    .B(\reg_module/_05477_ ),
    .Y(\reg_module/_06404_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13725_  (.A(\reg_module/_06395_ ),
    .B(\reg_module/_06404_ ),
    .C(\reg_module/_05400_ ),
    .Y(\reg_module/_06405_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13726_  (.A(\reg_module/_06386_ ),
    .B(\reg_module/_06405_ ),
    .Y(\reg_module/_06406_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13727_  (.A(\reg_module/_06406_ ),
    .B(\reg_module/_06255_ ),
    .Y(\reg_module/_06407_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13728_  (.A(\reg_module/_06331_ ),
    .B(\reg_module/gprf[305] ),
    .Y(\reg_module/_06408_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13729_  (.A(\reg_module/gprf[273] ),
    .B(net858),
    .Y(\reg_module/_06409_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13730_  (.A(\reg_module/_06408_ ),
    .B(net742),
    .C(\reg_module/_06409_ ),
    .Y(\reg_module/_06410_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13731_  (.A(\reg_module/_06194_ ),
    .B(\reg_module/gprf[369] ),
    .Y(\reg_module/_06411_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13732_  (.A(\reg_module/gprf[337] ),
    .B(net858),
    .Y(\reg_module/_06412_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13733_  (.A(\reg_module/_06411_ ),
    .B(\reg_module/_06104_ ),
    .C(\reg_module/_06412_ ),
    .Y(\reg_module/_06413_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13734_  (.A(\reg_module/_06410_ ),
    .B(\reg_module/_06413_ ),
    .Y(\reg_module/_06414_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13735_  (.A(\reg_module/_06414_ ),
    .B(net678),
    .Y(\reg_module/_06415_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13736_  (.A(\reg_module/_05043_ ),
    .X(\reg_module/_06416_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13737_  (.A(\reg_module/_06416_ ),
    .B(\reg_module/gprf[433] ),
    .Y(\reg_module/_06417_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13738_  (.A(\reg_module/gprf[401] ),
    .B(net854),
    .Y(\reg_module/_06418_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13739_  (.A(\reg_module/_06417_ ),
    .B(net739),
    .C(\reg_module/_06418_ ),
    .Y(\reg_module/_06419_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13740_  (.A(\reg_module/_06112_ ),
    .B(\reg_module/gprf[497] ),
    .Y(\reg_module/_06420_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13741_  (.A(\reg_module/gprf[465] ),
    .B(net853),
    .Y(\reg_module/_06421_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13742_  (.A(\reg_module/_06420_ ),
    .B(\reg_module/_06188_ ),
    .C(\reg_module/_06421_ ),
    .Y(\reg_module/_06422_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13743_  (.A(\reg_module/_06419_ ),
    .B(\reg_module/_06422_ ),
    .Y(\reg_module/_06423_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13744_  (.A(\reg_module/_06423_ ),
    .B(\reg_module/_06117_ ),
    .Y(\reg_module/_06424_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13745_  (.A(\reg_module/_06415_ ),
    .B(\reg_module/_06424_ ),
    .C(\reg_module/_06039_ ),
    .Y(\reg_module/_06425_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13746_  (.A(\reg_module/_05034_ ),
    .X(\reg_module/_06426_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13747_  (.A(\reg_module/_06426_ ),
    .B(\reg_module/gprf[49] ),
    .Y(\reg_module/_06427_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13748_  (.A(\reg_module/gprf[17] ),
    .B(net876),
    .Y(\reg_module/_06428_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13749_  (.A(\reg_module/_06427_ ),
    .B(net750),
    .C(\reg_module/_06428_ ),
    .Y(\reg_module/_06429_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_13750_  (.A(\reg_module/_05108_ ),
    .X(\reg_module/_06430_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13751_  (.A(\reg_module/_06430_ ),
    .B(\reg_module/gprf[113] ),
    .Y(\reg_module/_06431_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13752_  (.A(\reg_module/gprf[81] ),
    .B(net876),
    .Y(\reg_module/_06432_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13753_  (.A(\reg_module/_06431_ ),
    .B(\reg_module/_06353_ ),
    .C(\reg_module/_06432_ ),
    .Y(\reg_module/_06433_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13754_  (.A(\reg_module/_06429_ ),
    .B(\reg_module/_06433_ ),
    .Y(\reg_module/_06434_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13755_  (.A(\reg_module/_06434_ ),
    .B(net683),
    .Y(\reg_module/_06435_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13756_  (.A(\reg_module/_06282_ ),
    .B(\reg_module/gprf[177] ),
    .Y(\reg_module/_06436_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13757_  (.A(\reg_module/gprf[145] ),
    .B(net867),
    .Y(\reg_module/_06437_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13758_  (.A(\reg_module/_06436_ ),
    .B(net746),
    .C(\reg_module/_06437_ ),
    .Y(\reg_module/_06438_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13759_  (.A(\reg_module/_06286_ ),
    .B(\reg_module/gprf[241] ),
    .Y(\reg_module/_06439_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13760_  (.A(\reg_module/gprf[209] ),
    .B(net868),
    .Y(\reg_module/_06440_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13761_  (.A(\reg_module/_06439_ ),
    .B(\reg_module/_06362_ ),
    .C(\reg_module/_06440_ ),
    .Y(\reg_module/_06441_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13762_  (.A(\reg_module/_06438_ ),
    .B(\reg_module/_06441_ ),
    .Y(\reg_module/_06442_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13763_  (.A(\reg_module/_06442_ ),
    .B(\reg_module/_06056_ ),
    .Y(\reg_module/_06443_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13764_  (.A(\reg_module/_06435_ ),
    .B(\reg_module/_06443_ ),
    .C(net651),
    .Y(\reg_module/_06444_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13765_  (.A(\reg_module/_06425_ ),
    .B(\reg_module/_06444_ ),
    .Y(\reg_module/_06445_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13766_  (.A(\reg_module/_06445_ ),
    .B(net636),
    .Y(\reg_module/_06446_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13767_  (.A(\reg_module/_06407_ ),
    .B(\reg_module/_06446_ ),
    .Y(\wRs1Data[17] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13768_  (.A(\reg_module/_06214_ ),
    .B(\reg_module/gprf[818] ),
    .Y(\reg_module/_06447_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13769_  (.A(\reg_module/gprf[786] ),
    .B(net804),
    .Y(\reg_module/_06448_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13770_  (.A(\reg_module/_06447_ ),
    .B(net713),
    .C(\reg_module/_06448_ ),
    .Y(\reg_module/_06449_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13771_  (.A(\reg_module/_06218_ ),
    .B(\reg_module/gprf[882] ),
    .Y(\reg_module/_06450_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13772_  (.A(\reg_module/gprf[850] ),
    .B(net804),
    .Y(\reg_module/_06451_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13773_  (.A(\reg_module/_06450_ ),
    .B(\reg_module/_06220_ ),
    .C(\reg_module/_06451_ ),
    .Y(\reg_module/_06452_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13774_  (.A(\reg_module/_06449_ ),
    .B(\reg_module/_06452_ ),
    .Y(\reg_module/_06453_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13775_  (.A(\reg_module/_06453_ ),
    .B(net666),
    .Y(\reg_module/_06454_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13776_  (.A(\reg_module/_06069_ ),
    .B(\reg_module/gprf[946] ),
    .Y(\reg_module/_06455_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13777_  (.A(\reg_module/gprf[914] ),
    .B(net798),
    .Y(\reg_module/_06456_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13778_  (.A(\reg_module/_06455_ ),
    .B(net710),
    .C(\reg_module/_06456_ ),
    .Y(\reg_module/_06457_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13779_  (.A(\reg_module/_06073_ ),
    .B(\reg_module/gprf[1010] ),
    .Y(\reg_module/_06458_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13780_  (.A(\reg_module/gprf[978] ),
    .B(net846),
    .Y(\reg_module/_06459_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13781_  (.A(\reg_module/_06458_ ),
    .B(\reg_module/_06229_ ),
    .C(\reg_module/_06459_ ),
    .Y(\reg_module/_06460_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13782_  (.A(\reg_module/_06457_ ),
    .B(\reg_module/_06460_ ),
    .Y(\reg_module/_06461_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13783_  (.A(\reg_module/_05091_ ),
    .X(\reg_module/_06462_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13784_  (.A(\reg_module/_06461_ ),
    .B(\reg_module/_06462_ ),
    .Y(\reg_module/_06463_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13785_  (.A(\reg_module/_06454_ ),
    .B(\reg_module/_06463_ ),
    .C(\reg_module/_06234_ ),
    .Y(\reg_module/_06464_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13786_  (.A(\reg_module/_06156_ ),
    .B(\reg_module/gprf[690] ),
    .Y(\reg_module/_06465_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13787_  (.A(\reg_module/gprf[658] ),
    .B(net846),
    .Y(\reg_module/_06466_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13788_  (.A(\reg_module/_06465_ ),
    .B(net735),
    .C(\reg_module/_06466_ ),
    .Y(\reg_module/_06467_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13789_  (.A(\reg_module/_06083_ ),
    .B(\reg_module/gprf[754] ),
    .Y(\reg_module/_06468_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13790_  (.A(\reg_module/gprf[722] ),
    .B(net851),
    .Y(\reg_module/_06469_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13791_  (.A(\reg_module/_06468_ ),
    .B(\reg_module/_06391_ ),
    .C(\reg_module/_06469_ ),
    .Y(\reg_module/_06470_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13792_  (.A(\reg_module/_06467_ ),
    .B(\reg_module/_06470_ ),
    .Y(\reg_module/_06471_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13793_  (.A(\reg_module/_06471_ ),
    .B(\reg_module/_05856_ ),
    .Y(\reg_module/_06472_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13794_  (.A(\reg_module/_06244_ ),
    .B(\reg_module/gprf[562] ),
    .Y(\reg_module/_06473_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13795_  (.A(\reg_module/gprf[530] ),
    .B(net803),
    .Y(\reg_module/_06474_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13796_  (.A(\reg_module/_06473_ ),
    .B(net713),
    .C(\reg_module/_06474_ ),
    .Y(\reg_module/_06475_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13797_  (.A(\reg_module/_06399_ ),
    .B(\reg_module/gprf[626] ),
    .Y(\reg_module/_06476_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13798_  (.A(\reg_module/_05051_ ),
    .X(\reg_module/_06477_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13799_  (.A(\reg_module/gprf[594] ),
    .B(net804),
    .Y(\reg_module/_06478_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13800_  (.A(\reg_module/_06476_ ),
    .B(\reg_module/_06477_ ),
    .C(\reg_module/_06478_ ),
    .Y(\reg_module/_06479_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13801_  (.A(\reg_module/_06475_ ),
    .B(\reg_module/_06479_ ),
    .Y(\reg_module/_06480_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13802_  (.A(\reg_module/_06480_ ),
    .B(net667),
    .Y(\reg_module/_06481_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13803_  (.A(\reg_module/_06472_ ),
    .B(\reg_module/_06481_ ),
    .C(net643),
    .Y(\reg_module/_06482_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13804_  (.A(\reg_module/_06464_ ),
    .B(\reg_module/_06482_ ),
    .Y(\reg_module/_06483_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13805_  (.A(\reg_module/_06483_ ),
    .B(\reg_module/_06255_ ),
    .Y(\reg_module/_06484_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13806_  (.A(\reg_module/_06331_ ),
    .B(\reg_module/gprf[306] ),
    .Y(\reg_module/_06485_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13807_  (.A(\reg_module/gprf[274] ),
    .B(net854),
    .Y(\reg_module/_06486_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13808_  (.A(\reg_module/_06485_ ),
    .B(net740),
    .C(\reg_module/_06486_ ),
    .Y(\reg_module/_06487_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13809_  (.A(\reg_module/_06426_ ),
    .B(\reg_module/gprf[370] ),
    .Y(\reg_module/_06488_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13810_  (.A(\reg_module/gprf[338] ),
    .B(net852),
    .Y(\reg_module/_06489_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13811_  (.A(\reg_module/_06488_ ),
    .B(\reg_module/_06104_ ),
    .C(\reg_module/_06489_ ),
    .Y(\reg_module/_06490_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13812_  (.A(\reg_module/_06487_ ),
    .B(\reg_module/_06490_ ),
    .Y(\reg_module/_06491_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13813_  (.A(\reg_module/_06491_ ),
    .B(net678),
    .Y(\reg_module/_06492_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13814_  (.A(\reg_module/_06416_ ),
    .B(\reg_module/gprf[434] ),
    .Y(\reg_module/_06493_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13815_  (.A(\reg_module/gprf[402] ),
    .B(net852),
    .Y(\reg_module/_06494_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13816_  (.A(\reg_module/_06493_ ),
    .B(net739),
    .C(\reg_module/_06494_ ),
    .Y(\reg_module/_06495_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13817_  (.A(\reg_module/_06112_ ),
    .B(\reg_module/gprf[498] ),
    .Y(\reg_module/_06496_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13818_  (.A(\reg_module/gprf[466] ),
    .B(net855),
    .Y(\reg_module/_06497_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13819_  (.A(\reg_module/_06496_ ),
    .B(\reg_module/_06188_ ),
    .C(\reg_module/_06497_ ),
    .Y(\reg_module/_06498_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13820_  (.A(\reg_module/_06495_ ),
    .B(\reg_module/_06498_ ),
    .Y(\reg_module/_06499_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13821_  (.A(\reg_module/_06499_ ),
    .B(\reg_module/_06117_ ),
    .Y(\reg_module/_06500_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13822_  (.A(\reg_module/_05094_ ),
    .X(\reg_module/_06501_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13823_  (.A(\reg_module/_06492_ ),
    .B(\reg_module/_06500_ ),
    .C(\reg_module/_06501_ ),
    .Y(\reg_module/_06502_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13824_  (.A(\reg_module/_06426_ ),
    .B(\reg_module/gprf[50] ),
    .Y(\reg_module/_06503_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13825_  (.A(\reg_module/gprf[18] ),
    .B(net852),
    .Y(\reg_module/_06504_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13826_  (.A(\reg_module/_06503_ ),
    .B(net739),
    .C(\reg_module/_06504_ ),
    .Y(\reg_module/_06505_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13827_  (.A(\reg_module/_06430_ ),
    .B(\reg_module/gprf[114] ),
    .Y(\reg_module/_06506_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13828_  (.A(\reg_module/gprf[82] ),
    .B(net852),
    .Y(\reg_module/_06507_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13829_  (.A(\reg_module/_06506_ ),
    .B(\reg_module/_06353_ ),
    .C(\reg_module/_06507_ ),
    .Y(\reg_module/_06508_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13830_  (.A(\reg_module/_06505_ ),
    .B(\reg_module/_06508_ ),
    .Y(\reg_module/_06509_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13831_  (.A(\reg_module/_06509_ ),
    .B(net678),
    .Y(\reg_module/_06510_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13832_  (.A(\reg_module/_06282_ ),
    .B(\reg_module/gprf[178] ),
    .Y(\reg_module/_06511_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13833_  (.A(\reg_module/gprf[146] ),
    .B(net845),
    .Y(\reg_module/_06512_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13834_  (.A(\reg_module/_06511_ ),
    .B(net735),
    .C(\reg_module/_06512_ ),
    .Y(\reg_module/_06513_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13835_  (.A(\reg_module/_06286_ ),
    .B(\reg_module/gprf[242] ),
    .Y(\reg_module/_06514_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13836_  (.A(\reg_module/gprf[210] ),
    .B(net845),
    .Y(\reg_module/_06515_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13837_  (.A(\reg_module/_06514_ ),
    .B(\reg_module/_06362_ ),
    .C(\reg_module/_06515_ ),
    .Y(\reg_module/_06516_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13838_  (.A(\reg_module/_06513_ ),
    .B(\reg_module/_06516_ ),
    .Y(\reg_module/_06517_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13839_  (.A(\reg_module/_05009_ ),
    .X(\reg_module/_06518_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13840_  (.A(\reg_module/_06517_ ),
    .B(\reg_module/_06518_ ),
    .Y(\reg_module/_06519_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13841_  (.A(\reg_module/_06510_ ),
    .B(\reg_module/_06519_ ),
    .C(net653),
    .Y(\reg_module/_06520_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13842_  (.A(\reg_module/_06502_ ),
    .B(\reg_module/_06520_ ),
    .Y(\reg_module/_06521_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13843_  (.A(\reg_module/_06521_ ),
    .B(net636),
    .Y(\reg_module/_06522_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13844_  (.A(\reg_module/_06484_ ),
    .B(\reg_module/_06522_ ),
    .Y(\wRs1Data[18] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13845_  (.A(\reg_module/_06214_ ),
    .B(\reg_module/gprf[819] ),
    .Y(\reg_module/_06523_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13846_  (.A(\reg_module/gprf[787] ),
    .B(net805),
    .Y(\reg_module/_06524_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13847_  (.A(\reg_module/_06523_ ),
    .B(net714),
    .C(\reg_module/_06524_ ),
    .Y(\reg_module/_06525_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13848_  (.A(\reg_module/_06218_ ),
    .B(\reg_module/gprf[883] ),
    .Y(\reg_module/_06526_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13849_  (.A(\reg_module/gprf[851] ),
    .B(net806),
    .Y(\reg_module/_06527_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13850_  (.A(\reg_module/_06526_ ),
    .B(\reg_module/_06220_ ),
    .C(\reg_module/_06527_ ),
    .Y(\reg_module/_06528_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13851_  (.A(\reg_module/_06525_ ),
    .B(\reg_module/_06528_ ),
    .Y(\reg_module/_06529_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13852_  (.A(\reg_module/_06529_ ),
    .B(net666),
    .Y(\reg_module/_06530_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13853_  (.A(\reg_module/_05013_ ),
    .X(\reg_module/_06531_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13854_  (.A(\reg_module/_06531_ ),
    .B(\reg_module/gprf[947] ),
    .Y(\reg_module/_06532_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13855_  (.A(\reg_module/gprf[915] ),
    .B(net797),
    .Y(\reg_module/_06533_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13856_  (.A(\reg_module/_06532_ ),
    .B(net710),
    .C(\reg_module/_06533_ ),
    .Y(\reg_module/_06534_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13857_  (.A(\reg_module/_05100_ ),
    .X(\reg_module/_06535_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13858_  (.A(\reg_module/_06535_ ),
    .B(\reg_module/gprf[1011] ),
    .Y(\reg_module/_06536_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13859_  (.A(\reg_module/gprf[979] ),
    .B(net798),
    .Y(\reg_module/_06537_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13860_  (.A(\reg_module/_06536_ ),
    .B(\reg_module/_06229_ ),
    .C(\reg_module/_06537_ ),
    .Y(\reg_module/_06538_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13861_  (.A(\reg_module/_06534_ ),
    .B(\reg_module/_06538_ ),
    .Y(\reg_module/_06539_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13862_  (.A(\reg_module/_06539_ ),
    .B(\reg_module/_06462_ ),
    .Y(\reg_module/_06540_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13863_  (.A(\reg_module/_06530_ ),
    .B(\reg_module/_06540_ ),
    .C(\reg_module/_06234_ ),
    .Y(\reg_module/_06541_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13864_  (.A(\reg_module/_06156_ ),
    .B(\reg_module/gprf[691] ),
    .Y(\reg_module/_06542_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13865_  (.A(\reg_module/gprf[659] ),
    .B(net851),
    .Y(\reg_module/_06543_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13866_  (.A(\reg_module/_06542_ ),
    .B(net735),
    .C(\reg_module/_06543_ ),
    .Y(\reg_module/_06544_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13867_  (.A(\reg_module/_05078_ ),
    .X(\reg_module/_06545_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13868_  (.A(\reg_module/_06545_ ),
    .B(\reg_module/gprf[755] ),
    .Y(\reg_module/_06546_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13869_  (.A(\reg_module/gprf[723] ),
    .B(net798),
    .Y(\reg_module/_06547_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13870_  (.A(\reg_module/_06546_ ),
    .B(\reg_module/_06391_ ),
    .C(\reg_module/_06547_ ),
    .Y(\reg_module/_06548_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13871_  (.A(\reg_module/_06544_ ),
    .B(\reg_module/_06548_ ),
    .Y(\reg_module/_06549_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13872_  (.A(\reg_module/_05010_ ),
    .X(\reg_module/_06550_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13873_  (.A(\reg_module/_06549_ ),
    .B(\reg_module/_06550_ ),
    .Y(\reg_module/_06551_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13874_  (.A(\reg_module/_06244_ ),
    .B(\reg_module/gprf[563] ),
    .Y(\reg_module/_06552_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13875_  (.A(\reg_module/gprf[531] ),
    .B(net803),
    .Y(\reg_module/_06553_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13876_  (.A(\reg_module/_06552_ ),
    .B(net713),
    .C(\reg_module/_06553_ ),
    .Y(\reg_module/_06554_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13877_  (.A(\reg_module/_06399_ ),
    .B(\reg_module/gprf[627] ),
    .Y(\reg_module/_06555_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13878_  (.A(\reg_module/gprf[595] ),
    .B(net803),
    .Y(\reg_module/_06556_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13879_  (.A(\reg_module/_06555_ ),
    .B(\reg_module/_06477_ ),
    .C(\reg_module/_06556_ ),
    .Y(\reg_module/_06557_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13880_  (.A(\reg_module/_06554_ ),
    .B(\reg_module/_06557_ ),
    .Y(\reg_module/_06558_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13881_  (.A(\reg_module/_06558_ ),
    .B(net667),
    .Y(\reg_module/_06559_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13882_  (.A(\reg_module/_06551_ ),
    .B(\reg_module/_06559_ ),
    .C(net643),
    .Y(\reg_module/_06560_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13883_  (.A(\reg_module/_06541_ ),
    .B(\reg_module/_06560_ ),
    .Y(\reg_module/_06561_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13884_  (.A(\reg_module/_06561_ ),
    .B(\reg_module/_06255_ ),
    .Y(\reg_module/_06562_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13885_  (.A(\reg_module/_06331_ ),
    .B(\reg_module/gprf[307] ),
    .Y(\reg_module/_06563_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13886_  (.A(\reg_module/gprf[275] ),
    .B(net805),
    .Y(\reg_module/_06564_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13887_  (.A(\reg_module/_06563_ ),
    .B(net714),
    .C(\reg_module/_06564_ ),
    .Y(\reg_module/_06565_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13888_  (.A(\reg_module/_06426_ ),
    .B(\reg_module/gprf[371] ),
    .Y(\reg_module/_06566_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_13889_  (.A(\reg_module/_05037_ ),
    .X(\reg_module/_06567_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13890_  (.A(\reg_module/gprf[339] ),
    .B(net806),
    .Y(\reg_module/_06568_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13891_  (.A(\reg_module/_06566_ ),
    .B(\reg_module/_06567_ ),
    .C(\reg_module/_06568_ ),
    .Y(\reg_module/_06569_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13892_  (.A(\reg_module/_06565_ ),
    .B(\reg_module/_06569_ ),
    .Y(\reg_module/_06570_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13893_  (.A(\reg_module/_06570_ ),
    .B(net666),
    .Y(\reg_module/_06571_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13894_  (.A(\reg_module/_06416_ ),
    .B(\reg_module/gprf[435] ),
    .Y(\reg_module/_06572_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13895_  (.A(\reg_module/gprf[403] ),
    .B(net804),
    .Y(\reg_module/_06573_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13896_  (.A(\reg_module/_06572_ ),
    .B(net741),
    .C(\reg_module/_06573_ ),
    .Y(\reg_module/_06574_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13897_  (.A(\reg_module/_05083_ ),
    .X(\reg_module/_06575_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13898_  (.A(\reg_module/_06575_ ),
    .B(\reg_module/gprf[499] ),
    .Y(\reg_module/_06576_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13899_  (.A(\reg_module/gprf[467] ),
    .B(net855),
    .Y(\reg_module/_06577_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13900_  (.A(\reg_module/_06576_ ),
    .B(\reg_module/_06188_ ),
    .C(\reg_module/_06577_ ),
    .Y(\reg_module/_06578_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13901_  (.A(\reg_module/_06574_ ),
    .B(\reg_module/_06578_ ),
    .Y(\reg_module/_06579_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_13902_  (.A(\reg_module/_05056_ ),
    .X(\reg_module/_06580_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13903_  (.A(\reg_module/_06579_ ),
    .B(\reg_module/_06580_ ),
    .Y(\reg_module/_06581_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13904_  (.A(\reg_module/_06571_ ),
    .B(\reg_module/_06581_ ),
    .C(\reg_module/_06501_ ),
    .Y(\reg_module/_06582_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13905_  (.A(\reg_module/_06426_ ),
    .B(\reg_module/gprf[51] ),
    .Y(\reg_module/_06583_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13906_  (.A(\reg_module/gprf[19] ),
    .B(net852),
    .Y(\reg_module/_06584_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13907_  (.A(\reg_module/_06583_ ),
    .B(net739),
    .C(\reg_module/_06584_ ),
    .Y(\reg_module/_06585_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13908_  (.A(\reg_module/_06430_ ),
    .B(\reg_module/gprf[115] ),
    .Y(\reg_module/_06586_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13909_  (.A(\reg_module/gprf[83] ),
    .B(net852),
    .Y(\reg_module/_06587_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13910_  (.A(\reg_module/_06586_ ),
    .B(\reg_module/_06353_ ),
    .C(\reg_module/_06587_ ),
    .Y(\reg_module/_06588_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13911_  (.A(\reg_module/_06585_ ),
    .B(\reg_module/_06588_ ),
    .Y(\reg_module/_06589_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13912_  (.A(\reg_module/_06589_ ),
    .B(net667),
    .Y(\reg_module/_06590_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13913_  (.A(\reg_module/_06282_ ),
    .B(\reg_module/gprf[179] ),
    .Y(\reg_module/_06591_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13914_  (.A(\reg_module/gprf[147] ),
    .B(net795),
    .Y(\reg_module/_06592_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13915_  (.A(\reg_module/_06591_ ),
    .B(net709),
    .C(\reg_module/_06592_ ),
    .Y(\reg_module/_06593_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13916_  (.A(\reg_module/_06286_ ),
    .B(\reg_module/gprf[243] ),
    .Y(\reg_module/_06594_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13917_  (.A(\reg_module/gprf[211] ),
    .B(net845),
    .Y(\reg_module/_06595_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13918_  (.A(\reg_module/_06594_ ),
    .B(\reg_module/_06362_ ),
    .C(\reg_module/_06595_ ),
    .Y(\reg_module/_06596_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13919_  (.A(\reg_module/_06593_ ),
    .B(\reg_module/_06596_ ),
    .Y(\reg_module/_06597_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13920_  (.A(\reg_module/_06597_ ),
    .B(\reg_module/_06518_ ),
    .Y(\reg_module/_06598_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13921_  (.A(\reg_module/_06590_ ),
    .B(\reg_module/_06598_ ),
    .C(net644),
    .Y(\reg_module/_06599_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13922_  (.A(\reg_module/_06582_ ),
    .B(\reg_module/_06599_ ),
    .Y(\reg_module/_06600_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13923_  (.A(\reg_module/_06600_ ),
    .B(net636),
    .Y(\reg_module/_06601_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13924_  (.A(\reg_module/_06562_ ),
    .B(\reg_module/_06601_ ),
    .Y(\wRs1Data[19] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13925_  (.A(\reg_module/_06214_ ),
    .B(\reg_module/gprf[564] ),
    .Y(\reg_module/_06602_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13926_  (.A(\reg_module/gprf[532] ),
    .B(net804),
    .Y(\reg_module/_06603_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13927_  (.A(\reg_module/_06602_ ),
    .B(net713),
    .C(\reg_module/_06603_ ),
    .Y(\reg_module/_06604_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13928_  (.A(\reg_module/_06218_ ),
    .B(\reg_module/gprf[628] ),
    .Y(\reg_module/_06605_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13929_  (.A(\reg_module/gprf[596] ),
    .B(net803),
    .Y(\reg_module/_06606_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13930_  (.A(\reg_module/_06605_ ),
    .B(\reg_module/_06220_ ),
    .C(\reg_module/_06606_ ),
    .Y(\reg_module/_06607_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13931_  (.A(\reg_module/_06604_ ),
    .B(\reg_module/_06607_ ),
    .Y(\reg_module/_06608_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13932_  (.A(\reg_module/_06608_ ),
    .B(net666),
    .Y(\reg_module/_06609_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13933_  (.A(\reg_module/_06531_ ),
    .B(\reg_module/gprf[692] ),
    .Y(\reg_module/_06610_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13934_  (.A(\reg_module/gprf[660] ),
    .B(net798),
    .Y(\reg_module/_06611_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13935_  (.A(\reg_module/_06610_ ),
    .B(net710),
    .C(\reg_module/_06611_ ),
    .Y(\reg_module/_06612_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13936_  (.A(\reg_module/_06535_ ),
    .B(\reg_module/gprf[756] ),
    .Y(\reg_module/_06613_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13937_  (.A(\reg_module/gprf[724] ),
    .B(net798),
    .Y(\reg_module/_06614_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13938_  (.A(\reg_module/_06613_ ),
    .B(\reg_module/_06229_ ),
    .C(\reg_module/_06614_ ),
    .Y(\reg_module/_06615_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13939_  (.A(\reg_module/_06612_ ),
    .B(\reg_module/_06615_ ),
    .Y(\reg_module/_06616_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13940_  (.A(\reg_module/_06616_ ),
    .B(\reg_module/_06462_ ),
    .Y(\reg_module/_06617_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13941_  (.A(\reg_module/_06609_ ),
    .B(\reg_module/_06617_ ),
    .C(net644),
    .Y(\reg_module/_06618_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13942_  (.A(\reg_module/_05287_ ),
    .X(\reg_module/_06619_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13943_  (.A(\reg_module/_06619_ ),
    .B(\reg_module/gprf[820] ),
    .Y(\reg_module/_06620_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13944_  (.A(\reg_module/gprf[788] ),
    .B(net801),
    .Y(\reg_module/_06621_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13945_  (.A(\reg_module/_06620_ ),
    .B(net713),
    .C(\reg_module/_06621_ ),
    .Y(\reg_module/_06622_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13946_  (.A(\reg_module/_06545_ ),
    .B(\reg_module/gprf[884] ),
    .Y(\reg_module/_06623_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13947_  (.A(\reg_module/gprf[852] ),
    .B(net803),
    .Y(\reg_module/_06624_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13948_  (.A(\reg_module/_06623_ ),
    .B(\reg_module/_06391_ ),
    .C(\reg_module/_06624_ ),
    .Y(\reg_module/_06625_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13949_  (.A(\reg_module/_06622_ ),
    .B(\reg_module/_06625_ ),
    .Y(\reg_module/_06626_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13950_  (.A(\reg_module/_06626_ ),
    .B(net667),
    .Y(\reg_module/_06627_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13951_  (.A(\reg_module/_06244_ ),
    .B(\reg_module/gprf[948] ),
    .Y(\reg_module/_06628_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13952_  (.A(\reg_module/gprf[916] ),
    .B(net803),
    .Y(\reg_module/_06629_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13953_  (.A(\reg_module/_06628_ ),
    .B(net713),
    .C(\reg_module/_06629_ ),
    .Y(\reg_module/_06630_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13954_  (.A(\reg_module/_06399_ ),
    .B(\reg_module/gprf[1012] ),
    .Y(\reg_module/_06631_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13955_  (.A(\reg_module/gprf[980] ),
    .B(net800),
    .Y(\reg_module/_06632_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13956_  (.A(\reg_module/_06631_ ),
    .B(\reg_module/_06477_ ),
    .C(\reg_module/_06632_ ),
    .Y(\reg_module/_06633_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13957_  (.A(\reg_module/_06630_ ),
    .B(\reg_module/_06633_ ),
    .Y(\reg_module/_06634_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13958_  (.A(\reg_module/_06634_ ),
    .B(\reg_module/_05477_ ),
    .Y(\reg_module/_06635_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13959_  (.A(\reg_module/_06627_ ),
    .B(\reg_module/_06635_ ),
    .C(\reg_module/_05538_ ),
    .Y(\reg_module/_06636_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13960_  (.A(\reg_module/_06618_ ),
    .B(\reg_module/_06636_ ),
    .Y(\reg_module/_06637_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13961_  (.A(\reg_module/_06637_ ),
    .B(\reg_module/_06255_ ),
    .Y(\reg_module/_06638_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13962_  (.A(\reg_module/_06331_ ),
    .B(\reg_module/gprf[308] ),
    .Y(\reg_module/_06639_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13963_  (.A(\reg_module/gprf[276] ),
    .B(net802),
    .Y(\reg_module/_06640_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13964_  (.A(\reg_module/_06639_ ),
    .B(net712),
    .C(\reg_module/_06640_ ),
    .Y(\reg_module/_06641_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13965_  (.A(\reg_module/_06426_ ),
    .B(\reg_module/gprf[372] ),
    .Y(\reg_module/_06642_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13966_  (.A(\reg_module/gprf[340] ),
    .B(net802),
    .Y(\reg_module/_06643_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13967_  (.A(\reg_module/_06642_ ),
    .B(\reg_module/_06567_ ),
    .C(\reg_module/_06643_ ),
    .Y(\reg_module/_06644_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13968_  (.A(\reg_module/_06641_ ),
    .B(\reg_module/_06644_ ),
    .Y(\reg_module/_06645_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13969_  (.A(\reg_module/_06645_ ),
    .B(net668),
    .Y(\reg_module/_06646_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13970_  (.A(\reg_module/_06416_ ),
    .B(\reg_module/gprf[436] ),
    .Y(\reg_module/_06647_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13971_  (.A(\reg_module/gprf[404] ),
    .B(net788),
    .Y(\reg_module/_06648_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13972_  (.A(\reg_module/_06647_ ),
    .B(net706),
    .C(\reg_module/_06648_ ),
    .Y(\reg_module/_06649_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13973_  (.A(\reg_module/_06575_ ),
    .B(\reg_module/gprf[500] ),
    .Y(\reg_module/_06650_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_13974_  (.A(\reg_module/_05086_ ),
    .X(\reg_module/_06651_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13975_  (.A(\reg_module/gprf[468] ),
    .B(net788),
    .Y(\reg_module/_06652_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13976_  (.A(\reg_module/_06650_ ),
    .B(\reg_module/_06651_ ),
    .C(\reg_module/_06652_ ),
    .Y(\reg_module/_06653_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13977_  (.A(\reg_module/_06649_ ),
    .B(\reg_module/_06653_ ),
    .Y(\reg_module/_06654_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13978_  (.A(\reg_module/_06654_ ),
    .B(\reg_module/_06580_ ),
    .Y(\reg_module/_06655_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13979_  (.A(\reg_module/_06646_ ),
    .B(\reg_module/_06655_ ),
    .C(\reg_module/_06501_ ),
    .Y(\reg_module/_06656_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_13980_  (.A(\reg_module/_05034_ ),
    .X(\reg_module/_06657_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13981_  (.A(\reg_module/_06657_ ),
    .B(\reg_module/gprf[52] ),
    .Y(\reg_module/_06658_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13982_  (.A(\reg_module/gprf[20] ),
    .B(net805),
    .Y(\reg_module/_06659_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13983_  (.A(\reg_module/_06658_ ),
    .B(net714),
    .C(\reg_module/_06659_ ),
    .Y(\reg_module/_06660_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13984_  (.A(\reg_module/_06430_ ),
    .B(\reg_module/gprf[116] ),
    .Y(\reg_module/_06661_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13985_  (.A(\reg_module/gprf[84] ),
    .B(net805),
    .Y(\reg_module/_06662_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13986_  (.A(\reg_module/_06661_ ),
    .B(\reg_module/_06353_ ),
    .C(\reg_module/_06662_ ),
    .Y(\reg_module/_06663_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13987_  (.A(\reg_module/_06660_ ),
    .B(\reg_module/_06663_ ),
    .Y(\reg_module/_06664_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13988_  (.A(\reg_module/_06664_ ),
    .B(net666),
    .Y(\reg_module/_06665_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13989_  (.A(\reg_module/_06282_ ),
    .B(\reg_module/gprf[180] ),
    .Y(\reg_module/_06666_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13990_  (.A(\reg_module/gprf[148] ),
    .B(net795),
    .Y(\reg_module/_06667_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13991_  (.A(\reg_module/_06666_ ),
    .B(net709),
    .C(\reg_module/_06667_ ),
    .Y(\reg_module/_06668_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13992_  (.A(\reg_module/_06286_ ),
    .B(\reg_module/gprf[244] ),
    .Y(\reg_module/_06669_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13993_  (.A(\reg_module/gprf[212] ),
    .B(net796),
    .Y(\reg_module/_06670_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13994_  (.A(\reg_module/_06669_ ),
    .B(\reg_module/_06362_ ),
    .C(\reg_module/_06670_ ),
    .Y(\reg_module/_06671_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13995_  (.A(\reg_module/_06668_ ),
    .B(\reg_module/_06671_ ),
    .Y(\reg_module/_06672_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13996_  (.A(\reg_module/_06672_ ),
    .B(\reg_module/_06518_ ),
    .Y(\reg_module/_06673_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_13997_  (.A(\reg_module/_06665_ ),
    .B(\reg_module/_06673_ ),
    .C(net644),
    .Y(\reg_module/_06674_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13998_  (.A(\reg_module/_06656_ ),
    .B(\reg_module/_06674_ ),
    .Y(\reg_module/_06675_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_13999_  (.A(\reg_module/_06675_ ),
    .B(net638),
    .Y(\reg_module/_06676_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14000_  (.A(\reg_module/_06638_ ),
    .B(\reg_module/_06676_ ),
    .Y(\wRs1Data[20] ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14001_  (.A(\reg_module/_05002_ ),
    .X(\reg_module/_06677_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14002_  (.A(\reg_module/_06677_ ),
    .B(\reg_module/gprf[821] ),
    .Y(\reg_module/_06678_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14003_  (.A(\reg_module/gprf[789] ),
    .B(net801),
    .Y(\reg_module/_06679_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14004_  (.A(\reg_module/_06678_ ),
    .B(net712),
    .C(\reg_module/_06679_ ),
    .Y(\reg_module/_06680_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14005_  (.A(\reg_module/_05013_ ),
    .X(\reg_module/_06681_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14006_  (.A(\reg_module/_06681_ ),
    .B(\reg_module/gprf[885] ),
    .Y(\reg_module/_06682_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14007_  (.A(\reg_module/_05072_ ),
    .X(\reg_module/_06683_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14008_  (.A(\reg_module/gprf[853] ),
    .B(net801),
    .Y(\reg_module/_06684_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14009_  (.A(\reg_module/_06682_ ),
    .B(\reg_module/_06683_ ),
    .C(\reg_module/_06684_ ),
    .Y(\reg_module/_06685_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14010_  (.A(\reg_module/_06680_ ),
    .B(\reg_module/_06685_ ),
    .Y(\reg_module/_06686_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14011_  (.A(\reg_module/_06686_ ),
    .B(net665),
    .Y(\reg_module/_06687_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14012_  (.A(\reg_module/_06531_ ),
    .B(\reg_module/gprf[949] ),
    .Y(\reg_module/_06688_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14013_  (.A(\reg_module/gprf[917] ),
    .B(net797),
    .Y(\reg_module/_06689_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14014_  (.A(\reg_module/_06688_ ),
    .B(net710),
    .C(\reg_module/_06689_ ),
    .Y(\reg_module/_06690_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14015_  (.A(\reg_module/_06535_ ),
    .B(\reg_module/gprf[1013] ),
    .Y(\reg_module/_06691_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14016_  (.A(\reg_module/_05022_ ),
    .X(\reg_module/_06692_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14017_  (.A(\reg_module/gprf[981] ),
    .B(net793),
    .Y(\reg_module/_06693_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14018_  (.A(\reg_module/_06691_ ),
    .B(\reg_module/_06692_ ),
    .C(\reg_module/_06693_ ),
    .Y(\reg_module/_06694_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14019_  (.A(\reg_module/_06690_ ),
    .B(\reg_module/_06694_ ),
    .Y(\reg_module/_06695_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14020_  (.A(\reg_module/_06695_ ),
    .B(\reg_module/_06462_ ),
    .Y(\reg_module/_06696_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14021_  (.A(\reg_module/_06687_ ),
    .B(\reg_module/_06696_ ),
    .C(\reg_module/_06234_ ),
    .Y(\reg_module/_06697_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14022_  (.A(\reg_module/_06619_ ),
    .B(\reg_module/gprf[693] ),
    .Y(\reg_module/_06698_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14023_  (.A(\reg_module/gprf[661] ),
    .B(net797),
    .Y(\reg_module/_06699_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14024_  (.A(\reg_module/_06698_ ),
    .B(net710),
    .C(\reg_module/_06699_ ),
    .Y(\reg_module/_06700_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14025_  (.A(\reg_module/_06545_ ),
    .B(\reg_module/gprf[757] ),
    .Y(\reg_module/_06701_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14026_  (.A(\reg_module/gprf[725] ),
    .B(net797),
    .Y(\reg_module/_06702_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14027_  (.A(\reg_module/_06701_ ),
    .B(\reg_module/_06391_ ),
    .C(\reg_module/_06702_ ),
    .Y(\reg_module/_06703_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14028_  (.A(\reg_module/_06700_ ),
    .B(\reg_module/_06703_ ),
    .Y(\reg_module/_06704_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14029_  (.A(\reg_module/_06704_ ),
    .B(\reg_module/_06550_ ),
    .Y(\reg_module/_06705_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14030_  (.A(\reg_module/_05019_ ),
    .X(\reg_module/_06706_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14031_  (.A(\reg_module/_06706_ ),
    .B(\reg_module/gprf[565] ),
    .Y(\reg_module/_06707_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14032_  (.A(\reg_module/gprf[533] ),
    .B(net800),
    .Y(\reg_module/_06708_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14033_  (.A(\reg_module/_06707_ ),
    .B(net712),
    .C(\reg_module/_06708_ ),
    .Y(\reg_module/_06709_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14034_  (.A(\reg_module/_06399_ ),
    .B(\reg_module/gprf[629] ),
    .Y(\reg_module/_06710_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14035_  (.A(\reg_module/gprf[597] ),
    .B(net800),
    .Y(\reg_module/_06711_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14036_  (.A(\reg_module/_06710_ ),
    .B(\reg_module/_06477_ ),
    .C(\reg_module/_06711_ ),
    .Y(\reg_module/_06712_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14037_  (.A(\reg_module/_06709_ ),
    .B(\reg_module/_06712_ ),
    .Y(\reg_module/_06713_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14038_  (.A(\reg_module/_06713_ ),
    .B(net665),
    .Y(\reg_module/_06714_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14039_  (.A(\reg_module/_06705_ ),
    .B(\reg_module/_06714_ ),
    .C(net643),
    .Y(\reg_module/_06715_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14040_  (.A(\reg_module/_06697_ ),
    .B(\reg_module/_06715_ ),
    .Y(\reg_module/_06716_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_14041_  (.A(\reg_module/_05204_ ),
    .X(\reg_module/_06717_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14042_  (.A(\reg_module/_06716_ ),
    .B(\reg_module/_06717_ ),
    .Y(\reg_module/_06718_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14043_  (.A(\reg_module/_06331_ ),
    .B(\reg_module/gprf[309] ),
    .Y(\reg_module/_06719_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14044_  (.A(\reg_module/gprf[277] ),
    .B(net802),
    .Y(\reg_module/_06720_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14045_  (.A(\reg_module/_06719_ ),
    .B(net715),
    .C(\reg_module/_06720_ ),
    .Y(\reg_module/_06721_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14046_  (.A(\reg_module/_06657_ ),
    .B(\reg_module/gprf[373] ),
    .Y(\reg_module/_06722_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14047_  (.A(\reg_module/gprf[341] ),
    .B(net802),
    .Y(\reg_module/_06723_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14048_  (.A(\reg_module/_06722_ ),
    .B(\reg_module/_06567_ ),
    .C(\reg_module/_06723_ ),
    .Y(\reg_module/_06724_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14049_  (.A(\reg_module/_06721_ ),
    .B(\reg_module/_06724_ ),
    .Y(\reg_module/_06725_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14050_  (.A(\reg_module/_06725_ ),
    .B(net668),
    .Y(\reg_module/_06726_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14051_  (.A(\reg_module/_06416_ ),
    .B(\reg_module/gprf[437] ),
    .Y(\reg_module/_06727_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14052_  (.A(\reg_module/gprf[405] ),
    .B(net788),
    .Y(\reg_module/_06728_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14053_  (.A(\reg_module/_06727_ ),
    .B(net707),
    .C(\reg_module/_06728_ ),
    .Y(\reg_module/_06729_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14054_  (.A(\reg_module/_06575_ ),
    .B(\reg_module/gprf[501] ),
    .Y(\reg_module/_06730_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14055_  (.A(\reg_module/gprf[469] ),
    .B(net788),
    .Y(\reg_module/_06731_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14056_  (.A(\reg_module/_06730_ ),
    .B(\reg_module/_06651_ ),
    .C(\reg_module/_06731_ ),
    .Y(\reg_module/_06732_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14057_  (.A(\reg_module/_06729_ ),
    .B(\reg_module/_06732_ ),
    .Y(\reg_module/_06733_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14058_  (.A(\reg_module/_06733_ ),
    .B(\reg_module/_06580_ ),
    .Y(\reg_module/_06734_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14059_  (.A(\reg_module/_06726_ ),
    .B(\reg_module/_06734_ ),
    .C(\reg_module/_06501_ ),
    .Y(\reg_module/_06735_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14060_  (.A(\reg_module/_06657_ ),
    .B(\reg_module/gprf[53] ),
    .Y(\reg_module/_06736_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14061_  (.A(\reg_module/gprf[21] ),
    .B(net805),
    .Y(\reg_module/_06737_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14062_  (.A(\reg_module/_06736_ ),
    .B(net714),
    .C(\reg_module/_06737_ ),
    .Y(\reg_module/_06738_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14063_  (.A(\reg_module/_06430_ ),
    .B(\reg_module/gprf[117] ),
    .Y(\reg_module/_06739_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14064_  (.A(\reg_module/gprf[85] ),
    .B(net805),
    .Y(\reg_module/_06740_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14065_  (.A(\reg_module/_06739_ ),
    .B(\reg_module/_06353_ ),
    .C(\reg_module/_06740_ ),
    .Y(\reg_module/_06741_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14066_  (.A(\reg_module/_06738_ ),
    .B(\reg_module/_06741_ ),
    .Y(\reg_module/_06742_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14067_  (.A(\reg_module/_06742_ ),
    .B(net666),
    .Y(\reg_module/_06743_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14068_  (.A(\reg_module/_05083_ ),
    .X(\reg_module/_06744_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14069_  (.A(\reg_module/_06744_ ),
    .B(\reg_module/gprf[181] ),
    .Y(\reg_module/_06745_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14070_  (.A(\reg_module/gprf[149] ),
    .B(net795),
    .Y(\reg_module/_06746_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14071_  (.A(\reg_module/_06745_ ),
    .B(net709),
    .C(\reg_module/_06746_ ),
    .Y(\reg_module/_06747_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14072_  (.A(\reg_module/_05113_ ),
    .X(\reg_module/_06748_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14073_  (.A(\reg_module/_06748_ ),
    .B(\reg_module/gprf[245] ),
    .Y(\reg_module/_06749_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14074_  (.A(\reg_module/gprf[213] ),
    .B(net795),
    .Y(\reg_module/_06750_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14075_  (.A(\reg_module/_06749_ ),
    .B(\reg_module/_06362_ ),
    .C(\reg_module/_06750_ ),
    .Y(\reg_module/_06751_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14076_  (.A(\reg_module/_06747_ ),
    .B(\reg_module/_06751_ ),
    .Y(\reg_module/_06752_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14077_  (.A(\reg_module/_06752_ ),
    .B(\reg_module/_06518_ ),
    .Y(\reg_module/_06753_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14078_  (.A(\reg_module/_06743_ ),
    .B(\reg_module/_06753_ ),
    .C(net643),
    .Y(\reg_module/_06754_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14079_  (.A(\reg_module/_06735_ ),
    .B(\reg_module/_06754_ ),
    .Y(\reg_module/_06755_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14080_  (.A(\reg_module/_06755_ ),
    .B(net638),
    .Y(\reg_module/_06756_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14081_  (.A(\reg_module/_06718_ ),
    .B(\reg_module/_06756_ ),
    .Y(\wRs1Data[21] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14082_  (.A(\reg_module/_06677_ ),
    .B(\reg_module/gprf[822] ),
    .Y(\reg_module/_06757_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14083_  (.A(\reg_module/gprf[790] ),
    .B(net802),
    .Y(\reg_module/_06758_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14084_  (.A(\reg_module/_06757_ ),
    .B(net712),
    .C(\reg_module/_06758_ ),
    .Y(\reg_module/_06759_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14085_  (.A(\reg_module/_06681_ ),
    .B(\reg_module/gprf[886] ),
    .Y(\reg_module/_06760_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14086_  (.A(\reg_module/gprf[854] ),
    .B(net801),
    .Y(\reg_module/_06761_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14087_  (.A(\reg_module/_06760_ ),
    .B(\reg_module/_06683_ ),
    .C(\reg_module/_06761_ ),
    .Y(\reg_module/_06762_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14088_  (.A(\reg_module/_06759_ ),
    .B(\reg_module/_06762_ ),
    .Y(\reg_module/_06763_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14089_  (.A(\reg_module/_06763_ ),
    .B(net665),
    .Y(\reg_module/_06764_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14090_  (.A(\reg_module/_06531_ ),
    .B(\reg_module/gprf[950] ),
    .Y(\reg_module/_06765_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14091_  (.A(\reg_module/gprf[918] ),
    .B(net785),
    .Y(\reg_module/_06766_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14092_  (.A(\reg_module/_06765_ ),
    .B(net704),
    .C(\reg_module/_06766_ ),
    .Y(\reg_module/_06767_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14093_  (.A(\reg_module/_06535_ ),
    .B(\reg_module/gprf[1014] ),
    .Y(\reg_module/_06768_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14094_  (.A(\reg_module/gprf[982] ),
    .B(net785),
    .Y(\reg_module/_06769_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14095_  (.A(\reg_module/_06768_ ),
    .B(\reg_module/_06692_ ),
    .C(\reg_module/_06769_ ),
    .Y(\reg_module/_06770_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14096_  (.A(\reg_module/_06767_ ),
    .B(\reg_module/_06770_ ),
    .Y(\reg_module/_06771_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14097_  (.A(\reg_module/_06771_ ),
    .B(\reg_module/_06462_ ),
    .Y(\reg_module/_06772_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14098_  (.A(\reg_module/_06764_ ),
    .B(\reg_module/_06772_ ),
    .C(\reg_module/_06234_ ),
    .Y(\reg_module/_06773_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14099_  (.A(\reg_module/_06619_ ),
    .B(\reg_module/gprf[694] ),
    .Y(\reg_module/_06774_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14100_  (.A(\reg_module/gprf[662] ),
    .B(net797),
    .Y(\reg_module/_06775_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14101_  (.A(\reg_module/_06774_ ),
    .B(net710),
    .C(\reg_module/_06775_ ),
    .Y(\reg_module/_06776_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14102_  (.A(\reg_module/_06545_ ),
    .B(\reg_module/gprf[758] ),
    .Y(\reg_module/_06777_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14103_  (.A(\reg_module/gprf[726] ),
    .B(net797),
    .Y(\reg_module/_06778_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14104_  (.A(\reg_module/_06777_ ),
    .B(\reg_module/_06391_ ),
    .C(\reg_module/_06778_ ),
    .Y(\reg_module/_06779_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14105_  (.A(\reg_module/_06776_ ),
    .B(\reg_module/_06779_ ),
    .Y(\reg_module/_06780_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14106_  (.A(\reg_module/_06780_ ),
    .B(\reg_module/_06550_ ),
    .Y(\reg_module/_06781_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14107_  (.A(\reg_module/_06706_ ),
    .B(\reg_module/gprf[566] ),
    .Y(\reg_module/_06782_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14108_  (.A(\reg_module/gprf[534] ),
    .B(net801),
    .Y(\reg_module/_06783_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14109_  (.A(\reg_module/_06782_ ),
    .B(net712),
    .C(\reg_module/_06783_ ),
    .Y(\reg_module/_06784_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14110_  (.A(\reg_module/_06399_ ),
    .B(\reg_module/gprf[630] ),
    .Y(\reg_module/_06785_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14111_  (.A(\reg_module/gprf[598] ),
    .B(net800),
    .Y(\reg_module/_06786_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14112_  (.A(\reg_module/_06785_ ),
    .B(\reg_module/_06477_ ),
    .C(\reg_module/_06786_ ),
    .Y(\reg_module/_06787_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14113_  (.A(\reg_module/_06784_ ),
    .B(\reg_module/_06787_ ),
    .Y(\reg_module/_06788_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14114_  (.A(\reg_module/_06788_ ),
    .B(net665),
    .Y(\reg_module/_06789_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14115_  (.A(\reg_module/_06781_ ),
    .B(\reg_module/_06789_ ),
    .C(net643),
    .Y(\reg_module/_06790_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14116_  (.A(\reg_module/_06773_ ),
    .B(\reg_module/_06790_ ),
    .Y(\reg_module/_06791_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14117_  (.A(\reg_module/_06791_ ),
    .B(\reg_module/_06717_ ),
    .Y(\reg_module/_06792_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14118_  (.A(\reg_module/_05029_ ),
    .X(\reg_module/_06793_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14119_  (.A(\reg_module/_06793_ ),
    .B(\reg_module/gprf[310] ),
    .Y(\reg_module/_06794_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14120_  (.A(\reg_module/gprf[278] ),
    .B(net789),
    .Y(\reg_module/_06795_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14121_  (.A(\reg_module/_06794_ ),
    .B(net706),
    .C(\reg_module/_06795_ ),
    .Y(\reg_module/_06796_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14122_  (.A(\reg_module/_06657_ ),
    .B(\reg_module/gprf[374] ),
    .Y(\reg_module/_06797_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14123_  (.A(\reg_module/gprf[342] ),
    .B(net789),
    .Y(\reg_module/_06798_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14124_  (.A(\reg_module/_06797_ ),
    .B(\reg_module/_06567_ ),
    .C(\reg_module/_06798_ ),
    .Y(\reg_module/_06799_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14125_  (.A(\reg_module/_06796_ ),
    .B(\reg_module/_06799_ ),
    .Y(\reg_module/_06800_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14126_  (.A(\reg_module/_06800_ ),
    .B(net664),
    .Y(\reg_module/_06801_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14127_  (.A(\reg_module/_06416_ ),
    .B(\reg_module/gprf[438] ),
    .Y(\reg_module/_06802_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14128_  (.A(\reg_module/gprf[406] ),
    .B(net788),
    .Y(\reg_module/_06803_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14129_  (.A(\reg_module/_06802_ ),
    .B(net706),
    .C(\reg_module/_06803_ ),
    .Y(\reg_module/_06804_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14130_  (.A(\reg_module/_06575_ ),
    .B(\reg_module/gprf[502] ),
    .Y(\reg_module/_06805_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14131_  (.A(\reg_module/gprf[470] ),
    .B(net788),
    .Y(\reg_module/_06806_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14132_  (.A(\reg_module/_06805_ ),
    .B(\reg_module/_06651_ ),
    .C(\reg_module/_06806_ ),
    .Y(\reg_module/_06807_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14133_  (.A(\reg_module/_06804_ ),
    .B(\reg_module/_06807_ ),
    .Y(\reg_module/_06808_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14134_  (.A(\reg_module/_06808_ ),
    .B(\reg_module/_06580_ ),
    .Y(\reg_module/_06809_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14135_  (.A(\reg_module/_06801_ ),
    .B(\reg_module/_06809_ ),
    .C(\reg_module/_06501_ ),
    .Y(\reg_module/_06810_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14136_  (.A(\reg_module/_06657_ ),
    .B(\reg_module/gprf[54] ),
    .Y(\reg_module/_06811_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14137_  (.A(\reg_module/gprf[22] ),
    .B(net789),
    .Y(\reg_module/_06812_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14138_  (.A(\reg_module/_06811_ ),
    .B(net707),
    .C(\reg_module/_06812_ ),
    .Y(\reg_module/_06813_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14139_  (.A(\reg_module/_06430_ ),
    .B(\reg_module/gprf[118] ),
    .Y(\reg_module/_06814_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14140_  (.A(\reg_module/_04997_ ),
    .X(\reg_module/_06815_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14141_  (.A(\reg_module/gprf[86] ),
    .B(net789),
    .Y(\reg_module/_06816_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14142_  (.A(\reg_module/_06814_ ),
    .B(\reg_module/_06815_ ),
    .C(\reg_module/_06816_ ),
    .Y(\reg_module/_06817_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14143_  (.A(\reg_module/_06813_ ),
    .B(\reg_module/_06817_ ),
    .Y(\reg_module/_06818_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14144_  (.A(\reg_module/_06818_ ),
    .B(net664),
    .Y(\reg_module/_06819_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14145_  (.A(\reg_module/_06744_ ),
    .B(\reg_module/gprf[182] ),
    .Y(\reg_module/_06820_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14146_  (.A(\reg_module/gprf[150] ),
    .B(net795),
    .Y(\reg_module/_06821_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14147_  (.A(\reg_module/_06820_ ),
    .B(net709),
    .C(\reg_module/_06821_ ),
    .Y(\reg_module/_06822_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14148_  (.A(\reg_module/_06748_ ),
    .B(\reg_module/gprf[246] ),
    .Y(\reg_module/_06823_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14149_  (.A(\reg_module/_05071_ ),
    .X(\reg_module/_06824_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14150_  (.A(\reg_module/gprf[214] ),
    .B(net796),
    .Y(\reg_module/_06825_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14151_  (.A(\reg_module/_06823_ ),
    .B(\reg_module/_06824_ ),
    .C(\reg_module/_06825_ ),
    .Y(\reg_module/_06826_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14152_  (.A(\reg_module/_06822_ ),
    .B(\reg_module/_06826_ ),
    .Y(\reg_module/_06827_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_14153_  (.A(\reg_module/_06827_ ),
    .B(\reg_module/_06518_ ),
    .Y(\reg_module/_06828_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14154_  (.A(\reg_module/_06819_ ),
    .B(\reg_module/_06828_ ),
    .C(net646),
    .Y(\reg_module/_06829_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14155_  (.A(\reg_module/_06810_ ),
    .B(\reg_module/_06829_ ),
    .Y(\reg_module/_06830_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14156_  (.A(\reg_module/_06830_ ),
    .B(net638),
    .Y(\reg_module/_06831_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14157_  (.A(\reg_module/_06792_ ),
    .B(\reg_module/_06831_ ),
    .Y(\wRs1Data[22] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14158_  (.A(\reg_module/_06677_ ),
    .B(\reg_module/gprf[567] ),
    .Y(\reg_module/_06832_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14159_  (.A(\reg_module/gprf[535] ),
    .B(net800),
    .Y(\reg_module/_06833_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14160_  (.A(\reg_module/_06832_ ),
    .B(net712),
    .C(\reg_module/_06833_ ),
    .Y(\reg_module/_06834_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14161_  (.A(\reg_module/_06681_ ),
    .B(\reg_module/gprf[631] ),
    .Y(\reg_module/_06835_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14162_  (.A(\reg_module/gprf[599] ),
    .B(net800),
    .Y(\reg_module/_06836_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14163_  (.A(\reg_module/_06835_ ),
    .B(\reg_module/_06683_ ),
    .C(\reg_module/_06836_ ),
    .Y(\reg_module/_06837_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14164_  (.A(\reg_module/_06834_ ),
    .B(\reg_module/_06837_ ),
    .Y(\reg_module/_06838_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14165_  (.A(\reg_module/_06838_ ),
    .B(net665),
    .Y(\reg_module/_06839_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14166_  (.A(\reg_module/_06531_ ),
    .B(\reg_module/gprf[695] ),
    .Y(\reg_module/_06840_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14167_  (.A(\reg_module/gprf[663] ),
    .B(net793),
    .Y(\reg_module/_06841_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14168_  (.A(\reg_module/_06840_ ),
    .B(net711),
    .C(\reg_module/_06841_ ),
    .Y(\reg_module/_06842_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14169_  (.A(\reg_module/_06535_ ),
    .B(\reg_module/gprf[759] ),
    .Y(\reg_module/_06843_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14170_  (.A(\reg_module/gprf[727] ),
    .B(net792),
    .Y(\reg_module/_06844_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14171_  (.A(\reg_module/_06843_ ),
    .B(\reg_module/_06692_ ),
    .C(\reg_module/_06844_ ),
    .Y(\reg_module/_06845_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14172_  (.A(\reg_module/_06842_ ),
    .B(\reg_module/_06845_ ),
    .Y(\reg_module/_06846_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14173_  (.A(\reg_module/_06846_ ),
    .B(\reg_module/_06462_ ),
    .Y(\reg_module/_06847_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14174_  (.A(\reg_module/_06839_ ),
    .B(\reg_module/_06847_ ),
    .C(net643),
    .Y(\reg_module/_06848_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14175_  (.A(\reg_module/_06619_ ),
    .B(\reg_module/gprf[823] ),
    .Y(\reg_module/_06849_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14176_  (.A(\reg_module/gprf[791] ),
    .B(net793),
    .Y(\reg_module/_06850_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14177_  (.A(\reg_module/_06849_ ),
    .B(net711),
    .C(\reg_module/_06850_ ),
    .Y(\reg_module/_06851_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14178_  (.A(\reg_module/_06545_ ),
    .B(\reg_module/gprf[887] ),
    .Y(\reg_module/_06852_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14179_  (.A(\reg_module/_05022_ ),
    .X(\reg_module/_06853_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14180_  (.A(\reg_module/gprf[855] ),
    .B(net792),
    .Y(\reg_module/_06854_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14181_  (.A(\reg_module/_06852_ ),
    .B(\reg_module/_06853_ ),
    .C(\reg_module/_06854_ ),
    .Y(\reg_module/_06855_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14182_  (.A(\reg_module/_06851_ ),
    .B(\reg_module/_06855_ ),
    .Y(\reg_module/_06856_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14183_  (.A(\reg_module/_06856_ ),
    .B(net665),
    .Y(\reg_module/_06857_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14184_  (.A(\reg_module/_06706_ ),
    .B(\reg_module/gprf[951] ),
    .Y(\reg_module/_06858_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14185_  (.A(\reg_module/gprf[919] ),
    .B(net792),
    .Y(\reg_module/_06859_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14186_  (.A(\reg_module/_06858_ ),
    .B(net708),
    .C(\reg_module/_06859_ ),
    .Y(\reg_module/_06860_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14187_  (.A(\reg_module/_05048_ ),
    .X(\reg_module/_06861_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14188_  (.A(\reg_module/_06861_ ),
    .B(\reg_module/gprf[1015] ),
    .Y(\reg_module/_06862_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14189_  (.A(\reg_module/gprf[983] ),
    .B(net792),
    .Y(\reg_module/_06863_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14190_  (.A(\reg_module/_06862_ ),
    .B(\reg_module/_06477_ ),
    .C(\reg_module/_06863_ ),
    .Y(\reg_module/_06864_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14191_  (.A(\reg_module/_06860_ ),
    .B(\reg_module/_06864_ ),
    .Y(\reg_module/_06865_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14192_  (.A(\reg_module/_06865_ ),
    .B(\reg_module/_05362_ ),
    .Y(\reg_module/_06866_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14193_  (.A(\reg_module/_06857_ ),
    .B(\reg_module/_06866_ ),
    .C(\reg_module/_05538_ ),
    .Y(\reg_module/_06867_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14194_  (.A(\reg_module/_06848_ ),
    .B(\reg_module/_06867_ ),
    .Y(\reg_module/_06868_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14195_  (.A(\reg_module/_06868_ ),
    .B(\reg_module/_06717_ ),
    .Y(\reg_module/_06869_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14196_  (.A(\reg_module/_06793_ ),
    .B(\reg_module/gprf[311] ),
    .Y(\reg_module/_06870_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14197_  (.A(\reg_module/gprf[279] ),
    .B(net789),
    .Y(\reg_module/_06871_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14198_  (.A(\reg_module/_06870_ ),
    .B(net706),
    .C(\reg_module/_06871_ ),
    .Y(\reg_module/_06872_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14199_  (.A(\reg_module/_06657_ ),
    .B(\reg_module/gprf[375] ),
    .Y(\reg_module/_06873_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14200_  (.A(\reg_module/gprf[343] ),
    .B(net789),
    .Y(\reg_module/_06874_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14201_  (.A(\reg_module/_06873_ ),
    .B(\reg_module/_06567_ ),
    .C(\reg_module/_06874_ ),
    .Y(\reg_module/_06875_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14202_  (.A(\reg_module/_06872_ ),
    .B(\reg_module/_06875_ ),
    .Y(\reg_module/_06876_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14203_  (.A(\reg_module/_06876_ ),
    .B(net664),
    .Y(\reg_module/_06877_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14204_  (.A(\reg_module/_05043_ ),
    .X(\reg_module/_06878_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14205_  (.A(\reg_module/_06878_ ),
    .B(\reg_module/gprf[439] ),
    .Y(\reg_module/_06879_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14206_  (.A(\reg_module/gprf[407] ),
    .B(net790),
    .Y(\reg_module/_06880_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14207_  (.A(\reg_module/_06879_ ),
    .B(net706),
    .C(\reg_module/_06880_ ),
    .Y(\reg_module/_06881_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14208_  (.A(\reg_module/_06575_ ),
    .B(\reg_module/gprf[503] ),
    .Y(\reg_module/_06882_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14209_  (.A(\reg_module/gprf[471] ),
    .B(net790),
    .Y(\reg_module/_06883_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14210_  (.A(\reg_module/_06882_ ),
    .B(\reg_module/_06651_ ),
    .C(\reg_module/_06883_ ),
    .Y(\reg_module/_06884_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14211_  (.A(\reg_module/_06881_ ),
    .B(\reg_module/_06884_ ),
    .Y(\reg_module/_06885_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14212_  (.A(\reg_module/_06885_ ),
    .B(\reg_module/_06580_ ),
    .Y(\reg_module/_06886_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14213_  (.A(\reg_module/_06877_ ),
    .B(\reg_module/_06886_ ),
    .C(\reg_module/_06501_ ),
    .Y(\reg_module/_06887_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14214_  (.A(\reg_module/_05034_ ),
    .X(\reg_module/_06888_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14215_  (.A(\reg_module/_06888_ ),
    .B(\reg_module/gprf[55] ),
    .Y(\reg_module/_06889_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14216_  (.A(\reg_module/gprf[23] ),
    .B(net790),
    .Y(\reg_module/_06890_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14217_  (.A(\reg_module/_06889_ ),
    .B(net706),
    .C(\reg_module/_06890_ ),
    .Y(\reg_module/_06891_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_14218_  (.A(\reg_module/_05108_ ),
    .X(\reg_module/_06892_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14219_  (.A(\reg_module/_06892_ ),
    .B(\reg_module/gprf[119] ),
    .Y(\reg_module/_06893_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14220_  (.A(\reg_module/gprf[87] ),
    .B(net790),
    .Y(\reg_module/_06894_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14221_  (.A(\reg_module/_06893_ ),
    .B(\reg_module/_06815_ ),
    .C(\reg_module/_06894_ ),
    .Y(\reg_module/_06895_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14222_  (.A(\reg_module/_06891_ ),
    .B(\reg_module/_06895_ ),
    .Y(\reg_module/_06896_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14223_  (.A(\reg_module/_06896_ ),
    .B(net664),
    .Y(\reg_module/_06897_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14224_  (.A(\reg_module/_06744_ ),
    .B(\reg_module/gprf[183] ),
    .Y(\reg_module/_06898_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14225_  (.A(\reg_module/gprf[151] ),
    .B(net795),
    .Y(\reg_module/_06899_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14226_  (.A(\reg_module/_06898_ ),
    .B(net709),
    .C(\reg_module/_06899_ ),
    .Y(\reg_module/_06900_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14227_  (.A(\reg_module/_06748_ ),
    .B(\reg_module/gprf[247] ),
    .Y(\reg_module/_06901_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14228_  (.A(\reg_module/gprf[215] ),
    .B(net796),
    .Y(\reg_module/_06902_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14229_  (.A(\reg_module/_06901_ ),
    .B(\reg_module/_06824_ ),
    .C(\reg_module/_06902_ ),
    .Y(\reg_module/_06903_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14230_  (.A(\reg_module/_06900_ ),
    .B(\reg_module/_06903_ ),
    .Y(\reg_module/_06904_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_14231_  (.A(\reg_module/_06904_ ),
    .B(\reg_module/_06518_ ),
    .Y(\reg_module/_06905_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14232_  (.A(\reg_module/_06897_ ),
    .B(\reg_module/_06905_ ),
    .C(net646),
    .Y(\reg_module/_06906_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14233_  (.A(\reg_module/_06887_ ),
    .B(\reg_module/_06906_ ),
    .Y(\reg_module/_06907_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14234_  (.A(\reg_module/_06907_ ),
    .B(net638),
    .Y(\reg_module/_06908_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14235_  (.A(\reg_module/_06869_ ),
    .B(\reg_module/_06908_ ),
    .Y(\wRs1Data[23] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14236_  (.A(\reg_module/_06677_ ),
    .B(\reg_module/gprf[824] ),
    .Y(\reg_module/_06909_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14237_  (.A(\reg_module/gprf[792] ),
    .B(net794),
    .Y(\reg_module/_06910_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14238_  (.A(\reg_module/_06909_ ),
    .B(net708),
    .C(\reg_module/_06910_ ),
    .Y(\reg_module/_06911_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14239_  (.A(\reg_module/_06681_ ),
    .B(\reg_module/gprf[888] ),
    .Y(\reg_module/_06912_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14240_  (.A(\reg_module/gprf[856] ),
    .B(net794),
    .Y(\reg_module/_06913_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14241_  (.A(\reg_module/_06912_ ),
    .B(\reg_module/_06683_ ),
    .C(\reg_module/_06913_ ),
    .Y(\reg_module/_06914_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14242_  (.A(\reg_module/_06911_ ),
    .B(\reg_module/_06914_ ),
    .Y(\reg_module/_06915_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14243_  (.A(\reg_module/_06915_ ),
    .B(net669),
    .Y(\reg_module/_06916_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14244_  (.A(\reg_module/_06531_ ),
    .B(\reg_module/gprf[952] ),
    .Y(\reg_module/_06917_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14245_  (.A(\reg_module/gprf[920] ),
    .B(net786),
    .Y(\reg_module/_06918_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14246_  (.A(\reg_module/_06917_ ),
    .B(net704),
    .C(\reg_module/_06918_ ),
    .Y(\reg_module/_06919_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14247_  (.A(\reg_module/_06535_ ),
    .B(\reg_module/gprf[1016] ),
    .Y(\reg_module/_06920_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14248_  (.A(\reg_module/gprf[984] ),
    .B(net787),
    .Y(\reg_module/_06921_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14249_  (.A(\reg_module/_06920_ ),
    .B(\reg_module/_06692_ ),
    .C(\reg_module/_06921_ ),
    .Y(\reg_module/_06922_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14250_  (.A(\reg_module/_06919_ ),
    .B(\reg_module/_06922_ ),
    .Y(\reg_module/_06923_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14251_  (.A(\reg_module/_05091_ ),
    .X(\reg_module/_06924_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14252_  (.A(\reg_module/_06923_ ),
    .B(\reg_module/_06924_ ),
    .Y(\reg_module/_06925_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14253_  (.A(\reg_module/_05094_ ),
    .X(\reg_module/_06926_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14254_  (.A(\reg_module/_06916_ ),
    .B(\reg_module/_06925_ ),
    .C(\reg_module/_06926_ ),
    .Y(\reg_module/_06927_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14255_  (.A(\reg_module/_06619_ ),
    .B(\reg_module/gprf[696] ),
    .Y(\reg_module/_06928_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14256_  (.A(\reg_module/gprf[664] ),
    .B(net785),
    .Y(\reg_module/_06929_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14257_  (.A(\reg_module/_06928_ ),
    .B(net704),
    .C(\reg_module/_06929_ ),
    .Y(\reg_module/_06930_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14258_  (.A(\reg_module/_06545_ ),
    .B(\reg_module/gprf[760] ),
    .Y(\reg_module/_06931_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14259_  (.A(\reg_module/gprf[728] ),
    .B(net792),
    .Y(\reg_module/_06932_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14260_  (.A(\reg_module/_06931_ ),
    .B(\reg_module/_06853_ ),
    .C(\reg_module/_06932_ ),
    .Y(\reg_module/_06933_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14261_  (.A(\reg_module/_06930_ ),
    .B(\reg_module/_06933_ ),
    .Y(\reg_module/_06934_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14262_  (.A(\reg_module/_06934_ ),
    .B(\reg_module/_06550_ ),
    .Y(\reg_module/_06935_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14263_  (.A(\reg_module/_06706_ ),
    .B(\reg_module/gprf[568] ),
    .Y(\reg_module/_06936_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14264_  (.A(\reg_module/gprf[536] ),
    .B(net791),
    .Y(\reg_module/_06937_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14265_  (.A(\reg_module/_06936_ ),
    .B(net708),
    .C(\reg_module/_06937_ ),
    .Y(\reg_module/_06938_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14266_  (.A(\reg_module/_06861_ ),
    .B(\reg_module/gprf[632] ),
    .Y(\reg_module/_06939_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14267_  (.A(\reg_module/_05051_ ),
    .X(\reg_module/_06940_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14268_  (.A(\reg_module/gprf[600] ),
    .B(net791),
    .Y(\reg_module/_06941_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14269_  (.A(\reg_module/_06939_ ),
    .B(\reg_module/_06940_ ),
    .C(\reg_module/_06941_ ),
    .Y(\reg_module/_06942_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14270_  (.A(\reg_module/_06938_ ),
    .B(\reg_module/_06942_ ),
    .Y(\reg_module/_06943_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14271_  (.A(\reg_module/_06943_ ),
    .B(net669),
    .Y(\reg_module/_06944_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14272_  (.A(\reg_module/_06935_ ),
    .B(\reg_module/_06944_ ),
    .C(net645),
    .Y(\reg_module/_06945_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14273_  (.A(\reg_module/_06927_ ),
    .B(\reg_module/_06945_ ),
    .Y(\reg_module/_06946_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14274_  (.A(\reg_module/_06946_ ),
    .B(\reg_module/_06717_ ),
    .Y(\reg_module/_06947_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14275_  (.A(\reg_module/_06793_ ),
    .B(\reg_module/gprf[312] ),
    .Y(\reg_module/_06948_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14276_  (.A(\reg_module/gprf[280] ),
    .B(net785),
    .Y(\reg_module/_06949_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14277_  (.A(\reg_module/_06948_ ),
    .B(net705),
    .C(\reg_module/_06949_ ),
    .Y(\reg_module/_06950_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14278_  (.A(\reg_module/_06888_ ),
    .B(\reg_module/gprf[376] ),
    .Y(\reg_module/_06951_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14279_  (.A(\reg_module/gprf[344] ),
    .B(net785),
    .Y(\reg_module/_06952_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14280_  (.A(\reg_module/_06951_ ),
    .B(\reg_module/_06567_ ),
    .C(\reg_module/_06952_ ),
    .Y(\reg_module/_06953_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14281_  (.A(\reg_module/_06950_ ),
    .B(\reg_module/_06953_ ),
    .Y(\reg_module/_06954_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14282_  (.A(\reg_module/_06954_ ),
    .B(net663),
    .Y(\reg_module/_06955_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14283_  (.A(\reg_module/_06878_ ),
    .B(\reg_module/gprf[440] ),
    .Y(\reg_module/_06956_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14284_  (.A(\reg_module/gprf[408] ),
    .B(net787),
    .Y(\reg_module/_06957_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14285_  (.A(\reg_module/_06956_ ),
    .B(net703),
    .C(\reg_module/_06957_ ),
    .Y(\reg_module/_06958_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14286_  (.A(\reg_module/_06575_ ),
    .B(\reg_module/gprf[504] ),
    .Y(\reg_module/_06959_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14287_  (.A(\reg_module/gprf[472] ),
    .B(net784),
    .Y(\reg_module/_06960_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14288_  (.A(\reg_module/_06959_ ),
    .B(\reg_module/_06651_ ),
    .C(\reg_module/_06960_ ),
    .Y(\reg_module/_06961_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14289_  (.A(\reg_module/_06958_ ),
    .B(\reg_module/_06961_ ),
    .Y(\reg_module/_06962_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14290_  (.A(\reg_module/_06962_ ),
    .B(\reg_module/_06580_ ),
    .Y(\reg_module/_06963_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14291_  (.A(\reg_module/_05094_ ),
    .X(\reg_module/_06964_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14292_  (.A(\reg_module/_06955_ ),
    .B(\reg_module/_06963_ ),
    .C(\reg_module/_06964_ ),
    .Y(\reg_module/_06965_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14293_  (.A(\reg_module/_06888_ ),
    .B(\reg_module/gprf[56] ),
    .Y(\reg_module/_06966_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14294_  (.A(\reg_module/gprf[24] ),
    .B(net784),
    .Y(\reg_module/_06967_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14295_  (.A(\reg_module/_06966_ ),
    .B(net703),
    .C(\reg_module/_06967_ ),
    .Y(\reg_module/_06968_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14296_  (.A(\reg_module/_06892_ ),
    .B(\reg_module/gprf[120] ),
    .Y(\reg_module/_06969_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14297_  (.A(\reg_module/gprf[88] ),
    .B(net784),
    .Y(\reg_module/_06970_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14298_  (.A(\reg_module/_06969_ ),
    .B(\reg_module/_06815_ ),
    .C(\reg_module/_06970_ ),
    .Y(\reg_module/_06971_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14299_  (.A(\reg_module/_06968_ ),
    .B(\reg_module/_06971_ ),
    .Y(\reg_module/_06972_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14300_  (.A(\reg_module/_06972_ ),
    .B(net663),
    .Y(\reg_module/_06973_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14301_  (.A(\reg_module/_06744_ ),
    .B(\reg_module/gprf[184] ),
    .Y(\reg_module/_06974_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14302_  (.A(\reg_module/gprf[152] ),
    .B(net782),
    .Y(\reg_module/_06975_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14303_  (.A(\reg_module/_06974_ ),
    .B(net702),
    .C(\reg_module/_06975_ ),
    .Y(\reg_module/_06976_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14304_  (.A(\reg_module/_06748_ ),
    .B(\reg_module/gprf[248] ),
    .Y(\reg_module/_06977_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14305_  (.A(\reg_module/gprf[216] ),
    .B(net782),
    .Y(\reg_module/_06978_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14306_  (.A(\reg_module/_06977_ ),
    .B(\reg_module/_06824_ ),
    .C(\reg_module/_06978_ ),
    .Y(\reg_module/_06979_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14307_  (.A(\reg_module/_06976_ ),
    .B(\reg_module/_06979_ ),
    .Y(\reg_module/_06980_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14308_  (.A(\reg_module/_05009_ ),
    .X(\reg_module/_06981_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14309_  (.A(\reg_module/_06980_ ),
    .B(\reg_module/_06981_ ),
    .Y(\reg_module/_06982_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14310_  (.A(\reg_module/_06973_ ),
    .B(\reg_module/_06982_ ),
    .C(net646),
    .Y(\reg_module/_06983_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14311_  (.A(\reg_module/_06965_ ),
    .B(\reg_module/_06983_ ),
    .Y(\reg_module/_06984_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14312_  (.A(\reg_module/_06984_ ),
    .B(net638),
    .Y(\reg_module/_06985_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14313_  (.A(\reg_module/_06947_ ),
    .B(\reg_module/_06985_ ),
    .Y(\wRs1Data[24] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14314_  (.A(\reg_module/_06677_ ),
    .B(\reg_module/gprf[825] ),
    .Y(\reg_module/_06986_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14315_  (.A(\reg_module/gprf[793] ),
    .B(net796),
    .Y(\reg_module/_06987_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14316_  (.A(\reg_module/_06986_ ),
    .B(net709),
    .C(\reg_module/_06987_ ),
    .Y(\reg_module/_06988_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14317_  (.A(\reg_module/_06681_ ),
    .B(\reg_module/gprf[889] ),
    .Y(\reg_module/_06989_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14318_  (.A(\reg_module/gprf[857] ),
    .B(net796),
    .Y(\reg_module/_06990_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14319_  (.A(\reg_module/_06989_ ),
    .B(\reg_module/_06683_ ),
    .C(\reg_module/_06990_ ),
    .Y(\reg_module/_06991_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14320_  (.A(\reg_module/_06988_ ),
    .B(\reg_module/_06991_ ),
    .Y(\reg_module/_06992_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14321_  (.A(\reg_module/_06992_ ),
    .B(net669),
    .Y(\reg_module/_06993_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14322_  (.A(\reg_module/_05068_ ),
    .X(\reg_module/_06994_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14323_  (.A(\reg_module/_06994_ ),
    .B(\reg_module/gprf[953] ),
    .Y(\reg_module/_06995_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14324_  (.A(\reg_module/gprf[921] ),
    .B(net786),
    .Y(\reg_module/_06996_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14325_  (.A(\reg_module/_06995_ ),
    .B(net704),
    .C(\reg_module/_06996_ ),
    .Y(\reg_module/_06997_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14326_  (.A(\reg_module/_05100_ ),
    .X(\reg_module/_06998_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14327_  (.A(\reg_module/_06998_ ),
    .B(\reg_module/gprf[1017] ),
    .Y(\reg_module/_06999_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14328_  (.A(\reg_module/gprf[985] ),
    .B(net786),
    .Y(\reg_module/_07000_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14329_  (.A(\reg_module/_06999_ ),
    .B(\reg_module/_06692_ ),
    .C(\reg_module/_07000_ ),
    .Y(\reg_module/_07001_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14330_  (.A(\reg_module/_06997_ ),
    .B(\reg_module/_07001_ ),
    .Y(\reg_module/_07002_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14331_  (.A(\reg_module/_07002_ ),
    .B(\reg_module/_06924_ ),
    .Y(\reg_module/_07003_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14332_  (.A(\reg_module/_06993_ ),
    .B(\reg_module/_07003_ ),
    .C(\reg_module/_06926_ ),
    .Y(\reg_module/_07004_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14333_  (.A(\reg_module/_06619_ ),
    .B(\reg_module/gprf[697] ),
    .Y(\reg_module/_07005_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14334_  (.A(\reg_module/gprf[665] ),
    .B(net785),
    .Y(\reg_module/_07006_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14335_  (.A(\reg_module/_07005_ ),
    .B(net704),
    .C(\reg_module/_07006_ ),
    .Y(\reg_module/_07007_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14336_  (.A(\reg_module/_05078_ ),
    .X(\reg_module/_07008_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14337_  (.A(\reg_module/_07008_ ),
    .B(\reg_module/gprf[761] ),
    .Y(\reg_module/_07009_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14338_  (.A(\reg_module/gprf[729] ),
    .B(net792),
    .Y(\reg_module/_07010_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14339_  (.A(\reg_module/_07009_ ),
    .B(\reg_module/_06853_ ),
    .C(\reg_module/_07010_ ),
    .Y(\reg_module/_07011_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14340_  (.A(\reg_module/_07007_ ),
    .B(\reg_module/_07011_ ),
    .Y(\reg_module/_07012_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14341_  (.A(\reg_module/_07012_ ),
    .B(\reg_module/_06550_ ),
    .Y(\reg_module/_07013_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14342_  (.A(\reg_module/_06706_ ),
    .B(\reg_module/gprf[569] ),
    .Y(\reg_module/_07014_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14343_  (.A(\reg_module/gprf[537] ),
    .B(net791),
    .Y(\reg_module/_07015_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14344_  (.A(\reg_module/_07014_ ),
    .B(net708),
    .C(\reg_module/_07015_ ),
    .Y(\reg_module/_07016_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14345_  (.A(\reg_module/_06861_ ),
    .B(\reg_module/gprf[633] ),
    .Y(\reg_module/_07017_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14346_  (.A(\reg_module/gprf[601] ),
    .B(net791),
    .Y(\reg_module/_07018_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14347_  (.A(\reg_module/_07017_ ),
    .B(\reg_module/_06940_ ),
    .C(\reg_module/_07018_ ),
    .Y(\reg_module/_07019_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14348_  (.A(\reg_module/_07016_ ),
    .B(\reg_module/_07019_ ),
    .Y(\reg_module/_07020_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14349_  (.A(\reg_module/_07020_ ),
    .B(net669),
    .Y(\reg_module/_07021_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14350_  (.A(\reg_module/_07013_ ),
    .B(\reg_module/_07021_ ),
    .C(net645),
    .Y(\reg_module/_07022_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14351_  (.A(\reg_module/_07004_ ),
    .B(\reg_module/_07022_ ),
    .Y(\reg_module/_07023_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14352_  (.A(\reg_module/_07023_ ),
    .B(\reg_module/_06717_ ),
    .Y(\reg_module/_07024_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14353_  (.A(\reg_module/_06793_ ),
    .B(\reg_module/gprf[313] ),
    .Y(\reg_module/_07025_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14354_  (.A(\reg_module/gprf[281] ),
    .B(net786),
    .Y(\reg_module/_07026_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14355_  (.A(\reg_module/_07025_ ),
    .B(net702),
    .C(\reg_module/_07026_ ),
    .Y(\reg_module/_07027_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14356_  (.A(\reg_module/_06888_ ),
    .B(\reg_module/gprf[377] ),
    .Y(\reg_module/_07028_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14357_  (.A(\reg_module/_05037_ ),
    .X(\reg_module/_07029_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14358_  (.A(\reg_module/gprf[345] ),
    .B(net783),
    .Y(\reg_module/_07030_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14359_  (.A(\reg_module/_07028_ ),
    .B(\reg_module/_07029_ ),
    .C(\reg_module/_07030_ ),
    .Y(\reg_module/_07031_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14360_  (.A(\reg_module/_07027_ ),
    .B(\reg_module/_07031_ ),
    .Y(\reg_module/_07032_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14361_  (.A(\reg_module/_07032_ ),
    .B(net663),
    .Y(\reg_module/_07033_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14362_  (.A(\reg_module/_06878_ ),
    .B(\reg_module/gprf[441] ),
    .Y(\reg_module/_07034_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14363_  (.A(\reg_module/gprf[409] ),
    .B(net783),
    .Y(\reg_module/_07035_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14364_  (.A(\reg_module/_07034_ ),
    .B(net703),
    .C(\reg_module/_07035_ ),
    .Y(\reg_module/_07036_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14365_  (.A(\reg_module/_05048_ ),
    .X(\reg_module/_07037_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14366_  (.A(\reg_module/_07037_ ),
    .B(\reg_module/gprf[505] ),
    .Y(\reg_module/_07038_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14367_  (.A(\reg_module/gprf[473] ),
    .B(net784),
    .Y(\reg_module/_07039_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14368_  (.A(\reg_module/_07038_ ),
    .B(\reg_module/_06651_ ),
    .C(\reg_module/_07039_ ),
    .Y(\reg_module/_07040_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14369_  (.A(\reg_module/_07036_ ),
    .B(\reg_module/_07040_ ),
    .Y(\reg_module/_07041_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14370_  (.A(\reg_module/_05056_ ),
    .X(\reg_module/_07042_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14371_  (.A(\reg_module/_07041_ ),
    .B(\reg_module/_07042_ ),
    .Y(\reg_module/_07043_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14372_  (.A(\reg_module/_07033_ ),
    .B(\reg_module/_07043_ ),
    .C(\reg_module/_06964_ ),
    .Y(\reg_module/_07044_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14373_  (.A(\reg_module/_06888_ ),
    .B(\reg_module/gprf[57] ),
    .Y(\reg_module/_07045_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14374_  (.A(\reg_module/gprf[25] ),
    .B(net782),
    .Y(\reg_module/_07046_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14375_  (.A(\reg_module/_07045_ ),
    .B(net702),
    .C(\reg_module/_07046_ ),
    .Y(\reg_module/_07047_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14376_  (.A(\reg_module/_06892_ ),
    .B(\reg_module/gprf[121] ),
    .Y(\reg_module/_07048_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14377_  (.A(\reg_module/gprf[89] ),
    .B(net783),
    .Y(\reg_module/_07049_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14378_  (.A(\reg_module/_07048_ ),
    .B(\reg_module/_06815_ ),
    .C(\reg_module/_07049_ ),
    .Y(\reg_module/_07050_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14379_  (.A(\reg_module/_07047_ ),
    .B(\reg_module/_07050_ ),
    .Y(\reg_module/_07051_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14380_  (.A(\reg_module/_07051_ ),
    .B(net663),
    .Y(\reg_module/_07052_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14381_  (.A(\reg_module/_06744_ ),
    .B(\reg_module/gprf[185] ),
    .Y(\reg_module/_07053_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14382_  (.A(\reg_module/gprf[153] ),
    .B(net782),
    .Y(\reg_module/_07054_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14383_  (.A(\reg_module/_07053_ ),
    .B(net702),
    .C(\reg_module/_07054_ ),
    .Y(\reg_module/_07055_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14384_  (.A(\reg_module/_06748_ ),
    .B(\reg_module/gprf[249] ),
    .Y(\reg_module/_07056_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14385_  (.A(\reg_module/gprf[217] ),
    .B(net782),
    .Y(\reg_module/_07057_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14386_  (.A(\reg_module/_07056_ ),
    .B(\reg_module/_06824_ ),
    .C(\reg_module/_07057_ ),
    .Y(\reg_module/_07058_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14387_  (.A(\reg_module/_07055_ ),
    .B(\reg_module/_07058_ ),
    .Y(\reg_module/_07059_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14388_  (.A(\reg_module/_07059_ ),
    .B(\reg_module/_06981_ ),
    .Y(\reg_module/_07060_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14389_  (.A(\reg_module/_07052_ ),
    .B(\reg_module/_07060_ ),
    .C(net646),
    .Y(\reg_module/_07061_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14390_  (.A(\reg_module/_07044_ ),
    .B(\reg_module/_07061_ ),
    .Y(\reg_module/_07062_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14391_  (.A(\reg_module/_07062_ ),
    .B(net638),
    .Y(\reg_module/_07063_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14392_  (.A(\reg_module/_07024_ ),
    .B(\reg_module/_07063_ ),
    .Y(\wRs1Data[25] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14393_  (.A(\reg_module/_06677_ ),
    .B(\reg_module/gprf[570] ),
    .Y(\reg_module/_07064_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14394_  (.A(\reg_module/gprf[538] ),
    .B(net777),
    .Y(\reg_module/_07065_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14395_  (.A(\reg_module/_07064_ ),
    .B(net708),
    .C(\reg_module/_07065_ ),
    .Y(\reg_module/_07066_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14396_  (.A(\reg_module/_06681_ ),
    .B(\reg_module/gprf[634] ),
    .Y(\reg_module/_07067_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14397_  (.A(\reg_module/gprf[602] ),
    .B(net777),
    .Y(\reg_module/_07068_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14398_  (.A(\reg_module/_07067_ ),
    .B(\reg_module/_06683_ ),
    .C(\reg_module/_07068_ ),
    .Y(\reg_module/_07069_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14399_  (.A(\reg_module/_07066_ ),
    .B(\reg_module/_07069_ ),
    .Y(\reg_module/_07070_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14400_  (.A(\reg_module/_07070_ ),
    .B(net669),
    .Y(\reg_module/_07071_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14401_  (.A(\reg_module/_06994_ ),
    .B(\reg_module/gprf[698] ),
    .Y(\reg_module/_07072_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14402_  (.A(\reg_module/gprf[666] ),
    .B(net786),
    .Y(\reg_module/_07073_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14403_  (.A(\reg_module/_07072_ ),
    .B(net704),
    .C(\reg_module/_07073_ ),
    .Y(\reg_module/_07074_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14404_  (.A(\reg_module/_06998_ ),
    .B(\reg_module/gprf[762] ),
    .Y(\reg_module/_07075_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14405_  (.A(\reg_module/gprf[730] ),
    .B(net786),
    .Y(\reg_module/_07076_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14406_  (.A(\reg_module/_07075_ ),
    .B(\reg_module/_06692_ ),
    .C(\reg_module/_07076_ ),
    .Y(\reg_module/_07077_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14407_  (.A(\reg_module/_07074_ ),
    .B(\reg_module/_07077_ ),
    .Y(\reg_module/_07078_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14408_  (.A(\reg_module/_07078_ ),
    .B(\reg_module/_06924_ ),
    .Y(\reg_module/_07079_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14409_  (.A(\reg_module/_07071_ ),
    .B(\reg_module/_07079_ ),
    .C(net645),
    .Y(\reg_module/_07080_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14410_  (.A(\reg_module/_05287_ ),
    .X(\reg_module/_07081_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14411_  (.A(\reg_module/_07081_ ),
    .B(\reg_module/gprf[826] ),
    .Y(\reg_module/_07082_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14412_  (.A(\reg_module/gprf[794] ),
    .B(net780),
    .Y(\reg_module/_07083_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14413_  (.A(\reg_module/_07082_ ),
    .B(net699),
    .C(\reg_module/_07083_ ),
    .Y(\reg_module/_07084_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14414_  (.A(\reg_module/_07008_ ),
    .B(\reg_module/gprf[890] ),
    .Y(\reg_module/_07085_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14415_  (.A(\reg_module/gprf[858] ),
    .B(net777),
    .Y(\reg_module/_07086_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14416_  (.A(\reg_module/_07085_ ),
    .B(\reg_module/_06853_ ),
    .C(\reg_module/_07086_ ),
    .Y(\reg_module/_07087_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14417_  (.A(\reg_module/_07084_ ),
    .B(\reg_module/_07087_ ),
    .Y(\reg_module/_07088_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14418_  (.A(\reg_module/_07088_ ),
    .B(net660),
    .Y(\reg_module/_07089_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14419_  (.A(\reg_module/_06706_ ),
    .B(\reg_module/gprf[954] ),
    .Y(\reg_module/_07090_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14420_  (.A(\reg_module/gprf[922] ),
    .B(net791),
    .Y(\reg_module/_07091_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14421_  (.A(\reg_module/_07090_ ),
    .B(net708),
    .C(\reg_module/_07091_ ),
    .Y(\reg_module/_07092_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14422_  (.A(\reg_module/_06861_ ),
    .B(\reg_module/gprf[1018] ),
    .Y(\reg_module/_07093_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14423_  (.A(\reg_module/gprf[986] ),
    .B(net791),
    .Y(\reg_module/_07094_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14424_  (.A(\reg_module/_07093_ ),
    .B(\reg_module/_06940_ ),
    .C(\reg_module/_07094_ ),
    .Y(\reg_module/_07095_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14425_  (.A(\reg_module/_07092_ ),
    .B(\reg_module/_07095_ ),
    .Y(\reg_module/_07096_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14426_  (.A(\reg_module/_07096_ ),
    .B(\reg_module/_05362_ ),
    .Y(\reg_module/_07097_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14427_  (.A(\reg_module/_07089_ ),
    .B(\reg_module/_07097_ ),
    .C(\reg_module/_05538_ ),
    .Y(\reg_module/_07098_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14428_  (.A(\reg_module/_07080_ ),
    .B(\reg_module/_07098_ ),
    .Y(\reg_module/_07099_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14429_  (.A(\reg_module/_07099_ ),
    .B(\reg_module/_06717_ ),
    .Y(\reg_module/_07100_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14430_  (.A(\reg_module/_06793_ ),
    .B(\reg_module/gprf[314] ),
    .Y(\reg_module/_07101_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14431_  (.A(\reg_module/gprf[282] ),
    .B(net783),
    .Y(\reg_module/_07102_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14432_  (.A(\reg_module/_07101_ ),
    .B(net702),
    .C(\reg_module/_07102_ ),
    .Y(\reg_module/_07103_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14433_  (.A(\reg_module/_06888_ ),
    .B(\reg_module/gprf[378] ),
    .Y(\reg_module/_07104_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14434_  (.A(\reg_module/gprf[346] ),
    .B(net783),
    .Y(\reg_module/_07105_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14435_  (.A(\reg_module/_07104_ ),
    .B(\reg_module/_07029_ ),
    .C(\reg_module/_07105_ ),
    .Y(\reg_module/_07106_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14436_  (.A(\reg_module/_07103_ ),
    .B(\reg_module/_07106_ ),
    .Y(\reg_module/_07107_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14437_  (.A(\reg_module/_07107_ ),
    .B(net663),
    .Y(\reg_module/_07108_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14438_  (.A(\reg_module/_06878_ ),
    .B(\reg_module/gprf[442] ),
    .Y(\reg_module/_07109_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14439_  (.A(\reg_module/gprf[410] ),
    .B(net759),
    .Y(\reg_module/_07110_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14440_  (.A(\reg_module/_07109_ ),
    .B(net692),
    .C(\reg_module/_07110_ ),
    .Y(\reg_module/_07111_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14441_  (.A(\reg_module/_07037_ ),
    .B(\reg_module/gprf[506] ),
    .Y(\reg_module/_07112_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14442_  (.A(\reg_module/_05086_ ),
    .X(\reg_module/_07113_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14443_  (.A(\reg_module/gprf[474] ),
    .B(net759),
    .Y(\reg_module/_07114_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14444_  (.A(\reg_module/_07112_ ),
    .B(\reg_module/_07113_ ),
    .C(\reg_module/_07114_ ),
    .Y(\reg_module/_07115_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14445_  (.A(\reg_module/_07111_ ),
    .B(\reg_module/_07115_ ),
    .Y(\reg_module/_07116_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14446_  (.A(\reg_module/_07116_ ),
    .B(\reg_module/_07042_ ),
    .Y(\reg_module/_07117_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14447_  (.A(\reg_module/_07108_ ),
    .B(\reg_module/_07117_ ),
    .C(\reg_module/_06964_ ),
    .Y(\reg_module/_07118_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14448_  (.A(\reg_module/_05034_ ),
    .X(\reg_module/_07119_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14449_  (.A(\reg_module/_07119_ ),
    .B(\reg_module/gprf[58] ),
    .Y(\reg_module/_07120_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14450_  (.A(\reg_module/gprf[26] ),
    .B(net782),
    .Y(\reg_module/_07121_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14451_  (.A(\reg_module/_07120_ ),
    .B(net702),
    .C(\reg_module/_07121_ ),
    .Y(\reg_module/_07122_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14452_  (.A(\reg_module/_06892_ ),
    .B(\reg_module/gprf[122] ),
    .Y(\reg_module/_07123_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14453_  (.A(\reg_module/gprf[90] ),
    .B(net783),
    .Y(\reg_module/_07124_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14454_  (.A(\reg_module/_07123_ ),
    .B(\reg_module/_06815_ ),
    .C(\reg_module/_07124_ ),
    .Y(\reg_module/_07125_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14455_  (.A(\reg_module/_07122_ ),
    .B(\reg_module/_07125_ ),
    .Y(\reg_module/_07126_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14456_  (.A(\reg_module/_07126_ ),
    .B(net663),
    .Y(\reg_module/_07127_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14457_  (.A(\reg_module/_06744_ ),
    .B(\reg_module/gprf[186] ),
    .Y(\reg_module/_07128_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14458_  (.A(\reg_module/gprf[154] ),
    .B(net760),
    .Y(\reg_module/_07129_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14459_  (.A(\reg_module/_07128_ ),
    .B(net692),
    .C(\reg_module/_07129_ ),
    .Y(\reg_module/_07130_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14460_  (.A(\reg_module/_06748_ ),
    .B(\reg_module/gprf[250] ),
    .Y(\reg_module/_07131_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14461_  (.A(\reg_module/gprf[218] ),
    .B(net760),
    .Y(\reg_module/_07132_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14462_  (.A(\reg_module/_07131_ ),
    .B(\reg_module/_06824_ ),
    .C(\reg_module/_07132_ ),
    .Y(\reg_module/_07133_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14463_  (.A(\reg_module/_07130_ ),
    .B(\reg_module/_07133_ ),
    .Y(\reg_module/_07134_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14464_  (.A(\reg_module/_07134_ ),
    .B(\reg_module/_06981_ ),
    .Y(\reg_module/_07135_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14465_  (.A(\reg_module/_07127_ ),
    .B(\reg_module/_07135_ ),
    .C(net646),
    .Y(\reg_module/_07136_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14466_  (.A(\reg_module/_07118_ ),
    .B(\reg_module/_07136_ ),
    .Y(\reg_module/_07137_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14467_  (.A(\reg_module/_07137_ ),
    .B(net635),
    .Y(\reg_module/_07138_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14468_  (.A(\reg_module/_07100_ ),
    .B(\reg_module/_07138_ ),
    .Y(\wRs1Data[26] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14469_  (.A(\reg_module/_05003_ ),
    .B(\reg_module/gprf[827] ),
    .Y(\reg_module/_07139_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14470_  (.A(\reg_module/gprf[795] ),
    .B(net780),
    .Y(\reg_module/_07140_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14471_  (.A(\reg_module/_07139_ ),
    .B(net700),
    .C(\reg_module/_07140_ ),
    .Y(\reg_module/_07141_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14472_  (.A(\reg_module/_05014_ ),
    .B(\reg_module/gprf[891] ),
    .Y(\reg_module/_07142_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14473_  (.A(\reg_module/gprf[859] ),
    .B(net780),
    .Y(\reg_module/_07143_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14474_  (.A(\reg_module/_07142_ ),
    .B(\reg_module/_05073_ ),
    .C(\reg_module/_07143_ ),
    .Y(\reg_module/_07144_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14475_  (.A(\reg_module/_07141_ ),
    .B(\reg_module/_07144_ ),
    .Y(\reg_module/_07145_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14476_  (.A(\reg_module/_07145_ ),
    .B(net661),
    .Y(\reg_module/_07146_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14477_  (.A(\reg_module/_06994_ ),
    .B(\reg_module/gprf[955] ),
    .Y(\reg_module/_07147_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14478_  (.A(\reg_module/gprf[923] ),
    .B(net763),
    .Y(\reg_module/_07148_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14479_  (.A(\reg_module/_07147_ ),
    .B(net693),
    .C(\reg_module/_07148_ ),
    .Y(\reg_module/_07149_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14480_  (.A(\reg_module/_06998_ ),
    .B(\reg_module/gprf[1019] ),
    .Y(\reg_module/_07150_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14481_  (.A(\reg_module/gprf[987] ),
    .B(net762),
    .Y(\reg_module/_07151_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14482_  (.A(\reg_module/_07150_ ),
    .B(\reg_module/_04998_ ),
    .C(\reg_module/_07151_ ),
    .Y(\reg_module/_07152_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14483_  (.A(\reg_module/_07149_ ),
    .B(\reg_module/_07152_ ),
    .Y(\reg_module/_07153_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14484_  (.A(\reg_module/_07153_ ),
    .B(\reg_module/_06924_ ),
    .Y(\reg_module/_07154_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14485_  (.A(\reg_module/_07146_ ),
    .B(\reg_module/_07154_ ),
    .C(\reg_module/_06926_ ),
    .Y(\reg_module/_07155_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14486_  (.A(\reg_module/_07081_ ),
    .B(\reg_module/gprf[699] ),
    .Y(\reg_module/_07156_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14487_  (.A(\reg_module/gprf[667] ),
    .B(net777),
    .Y(\reg_module/_07157_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14488_  (.A(\reg_module/_07156_ ),
    .B(net700),
    .C(\reg_module/_07157_ ),
    .Y(\reg_module/_07158_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14489_  (.A(\reg_module/_07008_ ),
    .B(\reg_module/gprf[763] ),
    .Y(\reg_module/_07159_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14490_  (.A(\reg_module/gprf[731] ),
    .B(net777),
    .Y(\reg_module/_07160_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14491_  (.A(\reg_module/_07159_ ),
    .B(\reg_module/_06853_ ),
    .C(\reg_module/_07160_ ),
    .Y(\reg_module/_07161_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14492_  (.A(\reg_module/_07158_ ),
    .B(\reg_module/_07161_ ),
    .Y(\reg_module/_07162_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14493_  (.A(\reg_module/_07162_ ),
    .B(\reg_module/_06550_ ),
    .Y(\reg_module/_07163_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14494_  (.A(\reg_module/_05020_ ),
    .B(\reg_module/gprf[571] ),
    .Y(\reg_module/_07164_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14495_  (.A(\reg_module/gprf[539] ),
    .B(net777),
    .Y(\reg_module/_07165_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14496_  (.A(\reg_module/_07164_ ),
    .B(net698),
    .C(\reg_module/_07165_ ),
    .Y(\reg_module/_07166_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14497_  (.A(\reg_module/_06861_ ),
    .B(\reg_module/gprf[635] ),
    .Y(\reg_module/_07167_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14498_  (.A(\reg_module/gprf[603] ),
    .B(net778),
    .Y(\reg_module/_07168_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14499_  (.A(\reg_module/_07167_ ),
    .B(\reg_module/_06940_ ),
    .C(\reg_module/_07168_ ),
    .Y(\reg_module/_07169_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14500_  (.A(\reg_module/_07166_ ),
    .B(\reg_module/_07169_ ),
    .Y(\reg_module/_07170_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14501_  (.A(\reg_module/_07170_ ),
    .B(net660),
    .Y(\reg_module/_07171_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14502_  (.A(\reg_module/_07163_ ),
    .B(\reg_module/_07171_ ),
    .C(net641),
    .Y(\reg_module/_07172_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14503_  (.A(\reg_module/_07155_ ),
    .B(\reg_module/_07172_ ),
    .Y(\reg_module/_07173_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14504_  (.A(\reg_module/_07173_ ),
    .B(\reg_module/_05124_ ),
    .Y(\reg_module/_07174_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14505_  (.A(\reg_module/_06793_ ),
    .B(\reg_module/gprf[315] ),
    .Y(\reg_module/_07175_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14506_  (.A(\reg_module/gprf[283] ),
    .B(net759),
    .Y(\reg_module/_07176_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14507_  (.A(\reg_module/_07175_ ),
    .B(net691),
    .C(\reg_module/_07176_ ),
    .Y(\reg_module/_07177_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14508_  (.A(\reg_module/_07119_ ),
    .B(\reg_module/gprf[379] ),
    .Y(\reg_module/_07178_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14509_  (.A(\reg_module/gprf[347] ),
    .B(net759),
    .Y(\reg_module/_07179_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14510_  (.A(\reg_module/_07178_ ),
    .B(\reg_module/_07029_ ),
    .C(\reg_module/_07179_ ),
    .Y(\reg_module/_07180_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14511_  (.A(\reg_module/_07177_ ),
    .B(\reg_module/_07180_ ),
    .Y(\reg_module/_07181_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14512_  (.A(\reg_module/_07181_ ),
    .B(net657),
    .Y(\reg_module/_07182_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14513_  (.A(\reg_module/_06878_ ),
    .B(\reg_module/gprf[443] ),
    .Y(\reg_module/_07183_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14514_  (.A(\reg_module/gprf[411] ),
    .B(net759),
    .Y(\reg_module/_07184_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14515_  (.A(\reg_module/_07183_ ),
    .B(net692),
    .C(\reg_module/_07184_ ),
    .Y(\reg_module/_07185_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14516_  (.A(\reg_module/_07037_ ),
    .B(\reg_module/gprf[507] ),
    .Y(\reg_module/_07186_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14517_  (.A(\reg_module/gprf[475] ),
    .B(net759),
    .Y(\reg_module/_07187_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14518_  (.A(\reg_module/_07186_ ),
    .B(\reg_module/_07113_ ),
    .C(\reg_module/_07187_ ),
    .Y(\reg_module/_07188_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14519_  (.A(\reg_module/_07185_ ),
    .B(\reg_module/_07188_ ),
    .Y(\reg_module/_07189_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14520_  (.A(\reg_module/_07189_ ),
    .B(\reg_module/_07042_ ),
    .Y(\reg_module/_07190_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14521_  (.A(\reg_module/_07182_ ),
    .B(\reg_module/_07190_ ),
    .C(\reg_module/_06964_ ),
    .Y(\reg_module/_07191_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14522_  (.A(\reg_module/_07119_ ),
    .B(\reg_module/gprf[59] ),
    .Y(\reg_module/_07192_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14523_  (.A(\reg_module/gprf[27] ),
    .B(net760),
    .Y(\reg_module/_07193_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14524_  (.A(\reg_module/_07192_ ),
    .B(net692),
    .C(\reg_module/_07193_ ),
    .Y(\reg_module/_07194_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14525_  (.A(\reg_module/_06892_ ),
    .B(\reg_module/gprf[123] ),
    .Y(\reg_module/_07195_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14526_  (.A(\reg_module/gprf[91] ),
    .B(net761),
    .Y(\reg_module/_07196_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14527_  (.A(\reg_module/_07195_ ),
    .B(\reg_module/_06815_ ),
    .C(\reg_module/_07196_ ),
    .Y(\reg_module/_07197_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14528_  (.A(\reg_module/_07194_ ),
    .B(\reg_module/_07197_ ),
    .Y(\reg_module/_07198_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14529_  (.A(\reg_module/_07198_ ),
    .B(net657),
    .Y(\reg_module/_07199_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14530_  (.A(\reg_module/_05084_ ),
    .B(\reg_module/gprf[187] ),
    .Y(\reg_module/_07200_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14531_  (.A(\reg_module/gprf[155] ),
    .B(net760),
    .Y(\reg_module/_07201_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14532_  (.A(\reg_module/_07200_ ),
    .B(net692),
    .C(\reg_module/_07201_ ),
    .Y(\reg_module/_07202_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14533_  (.A(\reg_module/_05282_ ),
    .B(\reg_module/gprf[251] ),
    .Y(\reg_module/_07203_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14534_  (.A(\reg_module/gprf[219] ),
    .B(net760),
    .Y(\reg_module/_07204_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14535_  (.A(\reg_module/_07203_ ),
    .B(\reg_module/_06824_ ),
    .C(\reg_module/_07204_ ),
    .Y(\reg_module/_07205_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14536_  (.A(\reg_module/_07202_ ),
    .B(\reg_module/_07205_ ),
    .Y(\reg_module/_07206_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14537_  (.A(\reg_module/_07206_ ),
    .B(\reg_module/_06981_ ),
    .Y(\reg_module/_07207_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14538_  (.A(\reg_module/_07199_ ),
    .B(\reg_module/_07207_ ),
    .C(net642),
    .Y(\reg_module/_07208_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14539_  (.A(\reg_module/_07191_ ),
    .B(\reg_module/_07208_ ),
    .Y(\reg_module/_07209_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14540_  (.A(\reg_module/_07209_ ),
    .B(net635),
    .Y(\reg_module/_07210_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_14541_  (.A(\reg_module/_07174_ ),
    .B(\reg_module/_07210_ ),
    .Y(\wRs1Data[27] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14542_  (.A(\reg_module/_05003_ ),
    .B(\reg_module/gprf[828] ),
    .Y(\reg_module/_07211_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14543_  (.A(\reg_module/gprf[796] ),
    .B(net779),
    .Y(\reg_module/_07212_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14544_  (.A(\reg_module/_07211_ ),
    .B(net699),
    .C(\reg_module/_07212_ ),
    .Y(\reg_module/_07213_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14545_  (.A(\reg_module/_05014_ ),
    .B(\reg_module/gprf[892] ),
    .Y(\reg_module/_07214_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14546_  (.A(\reg_module/gprf[860] ),
    .B(net779),
    .Y(\reg_module/_07215_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14547_  (.A(\reg_module/_07214_ ),
    .B(\reg_module/_05073_ ),
    .C(\reg_module/_07215_ ),
    .Y(\reg_module/_07216_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14548_  (.A(\reg_module/_07213_ ),
    .B(\reg_module/_07216_ ),
    .Y(\reg_module/_07217_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14549_  (.A(\reg_module/_07217_ ),
    .B(net660),
    .Y(\reg_module/_07218_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14550_  (.A(\reg_module/_06994_ ),
    .B(\reg_module/gprf[956] ),
    .Y(\reg_module/_07219_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14551_  (.A(\reg_module/gprf[924] ),
    .B(net762),
    .Y(\reg_module/_07220_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14552_  (.A(\reg_module/_07219_ ),
    .B(net693),
    .C(\reg_module/_07220_ ),
    .Y(\reg_module/_07221_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14553_  (.A(\reg_module/_06998_ ),
    .B(\reg_module/gprf[1020] ),
    .Y(\reg_module/_07222_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14554_  (.A(\reg_module/gprf[988] ),
    .B(net762),
    .Y(\reg_module/_07223_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14555_  (.A(\reg_module/_07222_ ),
    .B(\reg_module/_04998_ ),
    .C(\reg_module/_07223_ ),
    .Y(\reg_module/_07224_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14556_  (.A(\reg_module/_07221_ ),
    .B(\reg_module/_07224_ ),
    .Y(\reg_module/_07225_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14557_  (.A(\reg_module/_07225_ ),
    .B(\reg_module/_06924_ ),
    .Y(\reg_module/_07226_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14558_  (.A(\reg_module/_07218_ ),
    .B(\reg_module/_07226_ ),
    .C(\reg_module/_06926_ ),
    .Y(\reg_module/_07227_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14559_  (.A(\reg_module/_07081_ ),
    .B(\reg_module/gprf[700] ),
    .Y(\reg_module/_07228_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14560_  (.A(\reg_module/gprf[668] ),
    .B(net775),
    .Y(\reg_module/_07229_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14561_  (.A(\reg_module/_07228_ ),
    .B(net698),
    .C(\reg_module/_07229_ ),
    .Y(\reg_module/_07230_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14562_  (.A(\reg_module/_07008_ ),
    .B(\reg_module/gprf[764] ),
    .Y(\reg_module/_07231_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14563_  (.A(\reg_module/gprf[732] ),
    .B(net775),
    .Y(\reg_module/_07232_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14564_  (.A(\reg_module/_07231_ ),
    .B(\reg_module/_06853_ ),
    .C(\reg_module/_07232_ ),
    .Y(\reg_module/_07233_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14565_  (.A(\reg_module/_07230_ ),
    .B(\reg_module/_07233_ ),
    .Y(\reg_module/_07234_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14566_  (.A(\reg_module/_07234_ ),
    .B(\reg_module/_05304_ ),
    .Y(\reg_module/_07235_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14567_  (.A(\reg_module/_05020_ ),
    .B(\reg_module/gprf[572] ),
    .Y(\reg_module/_07236_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14568_  (.A(\reg_module/gprf[540] ),
    .B(net776),
    .Y(\reg_module/_07237_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14569_  (.A(\reg_module/_07236_ ),
    .B(net698),
    .C(\reg_module/_07237_ ),
    .Y(\reg_module/_07238_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14570_  (.A(\reg_module/_06861_ ),
    .B(\reg_module/gprf[636] ),
    .Y(\reg_module/_07239_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14571_  (.A(\reg_module/gprf[604] ),
    .B(net775),
    .Y(\reg_module/_07240_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14572_  (.A(\reg_module/_07239_ ),
    .B(\reg_module/_06940_ ),
    .C(\reg_module/_07240_ ),
    .Y(\reg_module/_07241_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14573_  (.A(\reg_module/_07238_ ),
    .B(\reg_module/_07241_ ),
    .Y(\reg_module/_07242_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14574_  (.A(\reg_module/_07242_ ),
    .B(net659),
    .Y(\reg_module/_07243_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14575_  (.A(\reg_module/_07235_ ),
    .B(\reg_module/_07243_ ),
    .C(net640),
    .Y(\reg_module/_07244_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14576_  (.A(\reg_module/_07227_ ),
    .B(\reg_module/_07244_ ),
    .Y(\reg_module/_07245_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14577_  (.A(\reg_module/_07245_ ),
    .B(\reg_module/_05124_ ),
    .Y(\reg_module/_07246_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14578_  (.A(\reg_module/_05030_ ),
    .B(\reg_module/gprf[316] ),
    .Y(\reg_module/_07247_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14579_  (.A(\reg_module/gprf[284] ),
    .B(net762),
    .Y(\reg_module/_07248_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14580_  (.A(\reg_module/_07247_ ),
    .B(net693),
    .C(\reg_module/_07248_ ),
    .Y(\reg_module/_07249_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14581_  (.A(\reg_module/_07119_ ),
    .B(\reg_module/gprf[380] ),
    .Y(\reg_module/_07250_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14582_  (.A(\reg_module/gprf[348] ),
    .B(net758),
    .Y(\reg_module/_07251_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14583_  (.A(\reg_module/_07250_ ),
    .B(\reg_module/_07029_ ),
    .C(\reg_module/_07251_ ),
    .Y(\reg_module/_07252_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14584_  (.A(\reg_module/_07249_ ),
    .B(\reg_module/_07252_ ),
    .Y(\reg_module/_07253_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14585_  (.A(\reg_module/_07253_ ),
    .B(net657),
    .Y(\reg_module/_07254_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14586_  (.A(\reg_module/_06878_ ),
    .B(\reg_module/gprf[444] ),
    .Y(\reg_module/_07255_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14587_  (.A(\reg_module/gprf[412] ),
    .B(net758),
    .Y(\reg_module/_07256_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14588_  (.A(\reg_module/_07255_ ),
    .B(net691),
    .C(\reg_module/_07256_ ),
    .Y(\reg_module/_07257_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14589_  (.A(\reg_module/_07037_ ),
    .B(\reg_module/gprf[508] ),
    .Y(\reg_module/_07258_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14590_  (.A(\reg_module/gprf[476] ),
    .B(net758),
    .Y(\reg_module/_07259_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14591_  (.A(\reg_module/_07258_ ),
    .B(\reg_module/_07113_ ),
    .C(\reg_module/_07259_ ),
    .Y(\reg_module/_07260_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14592_  (.A(\reg_module/_07257_ ),
    .B(\reg_module/_07260_ ),
    .Y(\reg_module/_07261_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14593_  (.A(\reg_module/_07261_ ),
    .B(\reg_module/_07042_ ),
    .Y(\reg_module/_07262_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14594_  (.A(\reg_module/_07254_ ),
    .B(\reg_module/_07262_ ),
    .C(\reg_module/_06964_ ),
    .Y(\reg_module/_07263_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14595_  (.A(\reg_module/_07119_ ),
    .B(\reg_module/gprf[60] ),
    .Y(\reg_module/_07264_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14596_  (.A(\reg_module/gprf[28] ),
    .B(net757),
    .Y(\reg_module/_07265_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14597_  (.A(\reg_module/_07264_ ),
    .B(net691),
    .C(\reg_module/_07265_ ),
    .Y(\reg_module/_07266_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14598_  (.A(\reg_module/_06892_ ),
    .B(\reg_module/gprf[124] ),
    .Y(\reg_module/_07267_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14599_  (.A(\reg_module/gprf[92] ),
    .B(net758),
    .Y(\reg_module/_07268_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14600_  (.A(\reg_module/_07267_ ),
    .B(\reg_module/_05087_ ),
    .C(\reg_module/_07268_ ),
    .Y(\reg_module/_07269_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14601_  (.A(\reg_module/_07266_ ),
    .B(\reg_module/_07269_ ),
    .Y(\reg_module/_07270_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14602_  (.A(\reg_module/_07270_ ),
    .B(net656),
    .Y(\reg_module/_07271_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14603_  (.A(\reg_module/_05084_ ),
    .B(\reg_module/gprf[188] ),
    .Y(\reg_module/_07272_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14604_  (.A(\reg_module/gprf[156] ),
    .B(net757),
    .Y(\reg_module/_07273_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14605_  (.A(\reg_module/_07272_ ),
    .B(net691),
    .C(\reg_module/_07273_ ),
    .Y(\reg_module/_07274_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14606_  (.A(\reg_module/_05282_ ),
    .B(\reg_module/gprf[252] ),
    .Y(\reg_module/_07275_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14607_  (.A(\reg_module/gprf[220] ),
    .B(net757),
    .Y(\reg_module/_07276_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14608_  (.A(\reg_module/_07275_ ),
    .B(\reg_module/_05290_ ),
    .C(\reg_module/_07276_ ),
    .Y(\reg_module/_07277_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14609_  (.A(\reg_module/_07274_ ),
    .B(\reg_module/_07277_ ),
    .Y(\reg_module/_07278_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14610_  (.A(\reg_module/_07278_ ),
    .B(\reg_module/_06981_ ),
    .Y(\reg_module/_07279_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14611_  (.A(\reg_module/_07271_ ),
    .B(\reg_module/_07279_ ),
    .C(net642),
    .Y(\reg_module/_07280_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14612_  (.A(\reg_module/_07263_ ),
    .B(\reg_module/_07280_ ),
    .Y(\reg_module/_07281_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14613_  (.A(\reg_module/_07281_ ),
    .B(net632),
    .Y(\reg_module/_07282_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_14614_  (.A(\reg_module/_07246_ ),
    .B(\reg_module/_07282_ ),
    .Y(\wRs1Data[28] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14615_  (.A(\reg_module/_05003_ ),
    .B(\reg_module/gprf[573] ),
    .Y(\reg_module/_07283_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14616_  (.A(\reg_module/gprf[541] ),
    .B(net775),
    .Y(\reg_module/_07284_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14617_  (.A(\reg_module/_07283_ ),
    .B(net698),
    .C(\reg_module/_07284_ ),
    .Y(\reg_module/_07285_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14618_  (.A(\reg_module/_05014_ ),
    .B(\reg_module/gprf[637] ),
    .Y(\reg_module/_07286_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14619_  (.A(\reg_module/gprf[605] ),
    .B(net776),
    .Y(\reg_module/_07287_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14620_  (.A(\reg_module/_07286_ ),
    .B(\reg_module/_05073_ ),
    .C(\reg_module/_07287_ ),
    .Y(\reg_module/_07288_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14621_  (.A(\reg_module/_07285_ ),
    .B(\reg_module/_07288_ ),
    .Y(\reg_module/_07289_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14622_  (.A(\reg_module/_07289_ ),
    .B(net660),
    .Y(\reg_module/_07290_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14623_  (.A(\reg_module/_06994_ ),
    .B(\reg_module/gprf[701] ),
    .Y(\reg_module/_07291_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14624_  (.A(\reg_module/gprf[669] ),
    .B(net775),
    .Y(\reg_module/_07292_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14625_  (.A(\reg_module/_07291_ ),
    .B(net698),
    .C(\reg_module/_07292_ ),
    .Y(\reg_module/_07293_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14626_  (.A(\reg_module/_06998_ ),
    .B(\reg_module/gprf[765] ),
    .Y(\reg_module/_07294_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14627_  (.A(\reg_module/gprf[733] ),
    .B(net762),
    .Y(\reg_module/_07295_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14628_  (.A(\reg_module/_07294_ ),
    .B(\reg_module/_04998_ ),
    .C(\reg_module/_07295_ ),
    .Y(\reg_module/_07296_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14629_  (.A(\reg_module/_07293_ ),
    .B(\reg_module/_07296_ ),
    .Y(\reg_module/_07297_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14630_  (.A(\reg_module/_07297_ ),
    .B(\reg_module/_06924_ ),
    .Y(\reg_module/_07298_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14631_  (.A(\reg_module/_07290_ ),
    .B(\reg_module/_07298_ ),
    .C(net641),
    .Y(\reg_module/_07299_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14632_  (.A(\reg_module/_07081_ ),
    .B(\reg_module/gprf[829] ),
    .Y(\reg_module/_07300_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14633_  (.A(\reg_module/gprf[797] ),
    .B(net779),
    .Y(\reg_module/_07301_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14634_  (.A(\reg_module/_07300_ ),
    .B(net699),
    .C(\reg_module/_07301_ ),
    .Y(\reg_module/_07302_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14635_  (.A(\reg_module/_07008_ ),
    .B(\reg_module/gprf[893] ),
    .Y(\reg_module/_07303_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14636_  (.A(\reg_module/gprf[861] ),
    .B(net776),
    .Y(\reg_module/_07304_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14637_  (.A(\reg_module/_07303_ ),
    .B(\reg_module/_05023_ ),
    .C(\reg_module/_07304_ ),
    .Y(\reg_module/_07305_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14638_  (.A(\reg_module/_07302_ ),
    .B(\reg_module/_07305_ ),
    .Y(\reg_module/_07306_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14639_  (.A(\reg_module/_07306_ ),
    .B(net660),
    .Y(\reg_module/_07307_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14640_  (.A(\reg_module/_05020_ ),
    .B(\reg_module/gprf[957] ),
    .Y(\reg_module/_07308_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14641_  (.A(\reg_module/gprf[925] ),
    .B(net775),
    .Y(\reg_module/_07309_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14642_  (.A(\reg_module/_07308_ ),
    .B(net698),
    .C(\reg_module/_07309_ ),
    .Y(\reg_module/_07310_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14643_  (.A(\reg_module/_05114_ ),
    .B(\reg_module/gprf[1021] ),
    .Y(\reg_module/_07311_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14644_  (.A(\reg_module/gprf[989] ),
    .B(net767),
    .Y(\reg_module/_07312_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14645_  (.A(\reg_module/_07311_ ),
    .B(\reg_module/_06940_ ),
    .C(\reg_module/_07312_ ),
    .Y(\reg_module/_07313_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14646_  (.A(\reg_module/_07310_ ),
    .B(\reg_module/_07313_ ),
    .Y(\reg_module/_07314_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14647_  (.A(\reg_module/_07314_ ),
    .B(\reg_module/_05362_ ),
    .Y(\reg_module/_07315_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14648_  (.A(\reg_module/_07307_ ),
    .B(\reg_module/_07315_ ),
    .C(\reg_module/_05538_ ),
    .Y(\reg_module/_07316_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14649_  (.A(\reg_module/_07299_ ),
    .B(\reg_module/_07316_ ),
    .Y(\reg_module/_07317_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14650_  (.A(\reg_module/_07317_ ),
    .B(\reg_module/_05124_ ),
    .Y(\reg_module/_07318_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14651_  (.A(\reg_module/_05030_ ),
    .B(\reg_module/gprf[317] ),
    .Y(\reg_module/_07319_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14652_  (.A(\reg_module/gprf[285] ),
    .B(net762),
    .Y(\reg_module/_07320_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14653_  (.A(\reg_module/_07319_ ),
    .B(net693),
    .C(\reg_module/_07320_ ),
    .Y(\reg_module/_07321_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14654_  (.A(\reg_module/_07119_ ),
    .B(\reg_module/gprf[381] ),
    .Y(\reg_module/_07322_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14655_  (.A(\reg_module/gprf[349] ),
    .B(net758),
    .Y(\reg_module/_07323_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14656_  (.A(\reg_module/_07322_ ),
    .B(\reg_module/_07029_ ),
    .C(\reg_module/_07323_ ),
    .Y(\reg_module/_07324_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14657_  (.A(\reg_module/_07321_ ),
    .B(\reg_module/_07324_ ),
    .Y(\reg_module/_07325_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14658_  (.A(\reg_module/_07325_ ),
    .B(net657),
    .Y(\reg_module/_07326_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14659_  (.A(\reg_module/_05044_ ),
    .B(\reg_module/gprf[445] ),
    .Y(\reg_module/_07327_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14660_  (.A(\reg_module/gprf[413] ),
    .B(net757),
    .Y(\reg_module/_07328_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14661_  (.A(\reg_module/_07327_ ),
    .B(net691),
    .C(\reg_module/_07328_ ),
    .Y(\reg_module/_07329_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14662_  (.A(\reg_module/_07037_ ),
    .B(\reg_module/gprf[509] ),
    .Y(\reg_module/_07330_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14663_  (.A(\reg_module/gprf[477] ),
    .B(net758),
    .Y(\reg_module/_07331_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14664_  (.A(\reg_module/_07330_ ),
    .B(\reg_module/_07113_ ),
    .C(\reg_module/_07331_ ),
    .Y(\reg_module/_07332_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14665_  (.A(\reg_module/_07329_ ),
    .B(\reg_module/_07332_ ),
    .Y(\reg_module/_07333_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14666_  (.A(\reg_module/_07333_ ),
    .B(\reg_module/_07042_ ),
    .Y(\reg_module/_07334_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14667_  (.A(\reg_module/_07326_ ),
    .B(\reg_module/_07334_ ),
    .C(\reg_module/_06964_ ),
    .Y(\reg_module/_07335_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14668_  (.A(\reg_module/_05035_ ),
    .B(\reg_module/gprf[61] ),
    .Y(\reg_module/_07336_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14669_  (.A(\reg_module/gprf[29] ),
    .B(net756),
    .Y(\reg_module/_07337_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14670_  (.A(\reg_module/_07336_ ),
    .B(net690),
    .C(\reg_module/_07337_ ),
    .Y(\reg_module/_07338_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14671_  (.A(\reg_module/_05109_ ),
    .B(\reg_module/gprf[125] ),
    .Y(\reg_module/_07339_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14672_  (.A(\reg_module/gprf[93] ),
    .B(net756),
    .Y(\reg_module/_07340_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14673_  (.A(\reg_module/_07339_ ),
    .B(\reg_module/_05087_ ),
    .C(\reg_module/_07340_ ),
    .Y(\reg_module/_07341_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14674_  (.A(\reg_module/_07338_ ),
    .B(\reg_module/_07341_ ),
    .Y(\reg_module/_07342_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14675_  (.A(\reg_module/_07342_ ),
    .B(net656),
    .Y(\reg_module/_07343_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14676_  (.A(\reg_module/_05084_ ),
    .B(\reg_module/gprf[189] ),
    .Y(\reg_module/_07344_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14677_  (.A(\reg_module/gprf[157] ),
    .B(net757),
    .Y(\reg_module/_07345_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14678_  (.A(\reg_module/_07344_ ),
    .B(net691),
    .C(\reg_module/_07345_ ),
    .Y(\reg_module/_07346_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14679_  (.A(\reg_module/_05282_ ),
    .B(\reg_module/gprf[253] ),
    .Y(\reg_module/_07347_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14680_  (.A(\reg_module/gprf[221] ),
    .B(net757),
    .Y(\reg_module/_07348_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14681_  (.A(\reg_module/_07347_ ),
    .B(\reg_module/_05290_ ),
    .C(\reg_module/_07348_ ),
    .Y(\reg_module/_07349_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14682_  (.A(\reg_module/_07346_ ),
    .B(\reg_module/_07349_ ),
    .Y(\reg_module/_07350_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14683_  (.A(\reg_module/_07350_ ),
    .B(\reg_module/_06981_ ),
    .Y(\reg_module/_07351_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14684_  (.A(\reg_module/_07343_ ),
    .B(\reg_module/_07351_ ),
    .C(net642),
    .Y(\reg_module/_07352_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14685_  (.A(\reg_module/_07335_ ),
    .B(\reg_module/_07352_ ),
    .Y(\reg_module/_07353_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14686_  (.A(\reg_module/_07353_ ),
    .B(net632),
    .Y(\reg_module/_07354_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_14687_  (.A(\reg_module/_07318_ ),
    .B(\reg_module/_07354_ ),
    .Y(\wRs1Data[29] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14688_  (.A(\reg_module/_05003_ ),
    .B(\reg_module/gprf[830] ),
    .Y(\reg_module/_07355_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14689_  (.A(\reg_module/gprf[798] ),
    .B(net767),
    .Y(\reg_module/_07356_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14690_  (.A(\reg_module/_07355_ ),
    .B(net697),
    .C(\reg_module/_07356_ ),
    .Y(\reg_module/_07357_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14691_  (.A(\reg_module/_05014_ ),
    .B(\reg_module/gprf[894] ),
    .Y(\reg_module/_07358_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14692_  (.A(\reg_module/gprf[862] ),
    .B(net774),
    .Y(\reg_module/_07359_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14693_  (.A(\reg_module/_07358_ ),
    .B(\reg_module/_05073_ ),
    .C(\reg_module/_07359_ ),
    .Y(\reg_module/_07360_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14694_  (.A(\reg_module/_07357_ ),
    .B(\reg_module/_07360_ ),
    .Y(\reg_module/_07361_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14695_  (.A(\reg_module/_07361_ ),
    .B(net659),
    .Y(\reg_module/_07362_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14696_  (.A(\reg_module/_06994_ ),
    .B(\reg_module/gprf[958] ),
    .Y(\reg_module/_07363_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14697_  (.A(\reg_module/gprf[926] ),
    .B(net765),
    .Y(\reg_module/_07364_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14698_  (.A(\reg_module/_07363_ ),
    .B(net694),
    .C(\reg_module/_07364_ ),
    .Y(\reg_module/_07365_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14699_  (.A(\reg_module/_06998_ ),
    .B(\reg_module/gprf[1022] ),
    .Y(\reg_module/_07366_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14700_  (.A(\reg_module/gprf[990] ),
    .B(net765),
    .Y(\reg_module/_07367_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14701_  (.A(\reg_module/_07366_ ),
    .B(\reg_module/_04998_ ),
    .C(\reg_module/_07367_ ),
    .Y(\reg_module/_07368_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14702_  (.A(\reg_module/_07365_ ),
    .B(\reg_module/_07368_ ),
    .Y(\reg_module/_07369_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14703_  (.A(\reg_module/_07369_ ),
    .B(\reg_module/_05092_ ),
    .Y(\reg_module/_07370_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14704_  (.A(\reg_module/_07362_ ),
    .B(\reg_module/_07370_ ),
    .C(\reg_module/_06926_ ),
    .Y(\reg_module/_07371_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14705_  (.A(\reg_module/_07081_ ),
    .B(\reg_module/gprf[702] ),
    .Y(\reg_module/_07372_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14706_  (.A(\reg_module/gprf[670] ),
    .B(net765),
    .Y(\reg_module/_07373_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14707_  (.A(\reg_module/_07372_ ),
    .B(net694),
    .C(\reg_module/_07373_ ),
    .Y(\reg_module/_07374_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14708_  (.A(\reg_module/_07008_ ),
    .B(\reg_module/gprf[766] ),
    .Y(\reg_module/_07375_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14709_  (.A(\reg_module/gprf[734] ),
    .B(net765),
    .Y(\reg_module/_07376_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14710_  (.A(\reg_module/_07375_ ),
    .B(\reg_module/_05023_ ),
    .C(\reg_module/_07376_ ),
    .Y(\reg_module/_07377_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14711_  (.A(\reg_module/_07374_ ),
    .B(\reg_module/_07377_ ),
    .Y(\reg_module/_07378_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14712_  (.A(\reg_module/_07378_ ),
    .B(\reg_module/_05304_ ),
    .Y(\reg_module/_07379_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14713_  (.A(\reg_module/_05020_ ),
    .B(\reg_module/gprf[574] ),
    .Y(\reg_module/_07380_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14714_  (.A(\reg_module/gprf[542] ),
    .B(net765),
    .Y(\reg_module/_07381_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14715_  (.A(\reg_module/_07380_ ),
    .B(net694),
    .C(\reg_module/_07381_ ),
    .Y(\reg_module/_07382_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14716_  (.A(\reg_module/_05114_ ),
    .B(\reg_module/gprf[638] ),
    .Y(\reg_module/_07383_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14717_  (.A(\reg_module/gprf[606] ),
    .B(net767),
    .Y(\reg_module/_07384_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14718_  (.A(\reg_module/_07383_ ),
    .B(\reg_module/_05116_ ),
    .C(\reg_module/_07384_ ),
    .Y(\reg_module/_07385_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14719_  (.A(\reg_module/_07382_ ),
    .B(\reg_module/_07385_ ),
    .Y(\reg_module/_07386_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14720_  (.A(\reg_module/_07386_ ),
    .B(net659),
    .Y(\reg_module/_07387_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14721_  (.A(\reg_module/_07379_ ),
    .B(\reg_module/_07387_ ),
    .C(net640),
    .Y(\reg_module/_07388_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14722_  (.A(\reg_module/_07371_ ),
    .B(\reg_module/_07388_ ),
    .Y(\reg_module/_07389_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14723_  (.A(\reg_module/_07389_ ),
    .B(\reg_module/_05124_ ),
    .Y(\reg_module/_07390_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14724_  (.A(\reg_module/_05030_ ),
    .B(\reg_module/gprf[318] ),
    .Y(\reg_module/_07391_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14725_  (.A(\reg_module/gprf[286] ),
    .B(net754),
    .Y(\reg_module/_07392_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14726_  (.A(\reg_module/_07391_ ),
    .B(net690),
    .C(\reg_module/_07392_ ),
    .Y(\reg_module/_07393_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14727_  (.A(\reg_module/_05035_ ),
    .B(\reg_module/gprf[382] ),
    .Y(\reg_module/_07394_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14728_  (.A(\reg_module/gprf[350] ),
    .B(net754),
    .Y(\reg_module/_07395_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14729_  (.A(\reg_module/_07394_ ),
    .B(\reg_module/_07029_ ),
    .C(\reg_module/_07395_ ),
    .Y(\reg_module/_07396_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14730_  (.A(\reg_module/_07393_ ),
    .B(\reg_module/_07396_ ),
    .Y(\reg_module/_07397_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14731_  (.A(\reg_module/_07397_ ),
    .B(net656),
    .Y(\reg_module/_07398_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14732_  (.A(\reg_module/_05044_ ),
    .B(\reg_module/gprf[446] ),
    .Y(\reg_module/_07399_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14733_  (.A(\reg_module/gprf[414] ),
    .B(net756),
    .Y(\reg_module/_07400_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14734_  (.A(\reg_module/_07399_ ),
    .B(net690),
    .C(\reg_module/_07400_ ),
    .Y(\reg_module/_07401_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14735_  (.A(\reg_module/_07037_ ),
    .B(\reg_module/gprf[510] ),
    .Y(\reg_module/_07402_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14736_  (.A(\reg_module/gprf[478] ),
    .B(net756),
    .Y(\reg_module/_07403_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14737_  (.A(\reg_module/_07402_ ),
    .B(\reg_module/_07113_ ),
    .C(\reg_module/_07403_ ),
    .Y(\reg_module/_07404_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14738_  (.A(\reg_module/_07401_ ),
    .B(\reg_module/_07404_ ),
    .Y(\reg_module/_07405_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14739_  (.A(\reg_module/_07405_ ),
    .B(\reg_module/_07042_ ),
    .Y(\reg_module/_07406_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14740_  (.A(\reg_module/_07398_ ),
    .B(\reg_module/_07406_ ),
    .C(\reg_module/_05060_ ),
    .Y(\reg_module/_07407_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14741_  (.A(\reg_module/_05035_ ),
    .B(\reg_module/gprf[62] ),
    .Y(\reg_module/_07408_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14742_  (.A(\reg_module/gprf[30] ),
    .B(net755),
    .Y(\reg_module/_07409_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14743_  (.A(\reg_module/_07408_ ),
    .B(net689),
    .C(\reg_module/_07409_ ),
    .Y(\reg_module/_07410_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14744_  (.A(\reg_module/_05109_ ),
    .B(\reg_module/gprf[126] ),
    .Y(\reg_module/_07411_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14745_  (.A(\reg_module/gprf[94] ),
    .B(net756),
    .Y(\reg_module/_07412_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14746_  (.A(\reg_module/_07411_ ),
    .B(\reg_module/_05087_ ),
    .C(\reg_module/_07412_ ),
    .Y(\reg_module/_07413_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14747_  (.A(\reg_module/_07410_ ),
    .B(\reg_module/_07413_ ),
    .Y(\reg_module/_07414_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14748_  (.A(\reg_module/_07414_ ),
    .B(net656),
    .Y(\reg_module/_07415_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14749_  (.A(\reg_module/_05084_ ),
    .B(\reg_module/gprf[190] ),
    .Y(\reg_module/_07416_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14750_  (.A(\reg_module/gprf[158] ),
    .B(net755),
    .Y(\reg_module/_07417_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14751_  (.A(\reg_module/_07416_ ),
    .B(net689),
    .C(\reg_module/_07417_ ),
    .Y(\reg_module/_07418_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14752_  (.A(\reg_module/_05282_ ),
    .B(\reg_module/gprf[254] ),
    .Y(\reg_module/_07419_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14753_  (.A(\reg_module/gprf[222] ),
    .B(net755),
    .Y(\reg_module/_07420_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14754_  (.A(\reg_module/_07419_ ),
    .B(\reg_module/_05290_ ),
    .C(\reg_module/_07420_ ),
    .Y(\reg_module/_07421_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14755_  (.A(\reg_module/_07418_ ),
    .B(\reg_module/_07421_ ),
    .Y(\reg_module/_07422_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14756_  (.A(\reg_module/_07422_ ),
    .B(\reg_module/_05010_ ),
    .Y(\reg_module/_07423_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14757_  (.A(\reg_module/_07415_ ),
    .B(\reg_module/_07423_ ),
    .C(net642),
    .Y(\reg_module/_07424_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14758_  (.A(\reg_module/_07407_ ),
    .B(\reg_module/_07424_ ),
    .Y(\reg_module/_07425_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14759_  (.A(\reg_module/_07425_ ),
    .B(net632),
    .Y(\reg_module/_07426_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_14760_  (.A(\reg_module/_07390_ ),
    .B(\reg_module/_07426_ ),
    .Y(\wRs1Data[30] ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14761_  (.A(\reg_module/_05003_ ),
    .B(\reg_module/gprf[831] ),
    .Y(\reg_module/_07427_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14762_  (.A(\reg_module/gprf[799] ),
    .B(net771),
    .Y(\reg_module/_07428_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14763_  (.A(\reg_module/_07427_ ),
    .B(net696),
    .C(\reg_module/_07428_ ),
    .Y(\reg_module/_07429_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14764_  (.A(\reg_module/_05014_ ),
    .B(\reg_module/gprf[895] ),
    .Y(\reg_module/_07430_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14765_  (.A(\reg_module/gprf[863] ),
    .B(net767),
    .Y(\reg_module/_07431_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14766_  (.A(\reg_module/_07430_ ),
    .B(\reg_module/_05073_ ),
    .C(\reg_module/_07431_ ),
    .Y(\reg_module/_07432_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14767_  (.A(\reg_module/_07429_ ),
    .B(\reg_module/_07432_ ),
    .Y(\reg_module/_07433_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14768_  (.A(\reg_module/_07433_ ),
    .B(net659),
    .Y(\reg_module/_07434_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14769_  (.A(\reg_module/_05069_ ),
    .B(\reg_module/gprf[959] ),
    .Y(\reg_module/_07435_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14770_  (.A(\reg_module/gprf[927] ),
    .B(net766),
    .Y(\reg_module/_07436_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14771_  (.A(\reg_module/_07435_ ),
    .B(net694),
    .C(\reg_module/_07436_ ),
    .Y(\reg_module/_07437_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14772_  (.A(\reg_module/_05101_ ),
    .B(\reg_module/gprf[1023] ),
    .Y(\reg_module/_07438_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14773_  (.A(\reg_module/gprf[991] ),
    .B(net765),
    .Y(\reg_module/_07439_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14774_  (.A(\reg_module/_07438_ ),
    .B(\reg_module/_04998_ ),
    .C(\reg_module/_07439_ ),
    .Y(\reg_module/_07440_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14775_  (.A(\reg_module/_07437_ ),
    .B(\reg_module/_07440_ ),
    .Y(\reg_module/_07441_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14776_  (.A(\reg_module/_07441_ ),
    .B(\reg_module/_05092_ ),
    .Y(\reg_module/_07442_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14777_  (.A(\reg_module/_07434_ ),
    .B(\reg_module/_07442_ ),
    .C(\reg_module/_06926_ ),
    .Y(\reg_module/_07443_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14778_  (.A(\reg_module/_07081_ ),
    .B(\reg_module/gprf[703] ),
    .Y(\reg_module/_07444_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14779_  (.A(\reg_module/gprf[671] ),
    .B(net766),
    .Y(\reg_module/_07445_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14780_  (.A(\reg_module/_07444_ ),
    .B(net694),
    .C(\reg_module/_07445_ ),
    .Y(\reg_module/_07446_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14781_  (.A(\reg_module/_05079_ ),
    .B(\reg_module/gprf[767] ),
    .Y(\reg_module/_07447_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14782_  (.A(\reg_module/gprf[735] ),
    .B(net766),
    .Y(\reg_module/_07448_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14783_  (.A(\reg_module/_07447_ ),
    .B(\reg_module/_05023_ ),
    .C(\reg_module/_07448_ ),
    .Y(\reg_module/_07449_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14784_  (.A(\reg_module/_07446_ ),
    .B(\reg_module/_07449_ ),
    .Y(\reg_module/_07450_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14785_  (.A(\reg_module/_07450_ ),
    .B(\reg_module/_05304_ ),
    .Y(\reg_module/_07451_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14786_  (.A(\reg_module/_05020_ ),
    .B(\reg_module/gprf[575] ),
    .Y(\reg_module/_07452_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14787_  (.A(\reg_module/gprf[543] ),
    .B(net766),
    .Y(\reg_module/_07453_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14788_  (.A(\reg_module/_07452_ ),
    .B(net694),
    .C(\reg_module/_07453_ ),
    .Y(\reg_module/_07454_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14789_  (.A(\reg_module/_05114_ ),
    .B(\reg_module/gprf[639] ),
    .Y(\reg_module/_07455_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14790_  (.A(\reg_module/gprf[607] ),
    .B(net774),
    .Y(\reg_module/_07456_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14791_  (.A(\reg_module/_07455_ ),
    .B(\reg_module/_05116_ ),
    .C(\reg_module/_07456_ ),
    .Y(\reg_module/_07457_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14792_  (.A(\reg_module/_07454_ ),
    .B(\reg_module/_07457_ ),
    .Y(\reg_module/_07458_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14793_  (.A(\reg_module/_07458_ ),
    .B(net659),
    .Y(\reg_module/_07459_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14794_  (.A(\reg_module/_07451_ ),
    .B(\reg_module/_07459_ ),
    .C(net640),
    .Y(\reg_module/_07460_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14795_  (.A(\reg_module/_07443_ ),
    .B(\reg_module/_07460_ ),
    .Y(\reg_module/_07461_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14796_  (.A(\reg_module/_07461_ ),
    .B(\reg_module/_05124_ ),
    .Y(\reg_module/_07462_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14797_  (.A(\reg_module/_05030_ ),
    .B(\reg_module/gprf[319] ),
    .Y(\reg_module/_07463_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14798_  (.A(\reg_module/gprf[287] ),
    .B(net754),
    .Y(\reg_module/_07464_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14799_  (.A(\reg_module/_07463_ ),
    .B(net689),
    .C(\reg_module/_07464_ ),
    .Y(\reg_module/_07465_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14800_  (.A(\reg_module/_05035_ ),
    .B(\reg_module/gprf[383] ),
    .Y(\reg_module/_07466_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14801_  (.A(\reg_module/gprf[351] ),
    .B(net764),
    .Y(\reg_module/_07467_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14802_  (.A(\reg_module/_07466_ ),
    .B(\reg_module/_05038_ ),
    .C(\reg_module/_07467_ ),
    .Y(\reg_module/_07468_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14803_  (.A(\reg_module/_07465_ ),
    .B(\reg_module/_07468_ ),
    .Y(\reg_module/_07469_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14804_  (.A(\reg_module/_07469_ ),
    .B(net656),
    .Y(\reg_module/_07470_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14805_  (.A(\reg_module/_05044_ ),
    .B(\reg_module/gprf[447] ),
    .Y(\reg_module/_07471_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14806_  (.A(\reg_module/gprf[415] ),
    .B(net754),
    .Y(\reg_module/_07472_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14807_  (.A(\reg_module/_07471_ ),
    .B(net689),
    .C(\reg_module/_07472_ ),
    .Y(\reg_module/_07473_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14808_  (.A(\reg_module/_05049_ ),
    .B(\reg_module/gprf[511] ),
    .Y(\reg_module/_07474_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14809_  (.A(\reg_module/gprf[479] ),
    .B(net754),
    .Y(\reg_module/_07475_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14810_  (.A(\reg_module/_07474_ ),
    .B(\reg_module/_07113_ ),
    .C(\reg_module/_07475_ ),
    .Y(\reg_module/_07476_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14811_  (.A(\reg_module/_07473_ ),
    .B(\reg_module/_07476_ ),
    .Y(\reg_module/_07477_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14812_  (.A(\reg_module/_07477_ ),
    .B(\reg_module/_05057_ ),
    .Y(\reg_module/_07478_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14813_  (.A(\reg_module/_07470_ ),
    .B(\reg_module/_07478_ ),
    .C(\reg_module/_05060_ ),
    .Y(\reg_module/_07479_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14814_  (.A(\reg_module/_05035_ ),
    .B(\reg_module/gprf[63] ),
    .Y(\reg_module/_07480_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14815_  (.A(\reg_module/gprf[31] ),
    .B(net755),
    .Y(\reg_module/_07481_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14816_  (.A(\reg_module/_07480_ ),
    .B(net689),
    .C(\reg_module/_07481_ ),
    .Y(\reg_module/_07482_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14817_  (.A(\reg_module/_05109_ ),
    .B(\reg_module/gprf[127] ),
    .Y(\reg_module/_07483_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14818_  (.A(\reg_module/gprf[95] ),
    .B(net754),
    .Y(\reg_module/_07484_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14819_  (.A(\reg_module/_07483_ ),
    .B(\reg_module/_05087_ ),
    .C(\reg_module/_07484_ ),
    .Y(\reg_module/_07485_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14820_  (.A(\reg_module/_07482_ ),
    .B(\reg_module/_07485_ ),
    .Y(\reg_module/_07486_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14821_  (.A(\reg_module/_07486_ ),
    .B(net656),
    .Y(\reg_module/_07487_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14822_  (.A(\reg_module/_05084_ ),
    .B(\reg_module/gprf[191] ),
    .Y(\reg_module/_07488_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14823_  (.A(\reg_module/gprf[159] ),
    .B(net755),
    .Y(\reg_module/_07489_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14824_  (.A(\reg_module/_07488_ ),
    .B(net689),
    .C(\reg_module/_07489_ ),
    .Y(\reg_module/_07490_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14825_  (.A(\reg_module/_05282_ ),
    .B(\reg_module/gprf[255] ),
    .Y(\reg_module/_07491_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14826_  (.A(\reg_module/gprf[223] ),
    .B(net755),
    .Y(\reg_module/_07492_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14827_  (.A(\reg_module/_07491_ ),
    .B(\reg_module/_05290_ ),
    .C(\reg_module/_07492_ ),
    .Y(\reg_module/_07493_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14828_  (.A(\reg_module/_07490_ ),
    .B(\reg_module/_07493_ ),
    .Y(\reg_module/_07494_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14829_  (.A(\reg_module/_07494_ ),
    .B(\reg_module/_05010_ ),
    .Y(\reg_module/_07495_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14830_  (.A(\reg_module/_07487_ ),
    .B(\reg_module/_07495_ ),
    .C(net642),
    .Y(\reg_module/_07496_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14831_  (.A(\reg_module/_07479_ ),
    .B(\reg_module/_07496_ ),
    .Y(\reg_module/_07497_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14832_  (.A(\reg_module/_07497_ ),
    .B(net632),
    .Y(\reg_module/_07498_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_14833_  (.A(\reg_module/_07462_ ),
    .B(\reg_module/_07498_ ),
    .Y(\wRs1Data[31] ));
 sky130_fd_sc_hd__nand3_4 \reg_module/_14834_  (.A(net994),
    .B(net995),
    .C(net978),
    .Y(\reg_module/_07499_ ));
 sky130_fd_sc_hd__inv_4 \reg_module/_14835_  (.A(\reg_module/_07499_ ),
    .Y(\reg_module/_07500_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14836_  (.A(net962),
    .B(net964),
    .Y(\reg_module/_07501_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14837_  (.A(\reg_module/_07501_ ),
    .Y(\reg_module/_07502_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14838_  (.A(\reg_module/_07500_ ),
    .B(\reg_module/_07502_ ),
    .Y(\reg_module/_07503_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_14839_  (.A(net994),
    .B(net995),
    .Y(\reg_module/_07504_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_14840_  (.A(net962),
    .B(net978),
    .Y(\reg_module/_07505_ ));
 sky130_fd_sc_hd__inv_4 \reg_module/_14841_  (.A(net963),
    .Y(\reg_module/_07506_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_14842_  (.A(\reg_module/_07504_ ),
    .B(\reg_module/_07505_ ),
    .C(\reg_module/_07506_ ),
    .Y(\reg_module/_07507_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14843_  (.A(\reg_module/_07507_ ),
    .B(rRegWrEn2),
    .Y(\reg_module/_07508_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_14844_  (.A(\reg_module/_07503_ ),
    .B(\reg_module/_07508_ ),
    .Y(\reg_module/_07509_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_14845_  (.A(\reg_module/_07509_ ),
    .X(\reg_module/_07510_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14846_  (.A(\reg_module/_07510_ ),
    .X(\reg_module/_07511_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14847_  (.A(\reg_module/_07509_ ),
    .X(\reg_module/_07512_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14848_  (.A(net318),
    .Y(\reg_module/_07513_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14849_  (.A(\reg_module/_07513_ ),
    .X(\reg_module/_07514_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14850_  (.A(\reg_module/_07512_ ),
    .B(\reg_module/_07514_ ),
    .Y(\reg_module/_07515_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14851_  (.A1(net2017),
    .A2(\reg_module/_07511_ ),
    .B1(net1032),
    .C1(\reg_module/_07515_ ),
    .X(\reg_module/_00000_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14852_  (.A(net317),
    .Y(\reg_module/_07516_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_14853_  (.A(\reg_module/_07516_ ),
    .X(\reg_module/_07517_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14854_  (.A(\reg_module/_07512_ ),
    .B(\reg_module/_07517_ ),
    .Y(\reg_module/_07518_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14855_  (.A1(net2009),
    .A2(\reg_module/_07511_ ),
    .B1(net1032),
    .C1(\reg_module/_07518_ ),
    .X(\reg_module/_00001_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14856_  (.A(net316),
    .Y(\reg_module/_07519_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_14857_  (.A(\reg_module/_07519_ ),
    .X(\reg_module/_07520_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14858_  (.A(\reg_module/_07512_ ),
    .B(\reg_module/_07520_ ),
    .Y(\reg_module/_07521_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14859_  (.A1(net2000),
    .A2(\reg_module/_07511_ ),
    .B1(net1036),
    .C1(\reg_module/_07521_ ),
    .X(\reg_module/_00002_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14860_  (.A(net315),
    .Y(\reg_module/_07522_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14861_  (.A(\reg_module/_07522_ ),
    .X(\reg_module/_07523_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14862_  (.A(\reg_module/_07512_ ),
    .B(\reg_module/_07523_ ),
    .Y(\reg_module/_07524_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14863_  (.A1(net2013),
    .A2(\reg_module/_07511_ ),
    .B1(net1035),
    .C1(\reg_module/_07524_ ),
    .X(\reg_module/_00003_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_14864_  (.A(\reg_module/_07509_ ),
    .X(\reg_module/_07525_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14865_  (.A(\reg_module/_07525_ ),
    .X(\reg_module/_07526_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14866_  (.A(\wRegWrData[4] ),
    .Y(\reg_module/_07527_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14867_  (.A(\reg_module/_07527_ ),
    .X(\reg_module/_07528_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14868_  (.A(\reg_module/_07526_ ),
    .B(\reg_module/_07528_ ),
    .Y(\reg_module/_07529_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14869_  (.A1(net1910),
    .A2(\reg_module/_07511_ ),
    .B1(net1051),
    .C1(\reg_module/_07529_ ),
    .X(\reg_module/_00004_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14870_  (.A(net314),
    .Y(\reg_module/_07530_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14871_  (.A(\reg_module/_07530_ ),
    .X(\reg_module/_07531_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14872_  (.A(\reg_module/_07526_ ),
    .B(\reg_module/_07531_ ),
    .Y(\reg_module/_07532_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14873_  (.A1(net1909),
    .A2(\reg_module/_07511_ ),
    .B1(net1051),
    .C1(\reg_module/_07532_ ),
    .X(\reg_module/_00005_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_14874_  (.A(\reg_module/_07510_ ),
    .X(\reg_module/_07533_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14875_  (.A(\wRegWrData[6] ),
    .Y(\reg_module/_07534_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14876_  (.A(\reg_module/_07534_ ),
    .X(\reg_module/_07535_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14877_  (.A(\reg_module/_07526_ ),
    .B(\reg_module/_07535_ ),
    .Y(\reg_module/_07536_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14878_  (.A1(net1723),
    .A2(\reg_module/_07533_ ),
    .B1(net1054),
    .C1(\reg_module/_07536_ ),
    .X(\reg_module/_00006_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14879_  (.A(net313),
    .Y(\reg_module/_07537_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14880_  (.A(\reg_module/_07537_ ),
    .X(\reg_module/_07538_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14881_  (.A(\reg_module/_07526_ ),
    .B(\reg_module/_07538_ ),
    .Y(\reg_module/_07539_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14882_  (.A1(net1807),
    .A2(\reg_module/_07533_ ),
    .B1(net1054),
    .C1(\reg_module/_07539_ ),
    .X(\reg_module/_00007_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14883_  (.A(\wRegWrData[8] ),
    .Y(\reg_module/_07540_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14884_  (.A(\reg_module/_07540_ ),
    .X(\reg_module/_07541_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14885_  (.A(\reg_module/_07526_ ),
    .B(\reg_module/_07541_ ),
    .Y(\reg_module/_07542_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14886_  (.A1(net1831),
    .A2(\reg_module/_07533_ ),
    .B1(net1054),
    .C1(\reg_module/_07542_ ),
    .X(\reg_module/_00008_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14887_  (.A(net312),
    .Y(\reg_module/_07543_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14888_  (.A(\reg_module/_07543_ ),
    .X(\reg_module/_07544_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14889_  (.A(\reg_module/_07526_ ),
    .B(\reg_module/_07544_ ),
    .Y(\reg_module/_07545_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14890_  (.A1(net1946),
    .A2(\reg_module/_07533_ ),
    .B1(net1054),
    .C1(\reg_module/_07545_ ),
    .X(\reg_module/_00009_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_14891_  (.A(\reg_module/_07525_ ),
    .X(\reg_module/_07546_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14892_  (.A(net311),
    .Y(\reg_module/_07547_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14893_  (.A(\reg_module/_07547_ ),
    .X(\reg_module/_07548_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14894_  (.A(\reg_module/_07546_ ),
    .B(\reg_module/_07548_ ),
    .Y(\reg_module/_07549_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14895_  (.A1(net1961),
    .A2(\reg_module/_07533_ ),
    .B1(net1054),
    .C1(\reg_module/_07549_ ),
    .X(\reg_module/_00010_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14896_  (.A(net310),
    .Y(\reg_module/_07550_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14897_  (.A(\reg_module/_07550_ ),
    .X(\reg_module/_07551_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14898_  (.A(\reg_module/_07546_ ),
    .B(\reg_module/_07551_ ),
    .Y(\reg_module/_07552_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14899_  (.A1(net1950),
    .A2(\reg_module/_07533_ ),
    .B1(net1055),
    .C1(\reg_module/_07552_ ),
    .X(\reg_module/_00011_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_14900_  (.A(\reg_module/_07525_ ),
    .X(\reg_module/_07553_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14901_  (.A(\wRegWrData[12] ),
    .Y(\reg_module/_07554_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14902_  (.A(\reg_module/_07554_ ),
    .X(\reg_module/_07555_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14903_  (.A(\reg_module/_07546_ ),
    .B(\reg_module/_07555_ ),
    .Y(\reg_module/_07556_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14904_  (.A1(net1888),
    .A2(\reg_module/_07553_ ),
    .B1(net1065),
    .C1(\reg_module/_07556_ ),
    .X(\reg_module/_00012_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14905_  (.A(net309),
    .Y(\reg_module/_07557_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14906_  (.A(\reg_module/_07557_ ),
    .X(\reg_module/_07558_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14907_  (.A(\reg_module/_07546_ ),
    .B(\reg_module/_07558_ ),
    .Y(\reg_module/_07559_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14908_  (.A1(net1810),
    .A2(\reg_module/_07553_ ),
    .B1(net1065),
    .C1(\reg_module/_07559_ ),
    .X(\reg_module/_00013_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14909_  (.A(net308),
    .Y(\reg_module/_07560_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14910_  (.A(\reg_module/_07560_ ),
    .X(\reg_module/_07561_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14911_  (.A(\reg_module/_07546_ ),
    .B(\reg_module/_07561_ ),
    .Y(\reg_module/_07562_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14912_  (.A1(net1796),
    .A2(\reg_module/_07553_ ),
    .B1(net1065),
    .C1(\reg_module/_07562_ ),
    .X(\reg_module/_00014_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14913_  (.A(net306),
    .Y(\reg_module/_07563_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14914_  (.A(\reg_module/_07563_ ),
    .X(\reg_module/_07564_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14915_  (.A(\reg_module/_07546_ ),
    .B(\reg_module/_07564_ ),
    .Y(\reg_module/_07565_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14916_  (.A1(net1775),
    .A2(\reg_module/_07553_ ),
    .B1(net1065),
    .C1(\reg_module/_07565_ ),
    .X(\reg_module/_00015_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14917_  (.A(\reg_module/_07525_ ),
    .X(\reg_module/_07566_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14918_  (.A(\wRegWrData[16] ),
    .Y(\reg_module/_07567_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_14919_  (.A(\reg_module/_07567_ ),
    .X(\reg_module/_07568_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14920_  (.A(\reg_module/_07566_ ),
    .B(\reg_module/_07568_ ),
    .Y(\reg_module/_07569_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14921_  (.A1(net1926),
    .A2(\reg_module/_07553_ ),
    .B1(net1065),
    .C1(\reg_module/_07569_ ),
    .X(\reg_module/_00016_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14922_  (.A(net305),
    .Y(\reg_module/_07570_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_14923_  (.A(\reg_module/_07570_ ),
    .X(\reg_module/_07571_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14924_  (.A(\reg_module/_07566_ ),
    .B(\reg_module/_07571_ ),
    .Y(\reg_module/_07572_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14925_  (.A1(net2027),
    .A2(\reg_module/_07553_ ),
    .B1(net1067),
    .C1(\reg_module/_07572_ ),
    .X(\reg_module/_00017_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14926_  (.A(\reg_module/_07525_ ),
    .X(\reg_module/_07573_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14927_  (.A(net304),
    .Y(\reg_module/_07574_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14928_  (.A(\reg_module/_07574_ ),
    .X(\reg_module/_07575_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14929_  (.A(\reg_module/_07566_ ),
    .B(\reg_module/_07575_ ),
    .Y(\reg_module/_07576_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14930_  (.A1(net1947),
    .A2(\reg_module/_07573_ ),
    .B1(net1060),
    .C1(\reg_module/_07576_ ),
    .X(\reg_module/_00018_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14931_  (.A(net303),
    .Y(\reg_module/_07577_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_14932_  (.A(\reg_module/_07577_ ),
    .X(\reg_module/_07578_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14933_  (.A(\reg_module/_07566_ ),
    .B(\reg_module/_07578_ ),
    .Y(\reg_module/_07579_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14934_  (.A1(net1977),
    .A2(\reg_module/_07573_ ),
    .B1(net1058),
    .C1(\reg_module/_07579_ ),
    .X(\reg_module/_00019_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14935_  (.A(net302),
    .Y(\reg_module/_07580_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14936_  (.A(\reg_module/_07580_ ),
    .X(\reg_module/_07581_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14937_  (.A(\reg_module/_07566_ ),
    .B(\reg_module/_07581_ ),
    .Y(\reg_module/_07582_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14938_  (.A1(net1859),
    .A2(\reg_module/_07573_ ),
    .B1(net1058),
    .C1(\reg_module/_07582_ ),
    .X(\reg_module/_00020_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14939_  (.A(net301),
    .Y(\reg_module/_07583_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14940_  (.A(\reg_module/_07583_ ),
    .X(\reg_module/_07584_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14941_  (.A(\reg_module/_07566_ ),
    .B(\reg_module/_07584_ ),
    .Y(\reg_module/_07585_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14942_  (.A1(net1965),
    .A2(\reg_module/_07573_ ),
    .B1(net1062),
    .C1(\reg_module/_07585_ ),
    .X(\reg_module/_00021_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14943_  (.A(\reg_module/_07509_ ),
    .X(\reg_module/_07586_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14944_  (.A(net300),
    .Y(\reg_module/_07587_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14945_  (.A(\reg_module/_07587_ ),
    .X(\reg_module/_07588_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14946_  (.A(\reg_module/_07586_ ),
    .B(\reg_module/_07588_ ),
    .Y(\reg_module/_07589_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14947_  (.A1(net1948),
    .A2(\reg_module/_07573_ ),
    .B1(net1024),
    .C1(\reg_module/_07589_ ),
    .X(\reg_module/_00022_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14948_  (.A(net299),
    .Y(\reg_module/_07590_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_14949_  (.A(\reg_module/_07590_ ),
    .X(\reg_module/_07591_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14950_  (.A(\reg_module/_07586_ ),
    .B(\reg_module/_07591_ ),
    .Y(\reg_module/_07592_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14951_  (.A1(net1852),
    .A2(\reg_module/_07573_ ),
    .B1(net1024),
    .C1(\reg_module/_07592_ ),
    .X(\reg_module/_00023_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14952_  (.A(\reg_module/_07525_ ),
    .X(\reg_module/_07593_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14953_  (.A(net298),
    .Y(\reg_module/_07594_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14954_  (.A(\reg_module/_07594_ ),
    .X(\reg_module/_07595_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14955_  (.A(\reg_module/_07586_ ),
    .B(\reg_module/_07595_ ),
    .Y(\reg_module/_07596_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14956_  (.A1(net1713),
    .A2(\reg_module/_07593_ ),
    .B1(net1006),
    .C1(\reg_module/_07596_ ),
    .X(\reg_module/_00024_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14957_  (.A(net296),
    .Y(\reg_module/_07597_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14958_  (.A(\reg_module/_07597_ ),
    .X(\reg_module/_07598_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14959_  (.A(\reg_module/_07586_ ),
    .B(\reg_module/_07598_ ),
    .Y(\reg_module/_07599_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14960_  (.A1(net1787),
    .A2(\reg_module/_07593_ ),
    .B1(net1007),
    .C1(\reg_module/_07599_ ),
    .X(\reg_module/_00025_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14961_  (.A(net294),
    .Y(\reg_module/_07600_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14962_  (.A(\reg_module/_07600_ ),
    .X(\reg_module/_07601_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14963_  (.A(\reg_module/_07586_ ),
    .B(\reg_module/_07601_ ),
    .Y(\reg_module/_07602_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14964_  (.A1(net1799),
    .A2(\reg_module/_07593_ ),
    .B1(net1006),
    .C1(\reg_module/_07602_ ),
    .X(\reg_module/_00026_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14965_  (.A(net293),
    .Y(\reg_module/_07603_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14966_  (.A(\reg_module/_07603_ ),
    .X(\reg_module/_07604_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14967_  (.A(\reg_module/_07586_ ),
    .B(\reg_module/_07604_ ),
    .Y(\reg_module/_07605_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14968_  (.A1(net1850),
    .A2(\reg_module/_07593_ ),
    .B1(net1004),
    .C1(\reg_module/_07605_ ),
    .X(\reg_module/_00027_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14969_  (.A(net292),
    .Y(\reg_module/_07606_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14970_  (.A(\reg_module/_07606_ ),
    .X(\reg_module/_07607_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14971_  (.A(\reg_module/_07510_ ),
    .B(\reg_module/_07607_ ),
    .Y(\reg_module/_07608_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14972_  (.A1(net1726),
    .A2(\reg_module/_07593_ ),
    .B1(net1011),
    .C1(\reg_module/_07608_ ),
    .X(\reg_module/_00028_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14973_  (.A(net290),
    .Y(\reg_module/_07609_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14974_  (.A(\reg_module/_07609_ ),
    .X(\reg_module/_07610_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14975_  (.A(\reg_module/_07510_ ),
    .B(\reg_module/_07610_ ),
    .Y(\reg_module/_07611_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14976_  (.A1(net1768),
    .A2(\reg_module/_07593_ ),
    .B1(net1011),
    .C1(\reg_module/_07611_ ),
    .X(\reg_module/_00029_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14977_  (.A(net289),
    .Y(\reg_module/_07612_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_14978_  (.A(\reg_module/_07612_ ),
    .X(\reg_module/_07613_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14979_  (.A(\reg_module/_07510_ ),
    .B(\reg_module/_07613_ ),
    .Y(\reg_module/_07614_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14980_  (.A1(net1828),
    .A2(\reg_module/_07512_ ),
    .B1(net1010),
    .C1(\reg_module/_07614_ ),
    .X(\reg_module/_00030_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14981_  (.A(net287),
    .Y(\reg_module/_07615_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14982_  (.A(\reg_module/_07615_ ),
    .X(\reg_module/_07616_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14983_  (.A(\reg_module/_07510_ ),
    .B(\reg_module/_07616_ ),
    .Y(\reg_module/_07617_ ));
 sky130_fd_sc_hd__o211a_1 \reg_module/_14984_  (.A1(net1887),
    .A2(\reg_module/_07512_ ),
    .B1(net1010),
    .C1(\reg_module/_07617_ ),
    .X(\reg_module/_00031_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_14985_  (.A(\reg_module/_07501_ ),
    .B(\reg_module/_07499_ ),
    .Y(\reg_module/_07618_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_14986_  (.A(\reg_module/_07618_ ),
    .B(\reg_module/_07508_ ),
    .Y(\reg_module/_07619_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_14987_  (.A(\reg_module/_07619_ ),
    .X(\reg_module/_07620_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_14988_  (.A(\reg_module/_07500_ ),
    .B(net964),
    .Y(\reg_module/_07621_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14989_  (.A(net962),
    .Y(\reg_module/_07622_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14990_  (.A(\reg_module/_07621_ ),
    .B(\reg_module/_07622_ ),
    .Y(\reg_module/_07623_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_14991_  (.A(\reg_module/_07623_ ),
    .X(\reg_module/_07624_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_14992_  (.A(\reg_module/_07506_ ),
    .X(\reg_module/_07625_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_14993_  (.A(\reg_module/_07625_ ),
    .X(\reg_module/_07626_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_14994_  (.A(net995),
    .Y(\reg_module/_07627_ ));
 sky130_fd_sc_hd__and2_1 \reg_module/_14995_  (.A(\reg_module/_07627_ ),
    .B(net994),
    .X(\reg_module/_07628_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_14996_  (.A(\reg_module/_07628_ ),
    .B(net978),
    .Y(\reg_module/_07629_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_14997_  (.A(\reg_module/_07626_ ),
    .B(\reg_module/_07629_ ),
    .Y(\reg_module/_07630_ ));
 sky130_fd_sc_hd__nand3_2 \reg_module/_14998_  (.A(\reg_module/_07620_ ),
    .B(\reg_module/_07624_ ),
    .C(\reg_module/_07630_ ),
    .Y(\reg_module/_07631_ ));
 sky130_fd_sc_hd__buf_8 \reg_module/_14999_  (.A(\reg_module/_07631_ ),
    .X(\reg_module/_07632_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15000_  (.A(\reg_module/_07632_ ),
    .X(\reg_module/_07633_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15001_  (.A(\reg_module/_07633_ ),
    .B(net1997),
    .Y(\reg_module/_07634_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_15002_  (.A(\reg_module/_07506_ ),
    .B(\reg_module/_07499_ ),
    .Y(\reg_module/_07635_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15003_  (.A(net962),
    .B(\reg_module/_07635_ ),
    .Y(\reg_module/_07636_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15004_  (.A(\reg_module/_07503_ ),
    .B(\reg_module/_07507_ ),
    .C(rRegWrEn2),
    .Y(\reg_module/_07637_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15005_  (.A(\reg_module/_07636_ ),
    .B(\reg_module/_07637_ ),
    .Y(\reg_module/_07638_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_15006_  (.A(\reg_module/_07638_ ),
    .X(\reg_module/_07639_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_15007_  (.A(\reg_module/_07639_ ),
    .X(\reg_module/_07640_ ));
 sky130_fd_sc_hd__buf_8 \reg_module/_15008_  (.A(\reg_module/_07640_ ),
    .X(\reg_module/_07641_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_15009_  (.A(\reg_module/_07641_ ),
    .X(\reg_module/_07642_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15010_  (.A(\reg_module/_07499_ ),
    .B(\reg_module/_07506_ ),
    .Y(\reg_module/_07643_ ));
 sky130_fd_sc_hd__nand2_2 \reg_module/_15011_  (.A(\reg_module/_07621_ ),
    .B(\reg_module/_07643_ ),
    .Y(\reg_module/_07644_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_15012_  (.A(\reg_module/_07644_ ),
    .X(\reg_module/_07645_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15013_  (.A(\reg_module/_07645_ ),
    .X(\reg_module/_07646_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15014_  (.A(\reg_module/_07629_ ),
    .Y(\reg_module/_07647_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_15015_  (.A(\reg_module/_07647_ ),
    .X(\reg_module/_07648_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15016_  (.A(\reg_module/_07648_ ),
    .X(\reg_module/_07649_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15017_  (.A(\reg_module/_07649_ ),
    .B(net319),
    .Y(\reg_module/_07650_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15018_  (.A(\reg_module/_07646_ ),
    .B(\reg_module/_07650_ ),
    .Y(\reg_module/_07651_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15019_  (.A(\reg_module/_07642_ ),
    .B(\reg_module/_07651_ ),
    .Y(\reg_module/_07652_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15020_  (.A(net1038),
    .Y(\reg_module/_07653_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_15021_  (.A(\reg_module/_07653_ ),
    .X(\reg_module/_07654_ ));
 sky130_fd_sc_hd__buf_8 \reg_module/_15022_  (.A(\reg_module/_07654_ ),
    .X(\reg_module/_07655_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15023_  (.A(\reg_module/_07655_ ),
    .X(\reg_module/_07656_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15024_  (.A1(\reg_module/_07634_ ),
    .A2(\reg_module/_07652_ ),
    .B1(\reg_module/_07656_ ),
    .Y(\reg_module/_00032_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15025_  (.A(\reg_module/_07633_ ),
    .B(net1267),
    .Y(\reg_module/_07657_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15026_  (.A(\reg_module/_07649_ ),
    .B(net317),
    .Y(\reg_module/_07658_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15027_  (.A(\reg_module/_07646_ ),
    .B(\reg_module/_07658_ ),
    .Y(\reg_module/_07659_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15028_  (.A(\reg_module/_07642_ ),
    .B(\reg_module/_07659_ ),
    .Y(\reg_module/_07660_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15029_  (.A1(\reg_module/_07657_ ),
    .A2(\reg_module/_07660_ ),
    .B1(\reg_module/_07656_ ),
    .Y(\reg_module/_00033_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15030_  (.A(\reg_module/_07633_ ),
    .B(net1318),
    .Y(\reg_module/_07661_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_15031_  (.A(\reg_module/_07644_ ),
    .X(\reg_module/_07662_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15032_  (.A(\reg_module/_07662_ ),
    .X(\reg_module/_07663_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15033_  (.A(\reg_module/_07649_ ),
    .B(\wRegWrData[2] ),
    .Y(\reg_module/_07664_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15034_  (.A(\reg_module/_07663_ ),
    .B(\reg_module/_07664_ ),
    .Y(\reg_module/_07665_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15035_  (.A(\reg_module/_07642_ ),
    .B(\reg_module/_07665_ ),
    .Y(\reg_module/_07666_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15036_  (.A1(\reg_module/_07661_ ),
    .A2(\reg_module/_07666_ ),
    .B1(\reg_module/_07656_ ),
    .Y(\reg_module/_00034_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15037_  (.A(\reg_module/_07633_ ),
    .B(net1392),
    .Y(\reg_module/_07667_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15038_  (.A(\reg_module/_07649_ ),
    .B(net315),
    .Y(\reg_module/_07668_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15039_  (.A(\reg_module/_07663_ ),
    .B(\reg_module/_07668_ ),
    .Y(\reg_module/_07669_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15040_  (.A(\reg_module/_07642_ ),
    .B(\reg_module/_07669_ ),
    .Y(\reg_module/_07670_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15041_  (.A1(\reg_module/_07667_ ),
    .A2(\reg_module/_07670_ ),
    .B1(\reg_module/_07656_ ),
    .Y(\reg_module/_00035_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15042_  (.A(\reg_module/_07633_ ),
    .B(net1565),
    .Y(\reg_module/_07671_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15043_  (.A(\reg_module/_07649_ ),
    .B(\wRegWrData[4] ),
    .Y(\reg_module/_07672_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15044_  (.A(\reg_module/_07663_ ),
    .B(\reg_module/_07672_ ),
    .Y(\reg_module/_07673_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15045_  (.A(\reg_module/_07642_ ),
    .B(\reg_module/_07673_ ),
    .Y(\reg_module/_07674_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15046_  (.A1(\reg_module/_07671_ ),
    .A2(\reg_module/_07674_ ),
    .B1(\reg_module/_07656_ ),
    .Y(\reg_module/_00036_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15047_  (.A(\reg_module/_07633_ ),
    .B(net1606),
    .Y(\reg_module/_07675_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15048_  (.A(\reg_module/_07649_ ),
    .B(net314),
    .Y(\reg_module/_07676_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15049_  (.A(\reg_module/_07663_ ),
    .B(\reg_module/_07676_ ),
    .Y(\reg_module/_07677_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15050_  (.A(\reg_module/_07642_ ),
    .B(\reg_module/_07677_ ),
    .Y(\reg_module/_07678_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15051_  (.A1(\reg_module/_07675_ ),
    .A2(\reg_module/_07678_ ),
    .B1(\reg_module/_07656_ ),
    .Y(\reg_module/_00037_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15052_  (.A(\reg_module/_07632_ ),
    .X(\reg_module/_07679_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15053_  (.A(\reg_module/_07679_ ),
    .B(net1602),
    .Y(\reg_module/_07680_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15054_  (.A(\reg_module/_07641_ ),
    .X(\reg_module/_07681_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15055_  (.A(\reg_module/_07648_ ),
    .X(\reg_module/_07682_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15056_  (.A(\reg_module/_07682_ ),
    .B(\wRegWrData[6] ),
    .Y(\reg_module/_07683_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15057_  (.A(\reg_module/_07663_ ),
    .B(\reg_module/_07683_ ),
    .Y(\reg_module/_07684_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15058_  (.A(\reg_module/_07681_ ),
    .B(\reg_module/_07684_ ),
    .Y(\reg_module/_07685_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15059_  (.A(\reg_module/_07655_ ),
    .X(\reg_module/_07686_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15060_  (.A1(\reg_module/_07680_ ),
    .A2(\reg_module/_07685_ ),
    .B1(\reg_module/_07686_ ),
    .Y(\reg_module/_00038_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15061_  (.A(\reg_module/_07679_ ),
    .B(net1483),
    .Y(\reg_module/_07687_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15062_  (.A(\reg_module/_07682_ ),
    .B(net313),
    .Y(\reg_module/_07688_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15063_  (.A(\reg_module/_07663_ ),
    .B(\reg_module/_07688_ ),
    .Y(\reg_module/_07689_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15064_  (.A(\reg_module/_07681_ ),
    .B(\reg_module/_07689_ ),
    .Y(\reg_module/_07690_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15065_  (.A1(\reg_module/_07687_ ),
    .A2(\reg_module/_07690_ ),
    .B1(\reg_module/_07686_ ),
    .Y(\reg_module/_00039_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15066_  (.A(\reg_module/_07679_ ),
    .B(net1370),
    .Y(\reg_module/_07691_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15067_  (.A(\reg_module/_07662_ ),
    .X(\reg_module/_07692_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15068_  (.A(\reg_module/_07682_ ),
    .B(\wRegWrData[8] ),
    .Y(\reg_module/_07693_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15069_  (.A(\reg_module/_07692_ ),
    .B(\reg_module/_07693_ ),
    .Y(\reg_module/_07694_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15070_  (.A(\reg_module/_07681_ ),
    .B(\reg_module/_07694_ ),
    .Y(\reg_module/_07695_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15071_  (.A1(\reg_module/_07691_ ),
    .A2(\reg_module/_07695_ ),
    .B1(\reg_module/_07686_ ),
    .Y(\reg_module/_00040_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15072_  (.A(\reg_module/_07679_ ),
    .B(net1343),
    .Y(\reg_module/_07696_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15073_  (.A(\reg_module/_07682_ ),
    .B(net312),
    .Y(\reg_module/_07697_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15074_  (.A(\reg_module/_07692_ ),
    .B(\reg_module/_07697_ ),
    .Y(\reg_module/_07698_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15075_  (.A(\reg_module/_07681_ ),
    .B(\reg_module/_07698_ ),
    .Y(\reg_module/_07699_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15076_  (.A1(\reg_module/_07696_ ),
    .A2(\reg_module/_07699_ ),
    .B1(\reg_module/_07686_ ),
    .Y(\reg_module/_00041_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15077_  (.A(\reg_module/_07679_ ),
    .B(net1355),
    .Y(\reg_module/_07700_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15078_  (.A(\reg_module/_07682_ ),
    .B(net311),
    .Y(\reg_module/_07701_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15079_  (.A(\reg_module/_07692_ ),
    .B(\reg_module/_07701_ ),
    .Y(\reg_module/_07702_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15080_  (.A(\reg_module/_07681_ ),
    .B(\reg_module/_07702_ ),
    .Y(\reg_module/_07703_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15081_  (.A1(\reg_module/_07700_ ),
    .A2(\reg_module/_07703_ ),
    .B1(\reg_module/_07686_ ),
    .Y(\reg_module/_00042_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15082_  (.A(\reg_module/_07679_ ),
    .B(net1288),
    .Y(\reg_module/_07704_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15083_  (.A(\reg_module/_07682_ ),
    .B(\wRegWrData[11] ),
    .Y(\reg_module/_07705_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15084_  (.A(\reg_module/_07692_ ),
    .B(\reg_module/_07705_ ),
    .Y(\reg_module/_07706_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15085_  (.A(\reg_module/_07681_ ),
    .B(\reg_module/_07706_ ),
    .Y(\reg_module/_07707_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15086_  (.A1(\reg_module/_07704_ ),
    .A2(\reg_module/_07707_ ),
    .B1(\reg_module/_07686_ ),
    .Y(\reg_module/_00043_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15087_  (.A(\reg_module/_07632_ ),
    .X(\reg_module/_07708_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15088_  (.A(\reg_module/_07708_ ),
    .B(net1962),
    .Y(\reg_module/_07709_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15089_  (.A(\reg_module/_07641_ ),
    .X(\reg_module/_07710_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15090_  (.A(\reg_module/_07648_ ),
    .X(\reg_module/_07711_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15091_  (.A(\reg_module/_07711_ ),
    .B(\wRegWrData[12] ),
    .Y(\reg_module/_07712_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15092_  (.A(\reg_module/_07692_ ),
    .B(\reg_module/_07712_ ),
    .Y(\reg_module/_07713_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15093_  (.A(\reg_module/_07710_ ),
    .B(\reg_module/_07713_ ),
    .Y(\reg_module/_07714_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15094_  (.A(\reg_module/_07655_ ),
    .X(\reg_module/_07715_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15095_  (.A1(\reg_module/_07709_ ),
    .A2(\reg_module/_07714_ ),
    .B1(\reg_module/_07715_ ),
    .Y(\reg_module/_00044_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15096_  (.A(\reg_module/_07708_ ),
    .B(net1676),
    .Y(\reg_module/_07716_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15097_  (.A(\reg_module/_07711_ ),
    .B(net309),
    .Y(\reg_module/_07717_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15098_  (.A(\reg_module/_07692_ ),
    .B(\reg_module/_07717_ ),
    .Y(\reg_module/_07718_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15099_  (.A(\reg_module/_07710_ ),
    .B(\reg_module/_07718_ ),
    .Y(\reg_module/_07719_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15100_  (.A1(\reg_module/_07716_ ),
    .A2(\reg_module/_07719_ ),
    .B1(\reg_module/_07715_ ),
    .Y(\reg_module/_00045_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15101_  (.A(\reg_module/_07708_ ),
    .B(net1735),
    .Y(\reg_module/_07720_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15102_  (.A(\reg_module/_07662_ ),
    .X(\reg_module/_07721_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15103_  (.A(\reg_module/_07711_ ),
    .B(\wRegWrData[14] ),
    .Y(\reg_module/_07722_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15104_  (.A(\reg_module/_07721_ ),
    .B(\reg_module/_07722_ ),
    .Y(\reg_module/_07723_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15105_  (.A(\reg_module/_07710_ ),
    .B(\reg_module/_07723_ ),
    .Y(\reg_module/_07724_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15106_  (.A1(\reg_module/_07720_ ),
    .A2(\reg_module/_07724_ ),
    .B1(\reg_module/_07715_ ),
    .Y(\reg_module/_00046_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15107_  (.A(\reg_module/_07708_ ),
    .B(net1817),
    .Y(\reg_module/_07725_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15108_  (.A(\reg_module/_07711_ ),
    .B(net307),
    .Y(\reg_module/_07726_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15109_  (.A(\reg_module/_07721_ ),
    .B(\reg_module/_07726_ ),
    .Y(\reg_module/_07727_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15110_  (.A(\reg_module/_07710_ ),
    .B(\reg_module/_07727_ ),
    .Y(\reg_module/_07728_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15111_  (.A1(\reg_module/_07725_ ),
    .A2(\reg_module/_07728_ ),
    .B1(\reg_module/_07715_ ),
    .Y(\reg_module/_00047_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15112_  (.A(\reg_module/_07708_ ),
    .B(net1617),
    .Y(\reg_module/_07729_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15113_  (.A(\reg_module/_07711_ ),
    .B(\wRegWrData[16] ),
    .Y(\reg_module/_07730_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15114_  (.A(\reg_module/_07721_ ),
    .B(\reg_module/_07730_ ),
    .Y(\reg_module/_07731_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15115_  (.A(\reg_module/_07710_ ),
    .B(\reg_module/_07731_ ),
    .Y(\reg_module/_07732_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15116_  (.A1(\reg_module/_07729_ ),
    .A2(\reg_module/_07732_ ),
    .B1(\reg_module/_07715_ ),
    .Y(\reg_module/_00048_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15117_  (.A(\reg_module/_07708_ ),
    .B(net1569),
    .Y(\reg_module/_07733_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15118_  (.A(\reg_module/_07711_ ),
    .B(net305),
    .Y(\reg_module/_07734_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15119_  (.A(\reg_module/_07721_ ),
    .B(\reg_module/_07734_ ),
    .Y(\reg_module/_07735_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15120_  (.A(\reg_module/_07710_ ),
    .B(\reg_module/_07735_ ),
    .Y(\reg_module/_07736_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15121_  (.A1(\reg_module/_07733_ ),
    .A2(\reg_module/_07736_ ),
    .B1(\reg_module/_07715_ ),
    .Y(\reg_module/_00049_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15122_  (.A(\reg_module/_07632_ ),
    .X(\reg_module/_07737_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15123_  (.A(\reg_module/_07737_ ),
    .B(net2094),
    .Y(\reg_module/_07738_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15124_  (.A(\reg_module/_07641_ ),
    .X(\reg_module/_07739_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15125_  (.A(\reg_module/_07648_ ),
    .X(\reg_module/_07740_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15126_  (.A(\reg_module/_07740_ ),
    .B(net304),
    .Y(\reg_module/_07741_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15127_  (.A(\reg_module/_07721_ ),
    .B(\reg_module/_07741_ ),
    .Y(\reg_module/_07742_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15128_  (.A(\reg_module/_07739_ ),
    .B(\reg_module/_07742_ ),
    .Y(\reg_module/_07743_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15129_  (.A(\reg_module/_07655_ ),
    .X(\reg_module/_07744_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15130_  (.A1(\reg_module/_07738_ ),
    .A2(\reg_module/_07743_ ),
    .B1(\reg_module/_07744_ ),
    .Y(\reg_module/_00050_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15131_  (.A(\reg_module/_07737_ ),
    .B(net2016),
    .Y(\reg_module/_07745_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15132_  (.A(\reg_module/_07740_ ),
    .B(\wRegWrData[19] ),
    .Y(\reg_module/_07746_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15133_  (.A(\reg_module/_07721_ ),
    .B(\reg_module/_07746_ ),
    .Y(\reg_module/_07747_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15134_  (.A(\reg_module/_07739_ ),
    .B(\reg_module/_07747_ ),
    .Y(\reg_module/_07748_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15135_  (.A1(\reg_module/_07745_ ),
    .A2(\reg_module/_07748_ ),
    .B1(\reg_module/_07744_ ),
    .Y(\reg_module/_00051_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15136_  (.A(\reg_module/_07737_ ),
    .B(net1933),
    .Y(\reg_module/_07749_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15137_  (.A(\reg_module/_07662_ ),
    .X(\reg_module/_07750_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15138_  (.A(\reg_module/_07740_ ),
    .B(\wRegWrData[20] ),
    .Y(\reg_module/_07751_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15139_  (.A(\reg_module/_07750_ ),
    .B(\reg_module/_07751_ ),
    .Y(\reg_module/_07752_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15140_  (.A(\reg_module/_07739_ ),
    .B(\reg_module/_07752_ ),
    .Y(\reg_module/_07753_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15141_  (.A1(\reg_module/_07749_ ),
    .A2(\reg_module/_07753_ ),
    .B1(\reg_module/_07744_ ),
    .Y(\reg_module/_00052_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15142_  (.A(\reg_module/_07737_ ),
    .B(net2088),
    .Y(\reg_module/_07754_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15143_  (.A(\reg_module/_07740_ ),
    .B(\wRegWrData[21] ),
    .Y(\reg_module/_07755_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15144_  (.A(\reg_module/_07750_ ),
    .B(\reg_module/_07755_ ),
    .Y(\reg_module/_07756_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15145_  (.A(\reg_module/_07739_ ),
    .B(\reg_module/_07756_ ),
    .Y(\reg_module/_07757_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15146_  (.A1(\reg_module/_07754_ ),
    .A2(\reg_module/_07757_ ),
    .B1(\reg_module/_07744_ ),
    .Y(\reg_module/_00053_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15147_  (.A(\reg_module/_07737_ ),
    .B(net2020),
    .Y(\reg_module/_07758_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15148_  (.A(\reg_module/_07740_ ),
    .B(\wRegWrData[22] ),
    .Y(\reg_module/_07759_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15149_  (.A(\reg_module/_07750_ ),
    .B(\reg_module/_07759_ ),
    .Y(\reg_module/_07760_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15150_  (.A(\reg_module/_07739_ ),
    .B(\reg_module/_07760_ ),
    .Y(\reg_module/_07761_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15151_  (.A1(\reg_module/_07758_ ),
    .A2(\reg_module/_07761_ ),
    .B1(\reg_module/_07744_ ),
    .Y(\reg_module/_00054_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15152_  (.A(\reg_module/_07737_ ),
    .B(net2130),
    .Y(\reg_module/_07762_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15153_  (.A(\reg_module/_07740_ ),
    .B(\wRegWrData[23] ),
    .Y(\reg_module/_07763_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15154_  (.A(\reg_module/_07750_ ),
    .B(\reg_module/_07763_ ),
    .Y(\reg_module/_07764_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15155_  (.A(\reg_module/_07739_ ),
    .B(\reg_module/_07764_ ),
    .Y(\reg_module/_07765_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15156_  (.A1(\reg_module/_07762_ ),
    .A2(\reg_module/_07765_ ),
    .B1(\reg_module/_07744_ ),
    .Y(\reg_module/_00055_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15157_  (.A(\reg_module/_07631_ ),
    .X(\reg_module/_07766_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15158_  (.A(\reg_module/_07766_ ),
    .B(net1766),
    .Y(\reg_module/_07767_ ));
 sky130_fd_sc_hd__buf_8 \reg_module/_15159_  (.A(\reg_module/_07640_ ),
    .X(\reg_module/_07768_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15160_  (.A(\reg_module/_07768_ ),
    .X(\reg_module/_07769_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15161_  (.A(\reg_module/_07647_ ),
    .X(\reg_module/_07770_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15162_  (.A(\reg_module/_07770_ ),
    .B(net298),
    .Y(\reg_module/_07771_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15163_  (.A(\reg_module/_07750_ ),
    .B(\reg_module/_07771_ ),
    .Y(\reg_module/_07772_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15164_  (.A(\reg_module/_07769_ ),
    .B(\reg_module/_07772_ ),
    .Y(\reg_module/_07773_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_15165_  (.A(\reg_module/_07654_ ),
    .X(\reg_module/_07774_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15166_  (.A(\reg_module/_07774_ ),
    .X(\reg_module/_07775_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15167_  (.A1(\reg_module/_07767_ ),
    .A2(\reg_module/_07773_ ),
    .B1(\reg_module/_07775_ ),
    .Y(\reg_module/_00056_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15168_  (.A(\reg_module/_07766_ ),
    .B(net1521),
    .Y(\reg_module/_07776_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15169_  (.A(\reg_module/_07770_ ),
    .B(net296),
    .Y(\reg_module/_07777_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15170_  (.A(\reg_module/_07750_ ),
    .B(\reg_module/_07777_ ),
    .Y(\reg_module/_07778_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15171_  (.A(\reg_module/_07769_ ),
    .B(\reg_module/_07778_ ),
    .Y(\reg_module/_07779_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15172_  (.A1(\reg_module/_07776_ ),
    .A2(\reg_module/_07779_ ),
    .B1(\reg_module/_07775_ ),
    .Y(\reg_module/_00057_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15173_  (.A(\reg_module/_07766_ ),
    .B(net1397),
    .Y(\reg_module/_07780_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_15174_  (.A(\reg_module/_07644_ ),
    .X(\reg_module/_07781_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15175_  (.A(\reg_module/_07781_ ),
    .X(\reg_module/_07782_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15176_  (.A(\reg_module/_07770_ ),
    .B(net294),
    .Y(\reg_module/_07783_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15177_  (.A(\reg_module/_07782_ ),
    .B(\reg_module/_07783_ ),
    .Y(\reg_module/_07784_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15178_  (.A(\reg_module/_07769_ ),
    .B(\reg_module/_07784_ ),
    .Y(\reg_module/_07785_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15179_  (.A1(\reg_module/_07780_ ),
    .A2(\reg_module/_07785_ ),
    .B1(\reg_module/_07775_ ),
    .Y(\reg_module/_00058_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15180_  (.A(\reg_module/_07766_ ),
    .B(net1459),
    .Y(\reg_module/_07786_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15181_  (.A(\reg_module/_07770_ ),
    .B(\wRegWrData[27] ),
    .Y(\reg_module/_07787_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15182_  (.A(\reg_module/_07782_ ),
    .B(\reg_module/_07787_ ),
    .Y(\reg_module/_07788_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15183_  (.A(\reg_module/_07769_ ),
    .B(\reg_module/_07788_ ),
    .Y(\reg_module/_07789_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15184_  (.A1(\reg_module/_07786_ ),
    .A2(\reg_module/_07789_ ),
    .B1(\reg_module/_07775_ ),
    .Y(\reg_module/_00059_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15185_  (.A(\reg_module/_07766_ ),
    .B(net1680),
    .Y(\reg_module/_07790_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15186_  (.A(\reg_module/_07770_ ),
    .B(net292),
    .Y(\reg_module/_07791_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15187_  (.A(\reg_module/_07782_ ),
    .B(\reg_module/_07791_ ),
    .Y(\reg_module/_07792_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15188_  (.A(\reg_module/_07769_ ),
    .B(\reg_module/_07792_ ),
    .Y(\reg_module/_07793_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15189_  (.A1(\reg_module/_07790_ ),
    .A2(\reg_module/_07793_ ),
    .B1(\reg_module/_07775_ ),
    .Y(\reg_module/_00060_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15190_  (.A(\reg_module/_07766_ ),
    .B(net1855),
    .Y(\reg_module/_07794_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15191_  (.A(\reg_module/_07770_ ),
    .B(net290),
    .Y(\reg_module/_07795_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15192_  (.A(\reg_module/_07782_ ),
    .B(\reg_module/_07795_ ),
    .Y(\reg_module/_07796_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15193_  (.A(\reg_module/_07769_ ),
    .B(\reg_module/_07796_ ),
    .Y(\reg_module/_07797_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15194_  (.A1(\reg_module/_07794_ ),
    .A2(\reg_module/_07797_ ),
    .B1(\reg_module/_07775_ ),
    .Y(\reg_module/_00061_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15195_  (.A(\reg_module/_07632_ ),
    .B(net1994),
    .Y(\reg_module/_07798_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_15196_  (.A(\reg_module/_07768_ ),
    .X(\reg_module/_07799_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15197_  (.A(\reg_module/_07648_ ),
    .B(net289),
    .Y(\reg_module/_07800_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15198_  (.A(\reg_module/_07782_ ),
    .B(\reg_module/_07800_ ),
    .Y(\reg_module/_07801_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15199_  (.A(\reg_module/_07799_ ),
    .B(\reg_module/_07801_ ),
    .Y(\reg_module/_07802_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15200_  (.A(\reg_module/_07774_ ),
    .X(\reg_module/_07803_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15201_  (.A1(\reg_module/_07798_ ),
    .A2(\reg_module/_07802_ ),
    .B1(\reg_module/_07803_ ),
    .Y(\reg_module/_00062_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15202_  (.A(\reg_module/_07632_ ),
    .B(net1653),
    .Y(\reg_module/_07804_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15203_  (.A(\reg_module/_07648_ ),
    .B(net287),
    .Y(\reg_module/_07805_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15204_  (.A(\reg_module/_07782_ ),
    .B(\reg_module/_07805_ ),
    .Y(\reg_module/_07806_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15205_  (.A(\reg_module/_07799_ ),
    .B(\reg_module/_07806_ ),
    .Y(\reg_module/_07807_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15206_  (.A1(\reg_module/_07804_ ),
    .A2(\reg_module/_07807_ ),
    .B1(\reg_module/_07803_ ),
    .Y(\reg_module/_00063_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15207_  (.A(net994),
    .B(\reg_module/_07627_ ),
    .Y(\reg_module/_07808_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15208_  (.A(\reg_module/_07808_ ),
    .B(net978),
    .Y(\reg_module/_07809_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15209_  (.A(\reg_module/_07626_ ),
    .B(\reg_module/_07809_ ),
    .Y(\reg_module/_07810_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15210_  (.A(\reg_module/_07620_ ),
    .B(\reg_module/_07624_ ),
    .C(\reg_module/_07810_ ),
    .Y(\reg_module/_07811_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_15211_  (.A(\reg_module/_07811_ ),
    .X(\reg_module/_07812_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_15212_  (.A(\reg_module/_07812_ ),
    .X(\reg_module/_07813_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15213_  (.A(\reg_module/_07813_ ),
    .B(net1341),
    .Y(\reg_module/_07814_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15214_  (.A(\reg_module/_07781_ ),
    .X(\reg_module/_07815_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15215_  (.A(net978),
    .Y(\reg_module/_07816_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15216_  (.A(\reg_module/_07816_ ),
    .X(\reg_module/_07817_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15217_  (.A(\reg_module/_07817_ ),
    .X(\reg_module/_07818_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_15218_  (.A(\reg_module/_07808_ ),
    .X(\reg_module/_07819_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15219_  (.A(\reg_module/_07819_ ),
    .X(\reg_module/_07820_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15220_  (.A(\reg_module/_07820_ ),
    .B(net318),
    .Y(\reg_module/_07821_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15221_  (.A(\reg_module/_07818_ ),
    .B(\reg_module/_07821_ ),
    .X(\reg_module/_07822_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15222_  (.A(\reg_module/_07815_ ),
    .B(\reg_module/_07822_ ),
    .Y(\reg_module/_07823_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15223_  (.A(\reg_module/_07799_ ),
    .B(\reg_module/_07823_ ),
    .Y(\reg_module/_07824_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15224_  (.A1(\reg_module/_07814_ ),
    .A2(\reg_module/_07824_ ),
    .B1(\reg_module/_07803_ ),
    .Y(\reg_module/_00064_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15225_  (.A(\reg_module/_07813_ ),
    .B(net2029),
    .Y(\reg_module/_07825_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15226_  (.A(\reg_module/_07820_ ),
    .B(net317),
    .Y(\reg_module/_07826_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15227_  (.A(\reg_module/_07818_ ),
    .B(\reg_module/_07826_ ),
    .X(\reg_module/_07827_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15228_  (.A(\reg_module/_07815_ ),
    .B(\reg_module/_07827_ ),
    .Y(\reg_module/_07828_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15229_  (.A(\reg_module/_07799_ ),
    .B(\reg_module/_07828_ ),
    .Y(\reg_module/_07829_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15230_  (.A1(\reg_module/_07825_ ),
    .A2(\reg_module/_07829_ ),
    .B1(\reg_module/_07803_ ),
    .Y(\reg_module/_00065_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15231_  (.A(\reg_module/_07813_ ),
    .B(net1633),
    .Y(\reg_module/_07830_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15232_  (.A(\reg_module/_07820_ ),
    .B(net316),
    .Y(\reg_module/_07831_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15233_  (.A(\reg_module/_07818_ ),
    .B(\reg_module/_07831_ ),
    .X(\reg_module/_07832_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15234_  (.A(\reg_module/_07815_ ),
    .B(\reg_module/_07832_ ),
    .Y(\reg_module/_07833_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15235_  (.A(\reg_module/_07799_ ),
    .B(\reg_module/_07833_ ),
    .Y(\reg_module/_07834_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15236_  (.A1(\reg_module/_07830_ ),
    .A2(\reg_module/_07834_ ),
    .B1(\reg_module/_07803_ ),
    .Y(\reg_module/_00066_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15237_  (.A(\reg_module/_07813_ ),
    .B(net1919),
    .Y(\reg_module/_07835_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15238_  (.A(\reg_module/_07820_ ),
    .B(net315),
    .Y(\reg_module/_07836_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15239_  (.A(\reg_module/_07818_ ),
    .B(\reg_module/_07836_ ),
    .X(\reg_module/_07837_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15240_  (.A(\reg_module/_07815_ ),
    .B(\reg_module/_07837_ ),
    .Y(\reg_module/_07838_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15241_  (.A(\reg_module/_07799_ ),
    .B(\reg_module/_07838_ ),
    .Y(\reg_module/_07839_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15242_  (.A1(\reg_module/_07835_ ),
    .A2(\reg_module/_07839_ ),
    .B1(\reg_module/_07803_ ),
    .Y(\reg_module/_00067_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15243_  (.A(\reg_module/_07813_ ),
    .B(net1463),
    .Y(\reg_module/_07840_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_15244_  (.A(\reg_module/_07768_ ),
    .X(\reg_module/_07841_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_15245_  (.A(\reg_module/_07817_ ),
    .X(\reg_module/_07842_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_15246_  (.A(\reg_module/_07842_ ),
    .X(\reg_module/_07843_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15247_  (.A(\reg_module/_07820_ ),
    .B(\wRegWrData[4] ),
    .Y(\reg_module/_07844_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15248_  (.A(\reg_module/_07843_ ),
    .B(\reg_module/_07844_ ),
    .X(\reg_module/_07845_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15249_  (.A(\reg_module/_07815_ ),
    .B(\reg_module/_07845_ ),
    .Y(\reg_module/_07846_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15250_  (.A(\reg_module/_07841_ ),
    .B(\reg_module/_07846_ ),
    .Y(\reg_module/_07847_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15251_  (.A(\reg_module/_07774_ ),
    .X(\reg_module/_07848_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15252_  (.A1(\reg_module/_07840_ ),
    .A2(\reg_module/_07847_ ),
    .B1(\reg_module/_07848_ ),
    .Y(\reg_module/_00068_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15253_  (.A(\reg_module/_07813_ ),
    .B(net1572),
    .Y(\reg_module/_07849_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15254_  (.A(\reg_module/_07820_ ),
    .B(net314),
    .Y(\reg_module/_07850_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15255_  (.A(\reg_module/_07843_ ),
    .B(\reg_module/_07850_ ),
    .X(\reg_module/_07851_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15256_  (.A(\reg_module/_07815_ ),
    .B(\reg_module/_07851_ ),
    .Y(\reg_module/_07852_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15257_  (.A(\reg_module/_07841_ ),
    .B(\reg_module/_07852_ ),
    .Y(\reg_module/_07853_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15258_  (.A1(\reg_module/_07849_ ),
    .A2(\reg_module/_07853_ ),
    .B1(\reg_module/_07848_ ),
    .Y(\reg_module/_00069_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15259_  (.A(\reg_module/_07812_ ),
    .X(\reg_module/_07854_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15260_  (.A(\reg_module/_07854_ ),
    .B(net1486),
    .Y(\reg_module/_07855_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15261_  (.A(\reg_module/_07781_ ),
    .X(\reg_module/_07856_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15262_  (.A(\reg_module/_07819_ ),
    .X(\reg_module/_07857_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15263_  (.A(\reg_module/_07857_ ),
    .B(\wRegWrData[6] ),
    .Y(\reg_module/_07858_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15264_  (.A(\reg_module/_07843_ ),
    .B(\reg_module/_07858_ ),
    .X(\reg_module/_07859_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15265_  (.A(\reg_module/_07856_ ),
    .B(\reg_module/_07859_ ),
    .Y(\reg_module/_07860_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15266_  (.A(\reg_module/_07841_ ),
    .B(\reg_module/_07860_ ),
    .Y(\reg_module/_07861_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15267_  (.A1(\reg_module/_07855_ ),
    .A2(\reg_module/_07861_ ),
    .B1(\reg_module/_07848_ ),
    .Y(\reg_module/_00070_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15268_  (.A(\reg_module/_07854_ ),
    .B(net1434),
    .Y(\reg_module/_07862_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15269_  (.A(\reg_module/_07857_ ),
    .B(net313),
    .Y(\reg_module/_07863_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15270_  (.A(\reg_module/_07843_ ),
    .B(\reg_module/_07863_ ),
    .X(\reg_module/_07864_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15271_  (.A(\reg_module/_07856_ ),
    .B(\reg_module/_07864_ ),
    .Y(\reg_module/_07865_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15272_  (.A(\reg_module/_07841_ ),
    .B(\reg_module/_07865_ ),
    .Y(\reg_module/_07866_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15273_  (.A1(\reg_module/_07862_ ),
    .A2(\reg_module/_07866_ ),
    .B1(\reg_module/_07848_ ),
    .Y(\reg_module/_00071_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15274_  (.A(\reg_module/_07854_ ),
    .B(net1344),
    .Y(\reg_module/_07867_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15275_  (.A(\reg_module/_07857_ ),
    .B(\wRegWrData[8] ),
    .Y(\reg_module/_07868_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15276_  (.A(\reg_module/_07843_ ),
    .B(\reg_module/_07868_ ),
    .X(\reg_module/_07869_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15277_  (.A(\reg_module/_07856_ ),
    .B(\reg_module/_07869_ ),
    .Y(\reg_module/_07870_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15278_  (.A(\reg_module/_07841_ ),
    .B(\reg_module/_07870_ ),
    .Y(\reg_module/_07871_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15279_  (.A1(\reg_module/_07867_ ),
    .A2(\reg_module/_07871_ ),
    .B1(\reg_module/_07848_ ),
    .Y(\reg_module/_00072_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15280_  (.A(\reg_module/_07854_ ),
    .B(net1315),
    .Y(\reg_module/_07872_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15281_  (.A(\reg_module/_07857_ ),
    .B(net312),
    .Y(\reg_module/_07873_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15282_  (.A(\reg_module/_07843_ ),
    .B(\reg_module/_07873_ ),
    .X(\reg_module/_07874_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15283_  (.A(\reg_module/_07856_ ),
    .B(\reg_module/_07874_ ),
    .Y(\reg_module/_07875_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15284_  (.A(\reg_module/_07841_ ),
    .B(\reg_module/_07875_ ),
    .Y(\reg_module/_07876_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15285_  (.A1(\reg_module/_07872_ ),
    .A2(\reg_module/_07876_ ),
    .B1(\reg_module/_07848_ ),
    .Y(\reg_module/_00073_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15286_  (.A(\reg_module/_07854_ ),
    .B(net1575),
    .Y(\reg_module/_07877_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15287_  (.A(\reg_module/_07768_ ),
    .X(\reg_module/_07878_ ));
 sky130_fd_sc_hd__buf_1 \reg_module/_15288_  (.A(\reg_module/_07842_ ),
    .X(\reg_module/_07879_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15289_  (.A(\reg_module/_07857_ ),
    .B(net311),
    .Y(\reg_module/_07880_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15290_  (.A(\reg_module/_07879_ ),
    .B(\reg_module/_07880_ ),
    .X(\reg_module/_07881_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15291_  (.A(\reg_module/_07856_ ),
    .B(\reg_module/_07881_ ),
    .Y(\reg_module/_07882_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15292_  (.A(\reg_module/_07878_ ),
    .B(\reg_module/_07882_ ),
    .Y(\reg_module/_07883_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15293_  (.A(\reg_module/_07774_ ),
    .X(\reg_module/_07884_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15294_  (.A1(\reg_module/_07877_ ),
    .A2(\reg_module/_07883_ ),
    .B1(\reg_module/_07884_ ),
    .Y(\reg_module/_00074_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15295_  (.A(\reg_module/_07854_ ),
    .B(net1596),
    .Y(\reg_module/_07885_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15296_  (.A(\reg_module/_07857_ ),
    .B(net310),
    .Y(\reg_module/_07886_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15297_  (.A(\reg_module/_07879_ ),
    .B(\reg_module/_07886_ ),
    .X(\reg_module/_07887_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15298_  (.A(\reg_module/_07856_ ),
    .B(\reg_module/_07887_ ),
    .Y(\reg_module/_07888_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15299_  (.A(\reg_module/_07878_ ),
    .B(\reg_module/_07888_ ),
    .Y(\reg_module/_07889_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15300_  (.A1(\reg_module/_07885_ ),
    .A2(\reg_module/_07889_ ),
    .B1(\reg_module/_07884_ ),
    .Y(\reg_module/_00075_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15301_  (.A(\reg_module/_07812_ ),
    .X(\reg_module/_07890_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15302_  (.A(\reg_module/_07890_ ),
    .B(net1426),
    .Y(\reg_module/_07891_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_15303_  (.A(\reg_module/_07781_ ),
    .X(\reg_module/_07892_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_15304_  (.A(\reg_module/_07819_ ),
    .X(\reg_module/_07893_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15305_  (.A(\reg_module/_07893_ ),
    .B(\wRegWrData[12] ),
    .Y(\reg_module/_07894_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15306_  (.A(\reg_module/_07879_ ),
    .B(\reg_module/_07894_ ),
    .X(\reg_module/_07895_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15307_  (.A(\reg_module/_07892_ ),
    .B(\reg_module/_07895_ ),
    .Y(\reg_module/_07896_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15308_  (.A(\reg_module/_07878_ ),
    .B(\reg_module/_07896_ ),
    .Y(\reg_module/_07897_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15309_  (.A1(\reg_module/_07891_ ),
    .A2(\reg_module/_07897_ ),
    .B1(\reg_module/_07884_ ),
    .Y(\reg_module/_00076_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15310_  (.A(\reg_module/_07890_ ),
    .B(net1352),
    .Y(\reg_module/_07898_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15311_  (.A(\reg_module/_07893_ ),
    .B(net309),
    .Y(\reg_module/_07899_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15312_  (.A(\reg_module/_07879_ ),
    .B(\reg_module/_07899_ ),
    .X(\reg_module/_07900_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15313_  (.A(\reg_module/_07892_ ),
    .B(\reg_module/_07900_ ),
    .Y(\reg_module/_07901_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15314_  (.A(\reg_module/_07878_ ),
    .B(\reg_module/_07901_ ),
    .Y(\reg_module/_07902_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15315_  (.A1(\reg_module/_07898_ ),
    .A2(\reg_module/_07902_ ),
    .B1(\reg_module/_07884_ ),
    .Y(\reg_module/_00077_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15316_  (.A(\reg_module/_07890_ ),
    .B(net1313),
    .Y(\reg_module/_07903_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15317_  (.A(\reg_module/_07893_ ),
    .B(net308),
    .Y(\reg_module/_07904_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15318_  (.A(\reg_module/_07879_ ),
    .B(\reg_module/_07904_ ),
    .X(\reg_module/_07905_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15319_  (.A(\reg_module/_07892_ ),
    .B(\reg_module/_07905_ ),
    .Y(\reg_module/_07906_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15320_  (.A(\reg_module/_07878_ ),
    .B(\reg_module/_07906_ ),
    .Y(\reg_module/_07907_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15321_  (.A1(\reg_module/_07903_ ),
    .A2(\reg_module/_07907_ ),
    .B1(\reg_module/_07884_ ),
    .Y(\reg_module/_00078_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15322_  (.A(\reg_module/_07890_ ),
    .B(net1504),
    .Y(\reg_module/_07908_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15323_  (.A(\reg_module/_07893_ ),
    .B(net306),
    .Y(\reg_module/_07909_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15324_  (.A(\reg_module/_07879_ ),
    .B(\reg_module/_07909_ ),
    .X(\reg_module/_07910_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15325_  (.A(\reg_module/_07892_ ),
    .B(\reg_module/_07910_ ),
    .Y(\reg_module/_07911_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15326_  (.A(\reg_module/_07878_ ),
    .B(\reg_module/_07911_ ),
    .Y(\reg_module/_07912_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15327_  (.A1(\reg_module/_07908_ ),
    .A2(\reg_module/_07912_ ),
    .B1(\reg_module/_07884_ ),
    .Y(\reg_module/_00079_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15328_  (.A(\reg_module/_07890_ ),
    .B(net1732),
    .Y(\reg_module/_07913_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_15329_  (.A(\reg_module/_07768_ ),
    .X(\reg_module/_07914_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15330_  (.A(\reg_module/_07842_ ),
    .X(\reg_module/_07915_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15331_  (.A(\reg_module/_07893_ ),
    .B(\wRegWrData[16] ),
    .Y(\reg_module/_07916_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15332_  (.A(\reg_module/_07915_ ),
    .B(\reg_module/_07916_ ),
    .X(\reg_module/_07917_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15333_  (.A(\reg_module/_07892_ ),
    .B(\reg_module/_07917_ ),
    .Y(\reg_module/_07918_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15334_  (.A(\reg_module/_07914_ ),
    .B(\reg_module/_07918_ ),
    .Y(\reg_module/_07919_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_15335_  (.A(\reg_module/_07774_ ),
    .X(\reg_module/_07920_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15336_  (.A1(\reg_module/_07913_ ),
    .A2(\reg_module/_07919_ ),
    .B1(\reg_module/_07920_ ),
    .Y(\reg_module/_00080_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15337_  (.A(\reg_module/_07890_ ),
    .B(net1711),
    .Y(\reg_module/_07921_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15338_  (.A(\reg_module/_07893_ ),
    .B(net305),
    .Y(\reg_module/_07922_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15339_  (.A(\reg_module/_07915_ ),
    .B(\reg_module/_07922_ ),
    .X(\reg_module/_07923_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15340_  (.A(\reg_module/_07892_ ),
    .B(\reg_module/_07923_ ),
    .Y(\reg_module/_07924_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15341_  (.A(\reg_module/_07914_ ),
    .B(\reg_module/_07924_ ),
    .Y(\reg_module/_07925_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15342_  (.A1(\reg_module/_07921_ ),
    .A2(\reg_module/_07925_ ),
    .B1(\reg_module/_07920_ ),
    .Y(\reg_module/_00081_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15343_  (.A(\reg_module/_07812_ ),
    .X(\reg_module/_07926_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15344_  (.A(\reg_module/_07926_ ),
    .B(net1800),
    .Y(\reg_module/_07927_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15345_  (.A(\reg_module/_07781_ ),
    .X(\reg_module/_07928_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_15346_  (.A(\reg_module/_07819_ ),
    .X(\reg_module/_07929_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15347_  (.A(\reg_module/_07929_ ),
    .B(net304),
    .Y(\reg_module/_07930_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15348_  (.A(\reg_module/_07915_ ),
    .B(\reg_module/_07930_ ),
    .X(\reg_module/_07931_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15349_  (.A(\reg_module/_07928_ ),
    .B(\reg_module/_07931_ ),
    .Y(\reg_module/_07932_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15350_  (.A(\reg_module/_07914_ ),
    .B(\reg_module/_07932_ ),
    .Y(\reg_module/_07933_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15351_  (.A1(\reg_module/_07927_ ),
    .A2(\reg_module/_07933_ ),
    .B1(\reg_module/_07920_ ),
    .Y(\reg_module/_00082_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15352_  (.A(\reg_module/_07926_ ),
    .B(net1584),
    .Y(\reg_module/_07934_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15353_  (.A(\reg_module/_07929_ ),
    .B(net303),
    .Y(\reg_module/_07935_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15354_  (.A(\reg_module/_07915_ ),
    .B(\reg_module/_07935_ ),
    .X(\reg_module/_07936_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15355_  (.A(\reg_module/_07928_ ),
    .B(\reg_module/_07936_ ),
    .Y(\reg_module/_07937_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15356_  (.A(\reg_module/_07914_ ),
    .B(\reg_module/_07937_ ),
    .Y(\reg_module/_07938_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15357_  (.A1(\reg_module/_07934_ ),
    .A2(\reg_module/_07938_ ),
    .B1(\reg_module/_07920_ ),
    .Y(\reg_module/_00083_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15358_  (.A(\reg_module/_07926_ ),
    .B(net1439),
    .Y(\reg_module/_07939_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15359_  (.A(\reg_module/_07929_ ),
    .B(net302),
    .Y(\reg_module/_07940_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15360_  (.A(\reg_module/_07915_ ),
    .B(\reg_module/_07940_ ),
    .X(\reg_module/_07941_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15361_  (.A(\reg_module/_07928_ ),
    .B(\reg_module/_07941_ ),
    .Y(\reg_module/_07942_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15362_  (.A(\reg_module/_07914_ ),
    .B(\reg_module/_07942_ ),
    .Y(\reg_module/_07943_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15363_  (.A1(\reg_module/_07939_ ),
    .A2(\reg_module/_07943_ ),
    .B1(\reg_module/_07920_ ),
    .Y(\reg_module/_00084_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15364_  (.A(\reg_module/_07926_ ),
    .B(net1626),
    .Y(\reg_module/_07944_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15365_  (.A(\reg_module/_07929_ ),
    .B(net301),
    .Y(\reg_module/_07945_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15366_  (.A(\reg_module/_07915_ ),
    .B(\reg_module/_07945_ ),
    .X(\reg_module/_07946_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15367_  (.A(\reg_module/_07928_ ),
    .B(\reg_module/_07946_ ),
    .Y(\reg_module/_07947_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15368_  (.A(\reg_module/_07914_ ),
    .B(\reg_module/_07947_ ),
    .Y(\reg_module/_07948_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15369_  (.A1(\reg_module/_07944_ ),
    .A2(\reg_module/_07948_ ),
    .B1(\reg_module/_07920_ ),
    .Y(\reg_module/_00085_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15370_  (.A(\reg_module/_07926_ ),
    .B(net1875),
    .Y(\reg_module/_07949_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15371_  (.A(\reg_module/_07768_ ),
    .X(\reg_module/_07950_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_15372_  (.A(\reg_module/_07817_ ),
    .X(\reg_module/_07951_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15373_  (.A(\reg_module/_07929_ ),
    .B(net300),
    .Y(\reg_module/_07952_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15374_  (.A(\reg_module/_07951_ ),
    .B(\reg_module/_07952_ ),
    .X(\reg_module/_07953_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15375_  (.A(\reg_module/_07928_ ),
    .B(\reg_module/_07953_ ),
    .Y(\reg_module/_07954_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15376_  (.A(\reg_module/_07950_ ),
    .B(\reg_module/_07954_ ),
    .Y(\reg_module/_07955_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15377_  (.A(\reg_module/_07774_ ),
    .X(\reg_module/_07956_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15378_  (.A1(\reg_module/_07949_ ),
    .A2(\reg_module/_07955_ ),
    .B1(\reg_module/_07956_ ),
    .Y(\reg_module/_00086_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15379_  (.A(\reg_module/_07926_ ),
    .B(net1679),
    .Y(\reg_module/_07957_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15380_  (.A(\reg_module/_07929_ ),
    .B(net299),
    .Y(\reg_module/_07958_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15381_  (.A(\reg_module/_07951_ ),
    .B(\reg_module/_07958_ ),
    .X(\reg_module/_07959_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15382_  (.A(\reg_module/_07928_ ),
    .B(\reg_module/_07959_ ),
    .Y(\reg_module/_07960_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15383_  (.A(\reg_module/_07950_ ),
    .B(\reg_module/_07960_ ),
    .Y(\reg_module/_07961_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15384_  (.A1(\reg_module/_07957_ ),
    .A2(\reg_module/_07961_ ),
    .B1(\reg_module/_07956_ ),
    .Y(\reg_module/_00087_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15385_  (.A(\reg_module/_07811_ ),
    .X(\reg_module/_07962_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15386_  (.A(\reg_module/_07962_ ),
    .B(net1266),
    .Y(\reg_module/_07963_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15387_  (.A(\reg_module/_07781_ ),
    .X(\reg_module/_07964_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15388_  (.A(\reg_module/_07808_ ),
    .X(\reg_module/_07965_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15389_  (.A(\reg_module/_07965_ ),
    .B(net298),
    .Y(\reg_module/_07966_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15390_  (.A(\reg_module/_07951_ ),
    .B(\reg_module/_07966_ ),
    .X(\reg_module/_07967_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15391_  (.A(\reg_module/_07964_ ),
    .B(\reg_module/_07967_ ),
    .Y(\reg_module/_07968_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15392_  (.A(\reg_module/_07950_ ),
    .B(\reg_module/_07968_ ),
    .Y(\reg_module/_07969_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15393_  (.A1(\reg_module/_07963_ ),
    .A2(\reg_module/_07969_ ),
    .B1(\reg_module/_07956_ ),
    .Y(\reg_module/_00088_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15394_  (.A(\reg_module/_07962_ ),
    .B(net1449),
    .Y(\reg_module/_07970_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15395_  (.A(\reg_module/_07965_ ),
    .B(net296),
    .Y(\reg_module/_07971_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15396_  (.A(\reg_module/_07951_ ),
    .B(\reg_module/_07971_ ),
    .X(\reg_module/_07972_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15397_  (.A(\reg_module/_07964_ ),
    .B(\reg_module/_07972_ ),
    .Y(\reg_module/_07973_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15398_  (.A(\reg_module/_07950_ ),
    .B(\reg_module/_07973_ ),
    .Y(\reg_module/_07974_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15399_  (.A1(\reg_module/_07970_ ),
    .A2(\reg_module/_07974_ ),
    .B1(\reg_module/_07956_ ),
    .Y(\reg_module/_00089_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15400_  (.A(\reg_module/_07962_ ),
    .B(net1560),
    .Y(\reg_module/_07975_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15401_  (.A(\reg_module/_07965_ ),
    .B(net294),
    .Y(\reg_module/_07976_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15402_  (.A(\reg_module/_07951_ ),
    .B(\reg_module/_07976_ ),
    .X(\reg_module/_07977_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15403_  (.A(\reg_module/_07964_ ),
    .B(\reg_module/_07977_ ),
    .Y(\reg_module/_07978_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15404_  (.A(\reg_module/_07950_ ),
    .B(\reg_module/_07978_ ),
    .Y(\reg_module/_07979_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15405_  (.A1(\reg_module/_07975_ ),
    .A2(\reg_module/_07979_ ),
    .B1(\reg_module/_07956_ ),
    .Y(\reg_module/_00090_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15406_  (.A(\reg_module/_07962_ ),
    .B(net1631),
    .Y(\reg_module/_07980_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15407_  (.A(\reg_module/_07965_ ),
    .B(net293),
    .Y(\reg_module/_07981_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15408_  (.A(\reg_module/_07951_ ),
    .B(\reg_module/_07981_ ),
    .X(\reg_module/_07982_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15409_  (.A(\reg_module/_07964_ ),
    .B(\reg_module/_07982_ ),
    .Y(\reg_module/_07983_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15410_  (.A(\reg_module/_07950_ ),
    .B(\reg_module/_07983_ ),
    .Y(\reg_module/_07984_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15411_  (.A1(\reg_module/_07980_ ),
    .A2(\reg_module/_07984_ ),
    .B1(\reg_module/_07956_ ),
    .Y(\reg_module/_00091_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15412_  (.A(\reg_module/_07962_ ),
    .B(net1512),
    .Y(\reg_module/_07985_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_15413_  (.A(\reg_module/_07640_ ),
    .X(\reg_module/_07986_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_15414_  (.A(\reg_module/_07986_ ),
    .X(\reg_module/_07987_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15415_  (.A(\reg_module/_07817_ ),
    .X(\reg_module/_07988_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15416_  (.A(\reg_module/_07965_ ),
    .B(net292),
    .Y(\reg_module/_07989_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15417_  (.A(\reg_module/_07988_ ),
    .B(\reg_module/_07989_ ),
    .X(\reg_module/_07990_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15418_  (.A(\reg_module/_07964_ ),
    .B(\reg_module/_07990_ ),
    .Y(\reg_module/_07991_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15419_  (.A(\reg_module/_07987_ ),
    .B(\reg_module/_07991_ ),
    .Y(\reg_module/_07992_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15420_  (.A(\reg_module/_07653_ ),
    .X(\reg_module/_07993_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_15421_  (.A(\reg_module/_07993_ ),
    .X(\reg_module/_07994_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15422_  (.A(\reg_module/_07994_ ),
    .X(\reg_module/_07995_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15423_  (.A1(\reg_module/_07985_ ),
    .A2(\reg_module/_07992_ ),
    .B1(\reg_module/_07995_ ),
    .Y(\reg_module/_00092_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15424_  (.A(\reg_module/_07962_ ),
    .B(net1357),
    .Y(\reg_module/_07996_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15425_  (.A(\reg_module/_07965_ ),
    .B(net290),
    .Y(\reg_module/_07997_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15426_  (.A(\reg_module/_07988_ ),
    .B(\reg_module/_07997_ ),
    .X(\reg_module/_07998_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15427_  (.A(\reg_module/_07964_ ),
    .B(\reg_module/_07998_ ),
    .Y(\reg_module/_07999_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15428_  (.A(\reg_module/_07987_ ),
    .B(\reg_module/_07999_ ),
    .Y(\reg_module/_08000_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15429_  (.A1(\reg_module/_07996_ ),
    .A2(\reg_module/_08000_ ),
    .B1(\reg_module/_07995_ ),
    .Y(\reg_module/_00093_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15430_  (.A(\reg_module/_07812_ ),
    .B(net1761),
    .Y(\reg_module/_08001_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15431_  (.A(\reg_module/_07645_ ),
    .X(\reg_module/_08002_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15432_  (.A(\reg_module/_07819_ ),
    .B(net289),
    .Y(\reg_module/_08003_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15433_  (.A(\reg_module/_07988_ ),
    .B(\reg_module/_08003_ ),
    .X(\reg_module/_08004_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15434_  (.A(\reg_module/_08002_ ),
    .B(\reg_module/_08004_ ),
    .Y(\reg_module/_08005_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15435_  (.A(\reg_module/_07987_ ),
    .B(\reg_module/_08005_ ),
    .Y(\reg_module/_08006_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15436_  (.A1(\reg_module/_08001_ ),
    .A2(\reg_module/_08006_ ),
    .B1(\reg_module/_07995_ ),
    .Y(\reg_module/_00094_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15437_  (.A(\reg_module/_07812_ ),
    .B(net1383),
    .Y(\reg_module/_08007_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15438_  (.A(\reg_module/_07819_ ),
    .B(net287),
    .Y(\reg_module/_08008_ ));
 sky130_fd_sc_hd__or2_1 \reg_module/_15439_  (.A(\reg_module/_07988_ ),
    .B(\reg_module/_08008_ ),
    .X(\reg_module/_08009_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15440_  (.A(\reg_module/_08002_ ),
    .B(\reg_module/_08009_ ),
    .Y(\reg_module/_08010_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15441_  (.A(\reg_module/_07987_ ),
    .B(\reg_module/_08010_ ),
    .Y(\reg_module/_08011_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15442_  (.A1(\reg_module/_08007_ ),
    .A2(\reg_module/_08011_ ),
    .B1(\reg_module/_07995_ ),
    .Y(\reg_module/_00095_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15443_  (.A(\reg_module/_07504_ ),
    .Y(\reg_module/_08012_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15444_  (.A(\reg_module/_07816_ ),
    .B(\reg_module/_08012_ ),
    .Y(\reg_module/_08013_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15445_  (.A(\reg_module/_08013_ ),
    .B(net965),
    .Y(\reg_module/_08014_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15446_  (.A(\reg_module/_08014_ ),
    .Y(\reg_module/_08015_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15447_  (.A(\reg_module/_07620_ ),
    .B(\reg_module/_07624_ ),
    .C(\reg_module/_08015_ ),
    .Y(\reg_module/_08016_ ));
 sky130_fd_sc_hd__buf_8 \reg_module/_15448_  (.A(\reg_module/_08016_ ),
    .X(\reg_module/_08017_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_15449_  (.A(\reg_module/_08017_ ),
    .X(\reg_module/_08018_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15450_  (.A(\reg_module/_08018_ ),
    .B(net1371),
    .Y(\reg_module/_08019_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_15451_  (.A(\reg_module/_08013_ ),
    .X(\reg_module/_08020_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_15452_  (.A(\reg_module/_08020_ ),
    .X(\reg_module/_08021_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15453_  (.A(\reg_module/_08021_ ),
    .B(net318),
    .Y(\reg_module/_08022_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_15454_  (.A(\reg_module/_07662_ ),
    .X(\reg_module/_08023_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15455_  (.A(\reg_module/_08022_ ),
    .B(\reg_module/_08023_ ),
    .Y(\reg_module/_08024_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15456_  (.A(\reg_module/_07987_ ),
    .B(\reg_module/_08024_ ),
    .Y(\reg_module/_08025_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15457_  (.A1(\reg_module/_08019_ ),
    .A2(\reg_module/_08025_ ),
    .B1(\reg_module/_07995_ ),
    .Y(\reg_module/_00096_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15458_  (.A(\reg_module/_08018_ ),
    .B(net1983),
    .Y(\reg_module/_08026_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15459_  (.A(\reg_module/_08021_ ),
    .B(\wRegWrData[1] ),
    .Y(\reg_module/_08027_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_15460_  (.A(\reg_module/_07644_ ),
    .X(\reg_module/_08028_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_15461_  (.A(\reg_module/_08028_ ),
    .X(\reg_module/_08029_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15462_  (.A(\reg_module/_08027_ ),
    .B(\reg_module/_08029_ ),
    .Y(\reg_module/_08030_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15463_  (.A(\reg_module/_07987_ ),
    .B(\reg_module/_08030_ ),
    .Y(\reg_module/_08031_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15464_  (.A1(\reg_module/_08026_ ),
    .A2(\reg_module/_08031_ ),
    .B1(\reg_module/_07995_ ),
    .Y(\reg_module/_00097_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15465_  (.A(\reg_module/_08018_ ),
    .B(net2140),
    .Y(\reg_module/_08032_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_15466_  (.A(\reg_module/_07986_ ),
    .X(\reg_module/_08033_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15467_  (.A(\reg_module/_08021_ ),
    .B(net316),
    .Y(\reg_module/_08034_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15468_  (.A(\reg_module/_08034_ ),
    .B(\reg_module/_08029_ ),
    .Y(\reg_module/_08035_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15469_  (.A(\reg_module/_08033_ ),
    .B(\reg_module/_08035_ ),
    .Y(\reg_module/_08036_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15470_  (.A(\reg_module/_07994_ ),
    .X(\reg_module/_08037_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15471_  (.A1(\reg_module/_08032_ ),
    .A2(\reg_module/_08036_ ),
    .B1(\reg_module/_08037_ ),
    .Y(\reg_module/_00098_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15472_  (.A(\reg_module/_08018_ ),
    .B(net1991),
    .Y(\reg_module/_08038_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15473_  (.A(\reg_module/_08021_ ),
    .B(net315),
    .Y(\reg_module/_08039_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15474_  (.A(\reg_module/_08039_ ),
    .B(\reg_module/_08029_ ),
    .Y(\reg_module/_08040_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15475_  (.A(\reg_module/_08033_ ),
    .B(\reg_module/_08040_ ),
    .Y(\reg_module/_08041_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15476_  (.A1(\reg_module/_08038_ ),
    .A2(\reg_module/_08041_ ),
    .B1(\reg_module/_08037_ ),
    .Y(\reg_module/_00099_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15477_  (.A(\reg_module/_08018_ ),
    .B(net1433),
    .Y(\reg_module/_08042_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15478_  (.A(\reg_module/_08021_ ),
    .B(\wRegWrData[4] ),
    .Y(\reg_module/_08043_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15479_  (.A(\reg_module/_08043_ ),
    .B(\reg_module/_08029_ ),
    .Y(\reg_module/_08044_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15480_  (.A(\reg_module/_08033_ ),
    .B(\reg_module/_08044_ ),
    .Y(\reg_module/_08045_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15481_  (.A1(\reg_module/_08042_ ),
    .A2(\reg_module/_08045_ ),
    .B1(\reg_module/_08037_ ),
    .Y(\reg_module/_00100_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15482_  (.A(\reg_module/_08018_ ),
    .B(net1456),
    .Y(\reg_module/_08046_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15483_  (.A(\reg_module/_08021_ ),
    .B(\wRegWrData[5] ),
    .Y(\reg_module/_08047_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15484_  (.A(\reg_module/_08047_ ),
    .B(\reg_module/_08023_ ),
    .Y(\reg_module/_08048_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15485_  (.A(\reg_module/_08033_ ),
    .B(\reg_module/_08048_ ),
    .Y(\reg_module/_08049_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15486_  (.A1(\reg_module/_08046_ ),
    .A2(\reg_module/_08049_ ),
    .B1(\reg_module/_08037_ ),
    .Y(\reg_module/_00101_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15487_  (.A(\reg_module/_08017_ ),
    .X(\reg_module/_08050_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15488_  (.A(\reg_module/_08050_ ),
    .B(net1546),
    .Y(\reg_module/_08051_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15489_  (.A(\reg_module/_08020_ ),
    .X(\reg_module/_08052_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15490_  (.A(\reg_module/_08052_ ),
    .B(\wRegWrData[6] ),
    .Y(\reg_module/_08053_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15491_  (.A(\reg_module/_08053_ ),
    .B(\reg_module/_08029_ ),
    .Y(\reg_module/_08054_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15492_  (.A(\reg_module/_08033_ ),
    .B(\reg_module/_08054_ ),
    .Y(\reg_module/_08055_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15493_  (.A1(\reg_module/_08051_ ),
    .A2(\reg_module/_08055_ ),
    .B1(\reg_module/_08037_ ),
    .Y(\reg_module/_00102_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15494_  (.A(\reg_module/_08050_ ),
    .B(net1470),
    .Y(\reg_module/_08056_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15495_  (.A(\reg_module/_08052_ ),
    .B(\wRegWrData[7] ),
    .Y(\reg_module/_08057_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15496_  (.A(\reg_module/_08057_ ),
    .B(\reg_module/_08029_ ),
    .Y(\reg_module/_08058_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15497_  (.A(\reg_module/_08033_ ),
    .B(\reg_module/_08058_ ),
    .Y(\reg_module/_08059_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15498_  (.A1(\reg_module/_08056_ ),
    .A2(\reg_module/_08059_ ),
    .B1(\reg_module/_08037_ ),
    .Y(\reg_module/_00103_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15499_  (.A(\reg_module/_08050_ ),
    .B(net1668),
    .Y(\reg_module/_08060_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15500_  (.A(\reg_module/_07986_ ),
    .X(\reg_module/_08061_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15501_  (.A(\reg_module/_08052_ ),
    .B(\wRegWrData[8] ),
    .Y(\reg_module/_08062_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15502_  (.A(\reg_module/_08028_ ),
    .X(\reg_module/_08063_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15503_  (.A(\reg_module/_08062_ ),
    .B(\reg_module/_08063_ ),
    .Y(\reg_module/_08064_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15504_  (.A(\reg_module/_08061_ ),
    .B(\reg_module/_08064_ ),
    .Y(\reg_module/_08065_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15505_  (.A(\reg_module/_07994_ ),
    .X(\reg_module/_08066_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15506_  (.A1(\reg_module/_08060_ ),
    .A2(\reg_module/_08065_ ),
    .B1(\reg_module/_08066_ ),
    .Y(\reg_module/_00104_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15507_  (.A(\reg_module/_08050_ ),
    .B(net1533),
    .Y(\reg_module/_08067_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15508_  (.A(\reg_module/_08052_ ),
    .B(\wRegWrData[9] ),
    .Y(\reg_module/_08068_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15509_  (.A(\reg_module/_08068_ ),
    .B(\reg_module/_08063_ ),
    .Y(\reg_module/_08069_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15510_  (.A(\reg_module/_08061_ ),
    .B(\reg_module/_08069_ ),
    .Y(\reg_module/_08070_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15511_  (.A1(\reg_module/_08067_ ),
    .A2(\reg_module/_08070_ ),
    .B1(\reg_module/_08066_ ),
    .Y(\reg_module/_00105_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15512_  (.A(\reg_module/_08050_ ),
    .B(net1375),
    .Y(\reg_module/_08071_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15513_  (.A(\reg_module/_08052_ ),
    .B(\wRegWrData[10] ),
    .Y(\reg_module/_08072_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15514_  (.A(\reg_module/_08072_ ),
    .B(\reg_module/_08063_ ),
    .Y(\reg_module/_08073_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15515_  (.A(\reg_module/_08061_ ),
    .B(\reg_module/_08073_ ),
    .Y(\reg_module/_08074_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15516_  (.A1(\reg_module/_08071_ ),
    .A2(\reg_module/_08074_ ),
    .B1(\reg_module/_08066_ ),
    .Y(\reg_module/_00106_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15517_  (.A(\reg_module/_08050_ ),
    .B(net1646),
    .Y(\reg_module/_08075_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15518_  (.A(\reg_module/_08052_ ),
    .B(net310),
    .Y(\reg_module/_08076_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15519_  (.A(\reg_module/_08076_ ),
    .B(\reg_module/_08063_ ),
    .Y(\reg_module/_08077_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15520_  (.A(\reg_module/_08061_ ),
    .B(\reg_module/_08077_ ),
    .Y(\reg_module/_08078_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15521_  (.A1(\reg_module/_08075_ ),
    .A2(\reg_module/_08078_ ),
    .B1(\reg_module/_08066_ ),
    .Y(\reg_module/_00107_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15522_  (.A(\reg_module/_08017_ ),
    .X(\reg_module/_08079_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15523_  (.A(\reg_module/_08079_ ),
    .B(net1362),
    .Y(\reg_module/_08080_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15524_  (.A(\reg_module/_08020_ ),
    .X(\reg_module/_08081_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15525_  (.A(\reg_module/_08081_ ),
    .B(\wRegWrData[12] ),
    .Y(\reg_module/_08082_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15526_  (.A(\reg_module/_08082_ ),
    .B(\reg_module/_08023_ ),
    .Y(\reg_module/_08083_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15527_  (.A(\reg_module/_08061_ ),
    .B(\reg_module/_08083_ ),
    .Y(\reg_module/_08084_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15528_  (.A1(\reg_module/_08080_ ),
    .A2(\reg_module/_08084_ ),
    .B1(\reg_module/_08066_ ),
    .Y(\reg_module/_00108_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15529_  (.A(\reg_module/_08079_ ),
    .B(net1421),
    .Y(\reg_module/_08085_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15530_  (.A(\reg_module/_08081_ ),
    .B(\wRegWrData[13] ),
    .Y(\reg_module/_08086_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15531_  (.A(\reg_module/_08086_ ),
    .B(\reg_module/_08063_ ),
    .Y(\reg_module/_08087_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15532_  (.A(\reg_module/_08061_ ),
    .B(\reg_module/_08087_ ),
    .Y(\reg_module/_08088_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15533_  (.A1(\reg_module/_08085_ ),
    .A2(\reg_module/_08088_ ),
    .B1(\reg_module/_08066_ ),
    .Y(\reg_module/_00109_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15534_  (.A(\reg_module/_08079_ ),
    .B(net1435),
    .Y(\reg_module/_08089_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_15535_  (.A(\reg_module/_07986_ ),
    .X(\reg_module/_08090_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15536_  (.A(\reg_module/_08081_ ),
    .B(net308),
    .Y(\reg_module/_08091_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15537_  (.A(\reg_module/_08091_ ),
    .B(\reg_module/_08063_ ),
    .Y(\reg_module/_08092_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15538_  (.A(\reg_module/_08090_ ),
    .B(\reg_module/_08092_ ),
    .Y(\reg_module/_08093_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15539_  (.A(\reg_module/_07994_ ),
    .X(\reg_module/_08094_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15540_  (.A1(\reg_module/_08089_ ),
    .A2(\reg_module/_08093_ ),
    .B1(\reg_module/_08094_ ),
    .Y(\reg_module/_00110_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15541_  (.A(\reg_module/_08079_ ),
    .B(net1312),
    .Y(\reg_module/_08095_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15542_  (.A(\reg_module/_08081_ ),
    .B(net306),
    .Y(\reg_module/_08096_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_15543_  (.A(\reg_module/_08028_ ),
    .X(\reg_module/_08097_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15544_  (.A(\reg_module/_08096_ ),
    .B(\reg_module/_08097_ ),
    .Y(\reg_module/_08098_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15545_  (.A(\reg_module/_08090_ ),
    .B(\reg_module/_08098_ ),
    .Y(\reg_module/_08099_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15546_  (.A1(\reg_module/_08095_ ),
    .A2(\reg_module/_08099_ ),
    .B1(\reg_module/_08094_ ),
    .Y(\reg_module/_00111_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15547_  (.A(\reg_module/_08079_ ),
    .B(net1651),
    .Y(\reg_module/_08100_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15548_  (.A(\reg_module/_08081_ ),
    .B(\wRegWrData[16] ),
    .Y(\reg_module/_08101_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15549_  (.A(\reg_module/_08101_ ),
    .B(\reg_module/_08097_ ),
    .Y(\reg_module/_08102_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15550_  (.A(\reg_module/_08090_ ),
    .B(\reg_module/_08102_ ),
    .Y(\reg_module/_08103_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15551_  (.A1(\reg_module/_08100_ ),
    .A2(\reg_module/_08103_ ),
    .B1(\reg_module/_08094_ ),
    .Y(\reg_module/_00112_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15552_  (.A(\reg_module/_08079_ ),
    .B(net1405),
    .Y(\reg_module/_08104_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15553_  (.A(\reg_module/_08081_ ),
    .B(\wRegWrData[17] ),
    .Y(\reg_module/_08105_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15554_  (.A(\reg_module/_08105_ ),
    .B(\reg_module/_08097_ ),
    .Y(\reg_module/_08106_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15555_  (.A(\reg_module/_08090_ ),
    .B(\reg_module/_08106_ ),
    .Y(\reg_module/_08107_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15556_  (.A1(\reg_module/_08104_ ),
    .A2(\reg_module/_08107_ ),
    .B1(\reg_module/_08094_ ),
    .Y(\reg_module/_00113_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15557_  (.A(\reg_module/_08017_ ),
    .X(\reg_module/_08108_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15558_  (.A(\reg_module/_08108_ ),
    .B(net1536),
    .Y(\reg_module/_08109_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15559_  (.A(\reg_module/_08020_ ),
    .X(\reg_module/_08110_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15560_  (.A(\reg_module/_08110_ ),
    .B(\wRegWrData[18] ),
    .Y(\reg_module/_08111_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15561_  (.A(\reg_module/_08111_ ),
    .B(\reg_module/_08097_ ),
    .Y(\reg_module/_08112_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15562_  (.A(\reg_module/_08090_ ),
    .B(\reg_module/_08112_ ),
    .Y(\reg_module/_08113_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15563_  (.A1(\reg_module/_08109_ ),
    .A2(\reg_module/_08113_ ),
    .B1(\reg_module/_08094_ ),
    .Y(\reg_module/_00114_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15564_  (.A(\reg_module/_08108_ ),
    .B(net1303),
    .Y(\reg_module/_08114_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15565_  (.A(\reg_module/_08110_ ),
    .B(\wRegWrData[19] ),
    .Y(\reg_module/_08115_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15566_  (.A(\reg_module/_08115_ ),
    .B(\reg_module/_08097_ ),
    .Y(\reg_module/_08116_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15567_  (.A(\reg_module/_08090_ ),
    .B(\reg_module/_08116_ ),
    .Y(\reg_module/_08117_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15568_  (.A1(\reg_module/_08114_ ),
    .A2(\reg_module/_08117_ ),
    .B1(\reg_module/_08094_ ),
    .Y(\reg_module/_00115_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15569_  (.A(\reg_module/_08108_ ),
    .B(net1970),
    .Y(\reg_module/_08118_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_15570_  (.A(\reg_module/_07986_ ),
    .X(\reg_module/_08119_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15571_  (.A(\reg_module/_08110_ ),
    .B(net302),
    .Y(\reg_module/_08120_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15572_  (.A(\reg_module/_08120_ ),
    .B(\reg_module/_08097_ ),
    .Y(\reg_module/_08121_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15573_  (.A(\reg_module/_08119_ ),
    .B(\reg_module/_08121_ ),
    .Y(\reg_module/_08122_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15574_  (.A(\reg_module/_07994_ ),
    .X(\reg_module/_08123_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15575_  (.A1(\reg_module/_08118_ ),
    .A2(\reg_module/_08122_ ),
    .B1(\reg_module/_08123_ ),
    .Y(\reg_module/_00116_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15576_  (.A(\reg_module/_08108_ ),
    .B(net2031),
    .Y(\reg_module/_08124_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15577_  (.A(\reg_module/_08110_ ),
    .B(\wRegWrData[21] ),
    .Y(\reg_module/_08125_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15578_  (.A(\reg_module/_07662_ ),
    .X(\reg_module/_08126_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15579_  (.A(\reg_module/_08125_ ),
    .B(\reg_module/_08126_ ),
    .Y(\reg_module/_08127_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15580_  (.A(\reg_module/_08119_ ),
    .B(\reg_module/_08127_ ),
    .Y(\reg_module/_08128_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15581_  (.A1(\reg_module/_08124_ ),
    .A2(\reg_module/_08128_ ),
    .B1(\reg_module/_08123_ ),
    .Y(\reg_module/_00117_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15582_  (.A(\reg_module/_08108_ ),
    .B(net1641),
    .Y(\reg_module/_08129_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15583_  (.A(\reg_module/_08110_ ),
    .B(net300),
    .Y(\reg_module/_08130_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15584_  (.A(\reg_module/_08130_ ),
    .B(\reg_module/_08126_ ),
    .Y(\reg_module/_08131_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15585_  (.A(\reg_module/_08119_ ),
    .B(\reg_module/_08131_ ),
    .Y(\reg_module/_08132_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15586_  (.A1(\reg_module/_08129_ ),
    .A2(\reg_module/_08132_ ),
    .B1(\reg_module/_08123_ ),
    .Y(\reg_module/_00118_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15587_  (.A(\reg_module/_08108_ ),
    .B(net1539),
    .Y(\reg_module/_08133_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15588_  (.A(\reg_module/_08110_ ),
    .B(net299),
    .Y(\reg_module/_08134_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15589_  (.A(\reg_module/_08134_ ),
    .B(\reg_module/_08126_ ),
    .Y(\reg_module/_08135_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15590_  (.A(\reg_module/_08119_ ),
    .B(\reg_module/_08135_ ),
    .Y(\reg_module/_08136_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15591_  (.A1(\reg_module/_08133_ ),
    .A2(\reg_module/_08136_ ),
    .B1(\reg_module/_08123_ ),
    .Y(\reg_module/_00119_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15592_  (.A(\reg_module/_08016_ ),
    .X(\reg_module/_08137_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15593_  (.A(\reg_module/_08137_ ),
    .B(net1425),
    .Y(\reg_module/_08138_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15594_  (.A(\reg_module/_08013_ ),
    .X(\reg_module/_08139_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15595_  (.A(\reg_module/_08139_ ),
    .B(net298),
    .Y(\reg_module/_08140_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15596_  (.A(\reg_module/_08140_ ),
    .B(\reg_module/_08126_ ),
    .Y(\reg_module/_08141_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15597_  (.A(\reg_module/_08119_ ),
    .B(\reg_module/_08141_ ),
    .Y(\reg_module/_08142_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15598_  (.A1(\reg_module/_08138_ ),
    .A2(\reg_module/_08142_ ),
    .B1(\reg_module/_08123_ ),
    .Y(\reg_module/_00120_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15599_  (.A(\reg_module/_08137_ ),
    .B(net1625),
    .Y(\reg_module/_08143_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15600_  (.A(\reg_module/_08139_ ),
    .B(net296),
    .Y(\reg_module/_08144_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15601_  (.A(\reg_module/_08144_ ),
    .B(\reg_module/_08126_ ),
    .Y(\reg_module/_08145_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15602_  (.A(\reg_module/_08119_ ),
    .B(\reg_module/_08145_ ),
    .Y(\reg_module/_08146_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15603_  (.A1(\reg_module/_08143_ ),
    .A2(\reg_module/_08146_ ),
    .B1(\reg_module/_08123_ ),
    .Y(\reg_module/_00121_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15604_  (.A(\reg_module/_08137_ ),
    .B(net1864),
    .Y(\reg_module/_08147_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15605_  (.A(\reg_module/_07986_ ),
    .X(\reg_module/_08148_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15606_  (.A(\reg_module/_08139_ ),
    .B(net294),
    .Y(\reg_module/_08149_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15607_  (.A(\reg_module/_08149_ ),
    .B(\reg_module/_08126_ ),
    .Y(\reg_module/_08150_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15608_  (.A(\reg_module/_08148_ ),
    .B(\reg_module/_08150_ ),
    .Y(\reg_module/_08151_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15609_  (.A(\reg_module/_07994_ ),
    .X(\reg_module/_08152_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15610_  (.A1(\reg_module/_08147_ ),
    .A2(\reg_module/_08151_ ),
    .B1(\reg_module/_08152_ ),
    .Y(\reg_module/_00122_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15611_  (.A(\reg_module/_08137_ ),
    .B(net1811),
    .Y(\reg_module/_08153_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15612_  (.A(\reg_module/_08139_ ),
    .B(net293),
    .Y(\reg_module/_08154_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15613_  (.A(\reg_module/_08154_ ),
    .B(\reg_module/_07646_ ),
    .Y(\reg_module/_08155_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15614_  (.A(\reg_module/_08148_ ),
    .B(\reg_module/_08155_ ),
    .Y(\reg_module/_08156_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15615_  (.A1(\reg_module/_08153_ ),
    .A2(\reg_module/_08156_ ),
    .B1(\reg_module/_08152_ ),
    .Y(\reg_module/_00123_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15616_  (.A(\reg_module/_08137_ ),
    .B(net1247),
    .Y(\reg_module/_08157_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15617_  (.A(\reg_module/_08139_ ),
    .B(net292),
    .Y(\reg_module/_08158_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15618_  (.A(\reg_module/_08158_ ),
    .B(\reg_module/_08023_ ),
    .Y(\reg_module/_08159_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15619_  (.A(\reg_module/_08148_ ),
    .B(\reg_module/_08159_ ),
    .Y(\reg_module/_08160_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15620_  (.A1(\reg_module/_08157_ ),
    .A2(\reg_module/_08160_ ),
    .B1(\reg_module/_08152_ ),
    .Y(\reg_module/_00124_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15621_  (.A(\reg_module/_08137_ ),
    .B(net1581),
    .Y(\reg_module/_08161_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15622_  (.A(\reg_module/_08139_ ),
    .B(net290),
    .Y(\reg_module/_08162_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15623_  (.A(\reg_module/_08162_ ),
    .B(\reg_module/_07646_ ),
    .Y(\reg_module/_08163_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15624_  (.A(\reg_module/_08148_ ),
    .B(\reg_module/_08163_ ),
    .Y(\reg_module/_08164_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15625_  (.A1(\reg_module/_08161_ ),
    .A2(\reg_module/_08164_ ),
    .B1(\reg_module/_08152_ ),
    .Y(\reg_module/_00125_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15626_  (.A(\reg_module/_08017_ ),
    .B(net1414),
    .Y(\reg_module/_08165_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15627_  (.A(\reg_module/_08020_ ),
    .B(net289),
    .Y(\reg_module/_08166_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15628_  (.A(\reg_module/_08166_ ),
    .B(\reg_module/_07646_ ),
    .Y(\reg_module/_08167_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15629_  (.A(\reg_module/_08148_ ),
    .B(\reg_module/_08167_ ),
    .Y(\reg_module/_08168_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15630_  (.A1(\reg_module/_08165_ ),
    .A2(\reg_module/_08168_ ),
    .B1(\reg_module/_08152_ ),
    .Y(\reg_module/_00126_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15631_  (.A(\reg_module/_08017_ ),
    .B(net1302),
    .Y(\reg_module/_08169_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15632_  (.A(\reg_module/_08020_ ),
    .B(net287),
    .Y(\reg_module/_08170_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15633_  (.A(\reg_module/_08170_ ),
    .B(\reg_module/_07646_ ),
    .Y(\reg_module/_08171_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15634_  (.A(\reg_module/_08148_ ),
    .B(\reg_module/_08171_ ),
    .Y(\reg_module/_08172_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15635_  (.A1(\reg_module/_08169_ ),
    .A2(\reg_module/_08172_ ),
    .B1(\reg_module/_08152_ ),
    .Y(\reg_module/_00127_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15636_  (.A(net994),
    .B(net995),
    .Y(\reg_module/_08173_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15637_  (.A(net979),
    .B(\reg_module/_08173_ ),
    .Y(\reg_module/_08174_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15638_  (.A(\reg_module/_08174_ ),
    .B(net963),
    .Y(\reg_module/_08175_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15639_  (.A(\reg_module/_08175_ ),
    .Y(\reg_module/_08176_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15640_  (.A(\reg_module/_07638_ ),
    .B(\reg_module/_08176_ ),
    .Y(\reg_module/_08177_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_15641_  (.A(\reg_module/_08177_ ),
    .X(\reg_module/_08178_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15642_  (.A(\reg_module/_08178_ ),
    .X(\reg_module/_08179_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15643_  (.A(\reg_module/gprf[128] ),
    .Y(\reg_module/_08180_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15644_  (.A(\reg_module/_08179_ ),
    .B(\reg_module/_08180_ ),
    .Y(\reg_module/_08181_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15645_  (.A(\reg_module/_08181_ ),
    .Y(\reg_module/_08182_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_15646_  (.A(\reg_module/_07639_ ),
    .X(\reg_module/_08183_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_15647_  (.A(\reg_module/_08183_ ),
    .X(\reg_module/_08184_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_15648_  (.A(\reg_module/_08184_ ),
    .X(\reg_module/_08185_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_15649_  (.A(\reg_module/_08176_ ),
    .X(\reg_module/_08186_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15650_  (.A(\reg_module/_08186_ ),
    .X(\reg_module/_08187_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15651_  (.A(\reg_module/_08185_ ),
    .B(\reg_module/_07514_ ),
    .C(\reg_module/_08187_ ),
    .Y(\reg_module/_08188_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15652_  (.A(\reg_module/_08188_ ),
    .B(net1033),
    .Y(\reg_module/_08189_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15653_  (.A(\reg_module/_08182_ ),
    .B(\reg_module/_08189_ ),
    .Y(\reg_module/_00128_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15654_  (.A(net2217),
    .Y(\reg_module/_08190_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15655_  (.A(\reg_module/_08179_ ),
    .B(\reg_module/_08190_ ),
    .Y(\reg_module/_08191_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15656_  (.A(\reg_module/_08191_ ),
    .Y(\reg_module/_08192_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15657_  (.A(\reg_module/_08185_ ),
    .B(\reg_module/_07517_ ),
    .C(\reg_module/_08187_ ),
    .Y(\reg_module/_08193_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15658_  (.A(\reg_module/_08193_ ),
    .B(net1033),
    .Y(\reg_module/_08194_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15659_  (.A(\reg_module/_08192_ ),
    .B(\reg_module/_08194_ ),
    .Y(\reg_module/_00129_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15660_  (.A(\reg_module/gprf[130] ),
    .Y(\reg_module/_08195_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15661_  (.A(\reg_module/_08179_ ),
    .B(\reg_module/_08195_ ),
    .Y(\reg_module/_08196_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15662_  (.A(\reg_module/_08196_ ),
    .Y(\reg_module/_08197_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15663_  (.A(\reg_module/_08185_ ),
    .B(\reg_module/_07520_ ),
    .C(\reg_module/_08187_ ),
    .Y(\reg_module/_08198_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15664_  (.A(\reg_module/_08198_ ),
    .B(net1036),
    .Y(\reg_module/_08199_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15665_  (.A(\reg_module/_08197_ ),
    .B(\reg_module/_08199_ ),
    .Y(\reg_module/_00130_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15666_  (.A(\reg_module/gprf[131] ),
    .Y(\reg_module/_08200_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15667_  (.A(\reg_module/_08179_ ),
    .B(\reg_module/_08200_ ),
    .Y(\reg_module/_08201_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15668_  (.A(\reg_module/_08201_ ),
    .Y(\reg_module/_08202_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15669_  (.A(\reg_module/_08185_ ),
    .B(\reg_module/_07523_ ),
    .C(\reg_module/_08187_ ),
    .Y(\reg_module/_08203_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15670_  (.A(\reg_module/_08203_ ),
    .B(net1035),
    .Y(\reg_module/_08204_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15671_  (.A(\reg_module/_08202_ ),
    .B(\reg_module/_08204_ ),
    .Y(\reg_module/_00131_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15672_  (.A(net2189),
    .Y(\reg_module/_08205_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15673_  (.A(\reg_module/_08179_ ),
    .B(\reg_module/_08205_ ),
    .Y(\reg_module/_08206_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15674_  (.A(\reg_module/_08206_ ),
    .Y(\reg_module/_08207_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15675_  (.A(\reg_module/_08184_ ),
    .X(\reg_module/_08208_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15676_  (.A(\reg_module/_08208_ ),
    .B(\reg_module/_07528_ ),
    .C(\reg_module/_08187_ ),
    .Y(\reg_module/_08209_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15677_  (.A(\reg_module/_08209_ ),
    .B(net1047),
    .Y(\reg_module/_08210_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15678_  (.A(\reg_module/_08207_ ),
    .B(\reg_module/_08210_ ),
    .Y(\reg_module/_00132_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15679_  (.A(net2173),
    .Y(\reg_module/_08211_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15680_  (.A(\reg_module/_08179_ ),
    .B(\reg_module/_08211_ ),
    .Y(\reg_module/_08212_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15681_  (.A(\reg_module/_08212_ ),
    .Y(\reg_module/_08213_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15682_  (.A(\reg_module/_08208_ ),
    .B(\reg_module/_07531_ ),
    .C(\reg_module/_08187_ ),
    .Y(\reg_module/_08214_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15683_  (.A(\reg_module/_08214_ ),
    .B(net1047),
    .Y(\reg_module/_08215_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15684_  (.A(\reg_module/_08213_ ),
    .B(\reg_module/_08215_ ),
    .Y(\reg_module/_00133_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15685_  (.A(\reg_module/_08178_ ),
    .X(\reg_module/_08216_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15686_  (.A(\reg_module/gprf[134] ),
    .Y(\reg_module/_08217_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15687_  (.A(\reg_module/_08216_ ),
    .B(\reg_module/_08217_ ),
    .Y(\reg_module/_08218_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15688_  (.A(\reg_module/_08218_ ),
    .Y(\reg_module/_08219_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_15689_  (.A(\reg_module/_08186_ ),
    .X(\reg_module/_08220_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15690_  (.A(\reg_module/_08208_ ),
    .B(\reg_module/_07535_ ),
    .C(\reg_module/_08220_ ),
    .Y(\reg_module/_08221_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15691_  (.A(\reg_module/_08221_ ),
    .B(net1048),
    .Y(\reg_module/_08222_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15692_  (.A(\reg_module/_08219_ ),
    .B(\reg_module/_08222_ ),
    .Y(\reg_module/_00134_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15693_  (.A(net2214),
    .Y(\reg_module/_08223_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15694_  (.A(\reg_module/_08216_ ),
    .B(\reg_module/_08223_ ),
    .Y(\reg_module/_08224_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15695_  (.A(\reg_module/_08224_ ),
    .Y(\reg_module/_08225_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15696_  (.A(\reg_module/_08208_ ),
    .B(\reg_module/_07538_ ),
    .C(\reg_module/_08220_ ),
    .Y(\reg_module/_08226_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15697_  (.A(\reg_module/_08226_ ),
    .B(net1048),
    .Y(\reg_module/_08227_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15698_  (.A(\reg_module/_08225_ ),
    .B(\reg_module/_08227_ ),
    .Y(\reg_module/_00135_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15699_  (.A(\reg_module/gprf[136] ),
    .Y(\reg_module/_08228_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15700_  (.A(\reg_module/_08216_ ),
    .B(\reg_module/_08228_ ),
    .Y(\reg_module/_08229_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15701_  (.A(\reg_module/_08229_ ),
    .Y(\reg_module/_08230_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15702_  (.A(\reg_module/_08208_ ),
    .B(\reg_module/_07541_ ),
    .C(\reg_module/_08220_ ),
    .Y(\reg_module/_08231_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15703_  (.A(\reg_module/_08231_ ),
    .B(net1048),
    .Y(\reg_module/_08232_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15704_  (.A(\reg_module/_08230_ ),
    .B(\reg_module/_08232_ ),
    .Y(\reg_module/_00136_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15705_  (.A(\reg_module/gprf[137] ),
    .Y(\reg_module/_08233_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15706_  (.A(\reg_module/_08216_ ),
    .B(\reg_module/_08233_ ),
    .Y(\reg_module/_08234_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15707_  (.A(\reg_module/_08234_ ),
    .Y(\reg_module/_08235_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15708_  (.A(\reg_module/_08208_ ),
    .B(\reg_module/_07544_ ),
    .C(\reg_module/_08220_ ),
    .Y(\reg_module/_08236_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15709_  (.A(\reg_module/_08236_ ),
    .B(net1048),
    .Y(\reg_module/_08237_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15710_  (.A(\reg_module/_08235_ ),
    .B(\reg_module/_08237_ ),
    .Y(\reg_module/_00137_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15711_  (.A(net2205),
    .Y(\reg_module/_08238_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15712_  (.A(\reg_module/_08216_ ),
    .B(\reg_module/_08238_ ),
    .Y(\reg_module/_08239_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15713_  (.A(\reg_module/_08239_ ),
    .Y(\reg_module/_08240_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15714_  (.A(\reg_module/_08184_ ),
    .X(\reg_module/_08241_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15715_  (.A(\reg_module/_08241_ ),
    .B(\reg_module/_07548_ ),
    .C(\reg_module/_08220_ ),
    .Y(\reg_module/_08242_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15716_  (.A(\reg_module/_08242_ ),
    .B(net1054),
    .Y(\reg_module/_08243_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15717_  (.A(\reg_module/_08240_ ),
    .B(\reg_module/_08243_ ),
    .Y(\reg_module/_00138_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15718_  (.A(\reg_module/gprf[139] ),
    .Y(\reg_module/_08244_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15719_  (.A(\reg_module/_08216_ ),
    .B(\reg_module/_08244_ ),
    .Y(\reg_module/_08245_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15720_  (.A(\reg_module/_08245_ ),
    .Y(\reg_module/_08246_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15721_  (.A(\reg_module/_08241_ ),
    .B(\reg_module/_07551_ ),
    .C(\reg_module/_08220_ ),
    .Y(\reg_module/_08247_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15722_  (.A(\reg_module/_08247_ ),
    .B(net1048),
    .Y(\reg_module/_08248_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15723_  (.A(\reg_module/_08246_ ),
    .B(\reg_module/_08248_ ),
    .Y(\reg_module/_00139_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15724_  (.A(\reg_module/_08178_ ),
    .X(\reg_module/_08249_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15725_  (.A(net2203),
    .Y(\reg_module/_08250_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15726_  (.A(\reg_module/_08249_ ),
    .B(\reg_module/_08250_ ),
    .Y(\reg_module/_08251_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15727_  (.A(\reg_module/_08251_ ),
    .Y(\reg_module/_08252_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15728_  (.A(\reg_module/_08186_ ),
    .X(\reg_module/_08253_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15729_  (.A(\reg_module/_08241_ ),
    .B(\reg_module/_07555_ ),
    .C(\reg_module/_08253_ ),
    .Y(\reg_module/_08254_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15730_  (.A(\reg_module/_08254_ ),
    .B(net1063),
    .Y(\reg_module/_08255_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15731_  (.A(\reg_module/_08252_ ),
    .B(\reg_module/_08255_ ),
    .Y(\reg_module/_00140_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15732_  (.A(net2175),
    .Y(\reg_module/_08256_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15733_  (.A(\reg_module/_08249_ ),
    .B(\reg_module/_08256_ ),
    .Y(\reg_module/_08257_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15734_  (.A(\reg_module/_08257_ ),
    .Y(\reg_module/_08258_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15735_  (.A(\reg_module/_08241_ ),
    .B(\reg_module/_07558_ ),
    .C(\reg_module/_08253_ ),
    .Y(\reg_module/_08259_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15736_  (.A(\reg_module/_08259_ ),
    .B(net1064),
    .Y(\reg_module/_08260_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15737_  (.A(\reg_module/_08258_ ),
    .B(\reg_module/_08260_ ),
    .Y(\reg_module/_00141_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15738_  (.A(\reg_module/gprf[142] ),
    .Y(\reg_module/_08261_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15739_  (.A(\reg_module/_08249_ ),
    .B(\reg_module/_08261_ ),
    .Y(\reg_module/_08262_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15740_  (.A(\reg_module/_08262_ ),
    .Y(\reg_module/_08263_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15741_  (.A(\reg_module/_08241_ ),
    .B(\reg_module/_07561_ ),
    .C(\reg_module/_08253_ ),
    .Y(\reg_module/_08264_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15742_  (.A(\reg_module/_08264_ ),
    .B(net1063),
    .Y(\reg_module/_08265_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15743_  (.A(\reg_module/_08263_ ),
    .B(\reg_module/_08265_ ),
    .Y(\reg_module/_00142_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15744_  (.A(\reg_module/gprf[143] ),
    .Y(\reg_module/_08266_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15745_  (.A(\reg_module/_08249_ ),
    .B(\reg_module/_08266_ ),
    .Y(\reg_module/_08267_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15746_  (.A(\reg_module/_08267_ ),
    .Y(\reg_module/_08268_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15747_  (.A(\reg_module/_08241_ ),
    .B(\reg_module/_07564_ ),
    .C(\reg_module/_08253_ ),
    .Y(\reg_module/_08269_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15748_  (.A(\reg_module/_08269_ ),
    .B(net1064),
    .Y(\reg_module/_08270_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15749_  (.A(\reg_module/_08268_ ),
    .B(\reg_module/_08270_ ),
    .Y(\reg_module/_00143_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15750_  (.A(\reg_module/gprf[144] ),
    .Y(\reg_module/_08271_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15751_  (.A(\reg_module/_08249_ ),
    .B(\reg_module/_08271_ ),
    .Y(\reg_module/_08272_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15752_  (.A(\reg_module/_08272_ ),
    .Y(\reg_module/_08273_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_15753_  (.A(\reg_module/_08184_ ),
    .X(\reg_module/_08274_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15754_  (.A(\reg_module/_08274_ ),
    .B(\reg_module/_07568_ ),
    .C(\reg_module/_08253_ ),
    .Y(\reg_module/_08275_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15755_  (.A(\reg_module/_08275_ ),
    .B(net1055),
    .Y(\reg_module/_08276_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15756_  (.A(\reg_module/_08273_ ),
    .B(\reg_module/_08276_ ),
    .Y(\reg_module/_00144_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15757_  (.A(\reg_module/gprf[145] ),
    .Y(\reg_module/_08277_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15758_  (.A(\reg_module/_08249_ ),
    .B(\reg_module/_08277_ ),
    .Y(\reg_module/_08278_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15759_  (.A(\reg_module/_08278_ ),
    .Y(\reg_module/_08279_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15760_  (.A(\reg_module/_08274_ ),
    .B(\reg_module/_07571_ ),
    .C(\reg_module/_08253_ ),
    .Y(\reg_module/_08280_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15761_  (.A(\reg_module/_08280_ ),
    .B(net1055),
    .Y(\reg_module/_08281_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15762_  (.A(\reg_module/_08279_ ),
    .B(\reg_module/_08281_ ),
    .Y(\reg_module/_00145_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15763_  (.A(\reg_module/_08178_ ),
    .X(\reg_module/_08282_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15764_  (.A(\reg_module/gprf[146] ),
    .Y(\reg_module/_08283_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15765_  (.A(\reg_module/_08282_ ),
    .B(\reg_module/_08283_ ),
    .Y(\reg_module/_08284_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15766_  (.A(\reg_module/_08284_ ),
    .Y(\reg_module/_08285_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15767_  (.A(\reg_module/_08186_ ),
    .X(\reg_module/_08286_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15768_  (.A(\reg_module/_08274_ ),
    .B(\reg_module/_07575_ ),
    .C(\reg_module/_08286_ ),
    .Y(\reg_module/_08287_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15769_  (.A(\reg_module/_08287_ ),
    .B(net1039),
    .Y(\reg_module/_08288_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15770_  (.A(\reg_module/_08285_ ),
    .B(\reg_module/_08288_ ),
    .Y(\reg_module/_00146_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15771_  (.A(\reg_module/gprf[147] ),
    .Y(\reg_module/_08289_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15772_  (.A(\reg_module/_08282_ ),
    .B(\reg_module/_08289_ ),
    .Y(\reg_module/_08290_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15773_  (.A(\reg_module/_08290_ ),
    .Y(\reg_module/_08291_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15774_  (.A(\reg_module/_08274_ ),
    .B(\reg_module/_07578_ ),
    .C(\reg_module/_08286_ ),
    .Y(\reg_module/_08292_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15775_  (.A(\reg_module/_08292_ ),
    .B(net1039),
    .Y(\reg_module/_08293_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15776_  (.A(\reg_module/_08291_ ),
    .B(\reg_module/_08293_ ),
    .Y(\reg_module/_00147_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15777_  (.A(\reg_module/gprf[148] ),
    .Y(\reg_module/_08294_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15778_  (.A(\reg_module/_08282_ ),
    .B(\reg_module/_08294_ ),
    .Y(\reg_module/_08295_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15779_  (.A(\reg_module/_08295_ ),
    .Y(\reg_module/_08296_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15780_  (.A(\reg_module/_08274_ ),
    .B(\reg_module/_07581_ ),
    .C(\reg_module/_08286_ ),
    .Y(\reg_module/_08297_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15781_  (.A(\reg_module/_08297_ ),
    .B(net1039),
    .Y(\reg_module/_08298_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15782_  (.A(\reg_module/_08296_ ),
    .B(\reg_module/_08298_ ),
    .Y(\reg_module/_00148_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15783_  (.A(\reg_module/gprf[149] ),
    .Y(\reg_module/_08299_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15784_  (.A(\reg_module/_08282_ ),
    .B(\reg_module/_08299_ ),
    .Y(\reg_module/_08300_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15785_  (.A(\reg_module/_08300_ ),
    .Y(\reg_module/_08301_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15786_  (.A(\reg_module/_08274_ ),
    .B(\reg_module/_07584_ ),
    .C(\reg_module/_08286_ ),
    .Y(\reg_module/_08302_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15787_  (.A(\reg_module/_08302_ ),
    .B(net1039),
    .Y(\reg_module/_08303_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15788_  (.A(\reg_module/_08301_ ),
    .B(\reg_module/_08303_ ),
    .Y(\reg_module/_00149_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15789_  (.A(net2209),
    .Y(\reg_module/_08304_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15790_  (.A(\reg_module/_08282_ ),
    .B(\reg_module/_08304_ ),
    .Y(\reg_module/_08305_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15791_  (.A(\reg_module/_08305_ ),
    .Y(\reg_module/_08306_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15792_  (.A(\reg_module/_08184_ ),
    .X(\reg_module/_08307_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15793_  (.A(\reg_module/_08307_ ),
    .B(\reg_module/_07588_ ),
    .C(\reg_module/_08286_ ),
    .Y(\reg_module/_08308_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15794_  (.A(\reg_module/_08308_ ),
    .B(net1038),
    .Y(\reg_module/_08309_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15795_  (.A(\reg_module/_08306_ ),
    .B(\reg_module/_08309_ ),
    .Y(\reg_module/_00150_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15796_  (.A(\reg_module/gprf[151] ),
    .Y(\reg_module/_08310_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15797_  (.A(\reg_module/_08282_ ),
    .B(\reg_module/_08310_ ),
    .Y(\reg_module/_08311_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15798_  (.A(\reg_module/_08311_ ),
    .Y(\reg_module/_08312_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15799_  (.A(\reg_module/_08307_ ),
    .B(\reg_module/_07591_ ),
    .C(\reg_module/_08286_ ),
    .Y(\reg_module/_08313_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15800_  (.A(\reg_module/_08313_ ),
    .B(net1038),
    .Y(\reg_module/_08314_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15801_  (.A(\reg_module/_08312_ ),
    .B(\reg_module/_08314_ ),
    .Y(\reg_module/_00151_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15802_  (.A(\reg_module/_08177_ ),
    .X(\reg_module/_08315_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15803_  (.A(\reg_module/gprf[152] ),
    .Y(\reg_module/_08316_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15804_  (.A(\reg_module/_08315_ ),
    .B(\reg_module/_08316_ ),
    .Y(\reg_module/_08317_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15805_  (.A(\reg_module/_08317_ ),
    .Y(\reg_module/_08318_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15806_  (.A(\reg_module/_08176_ ),
    .X(\reg_module/_08319_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15807_  (.A(\reg_module/_08307_ ),
    .B(\reg_module/_07595_ ),
    .C(\reg_module/_08319_ ),
    .Y(\reg_module/_08320_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15808_  (.A(\reg_module/_08320_ ),
    .B(net1006),
    .Y(\reg_module/_08321_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15809_  (.A(\reg_module/_08318_ ),
    .B(\reg_module/_08321_ ),
    .Y(\reg_module/_00152_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15810_  (.A(net2223),
    .Y(\reg_module/_08322_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15811_  (.A(\reg_module/_08315_ ),
    .B(\reg_module/_08322_ ),
    .Y(\reg_module/_08323_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15812_  (.A(\reg_module/_08323_ ),
    .Y(\reg_module/_08324_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15813_  (.A(\reg_module/_08307_ ),
    .B(\reg_module/_07598_ ),
    .C(\reg_module/_08319_ ),
    .Y(\reg_module/_08325_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15814_  (.A(\reg_module/_08325_ ),
    .B(net1006),
    .Y(\reg_module/_08326_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15815_  (.A(\reg_module/_08324_ ),
    .B(\reg_module/_08326_ ),
    .Y(\reg_module/_00153_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15816_  (.A(\reg_module/gprf[154] ),
    .Y(\reg_module/_08327_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15817_  (.A(\reg_module/_08315_ ),
    .B(\reg_module/_08327_ ),
    .Y(\reg_module/_08328_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15818_  (.A(\reg_module/_08328_ ),
    .Y(\reg_module/_08329_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15819_  (.A(\reg_module/_08307_ ),
    .B(\reg_module/_07601_ ),
    .C(\reg_module/_08319_ ),
    .Y(\reg_module/_08330_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15820_  (.A(\reg_module/_08330_ ),
    .B(net1005),
    .Y(\reg_module/_08331_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15821_  (.A(\reg_module/_08329_ ),
    .B(\reg_module/_08331_ ),
    .Y(\reg_module/_00154_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15822_  (.A(net2206),
    .Y(\reg_module/_08332_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15823_  (.A(\reg_module/_08315_ ),
    .B(\reg_module/_08332_ ),
    .Y(\reg_module/_08333_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15824_  (.A(\reg_module/_08333_ ),
    .Y(\reg_module/_08334_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15825_  (.A(\reg_module/_08307_ ),
    .B(\reg_module/_07604_ ),
    .C(\reg_module/_08319_ ),
    .Y(\reg_module/_08335_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15826_  (.A(\reg_module/_08335_ ),
    .B(net1005),
    .Y(\reg_module/_08336_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15827_  (.A(\reg_module/_08334_ ),
    .B(\reg_module/_08336_ ),
    .Y(\reg_module/_00155_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15828_  (.A(\reg_module/gprf[156] ),
    .Y(\reg_module/_08337_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15829_  (.A(\reg_module/_08315_ ),
    .B(\reg_module/_08337_ ),
    .Y(\reg_module/_08338_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15830_  (.A(\reg_module/_08338_ ),
    .Y(\reg_module/_08339_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_15831_  (.A(\reg_module/_08184_ ),
    .X(\reg_module/_08340_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15832_  (.A(\reg_module/_08340_ ),
    .B(\reg_module/_07607_ ),
    .C(\reg_module/_08319_ ),
    .Y(\reg_module/_08341_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15833_  (.A(\reg_module/_08341_ ),
    .B(net1004),
    .Y(\reg_module/_08342_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15834_  (.A(\reg_module/_08339_ ),
    .B(\reg_module/_08342_ ),
    .Y(\reg_module/_00156_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15835_  (.A(net2174),
    .Y(\reg_module/_08343_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15836_  (.A(\reg_module/_08315_ ),
    .B(\reg_module/_08343_ ),
    .Y(\reg_module/_08344_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15837_  (.A(\reg_module/_08344_ ),
    .Y(\reg_module/_08345_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15838_  (.A(\reg_module/_08340_ ),
    .B(\reg_module/_07610_ ),
    .C(\reg_module/_08319_ ),
    .Y(\reg_module/_08346_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15839_  (.A(\reg_module/_08346_ ),
    .B(net1004),
    .Y(\reg_module/_08347_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15840_  (.A(\reg_module/_08345_ ),
    .B(\reg_module/_08347_ ),
    .Y(\reg_module/_00157_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15841_  (.A(net2184),
    .Y(\reg_module/_08348_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15842_  (.A(\reg_module/_08178_ ),
    .B(\reg_module/_08348_ ),
    .Y(\reg_module/_08349_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15843_  (.A(\reg_module/_08349_ ),
    .Y(\reg_module/_08350_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15844_  (.A(\reg_module/_08340_ ),
    .B(\reg_module/_07613_ ),
    .C(\reg_module/_08186_ ),
    .Y(\reg_module/_08351_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15845_  (.A(\reg_module/_08351_ ),
    .B(net1010),
    .Y(\reg_module/_08352_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15846_  (.A(\reg_module/_08350_ ),
    .B(\reg_module/_08352_ ),
    .Y(\reg_module/_00158_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15847_  (.A(net2204),
    .Y(\reg_module/_08353_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15848_  (.A(\reg_module/_08178_ ),
    .B(\reg_module/_08353_ ),
    .Y(\reg_module/_08354_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15849_  (.A(\reg_module/_08354_ ),
    .Y(\reg_module/_08355_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_15850_  (.A(\reg_module/_08340_ ),
    .B(\reg_module/_07616_ ),
    .C(\reg_module/_08186_ ),
    .Y(\reg_module/_08356_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15851_  (.A(\reg_module/_08356_ ),
    .B(net1012),
    .Y(\reg_module/_08357_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15852_  (.A(\reg_module/_08355_ ),
    .B(\reg_module/_08357_ ),
    .Y(\reg_module/_00159_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15853_  (.A(\reg_module/_07628_ ),
    .B(\reg_module/_07816_ ),
    .Y(\reg_module/_08358_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15854_  (.A(\reg_module/_07625_ ),
    .B(\reg_module/_08358_ ),
    .Y(\reg_module/_08359_ ));
 sky130_fd_sc_hd__nand3_2 \reg_module/_15855_  (.A(\reg_module/_07620_ ),
    .B(\reg_module/_07624_ ),
    .C(\reg_module/_08359_ ),
    .Y(\reg_module/_08360_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_15856_  (.A(\reg_module/_08360_ ),
    .X(\reg_module/_08361_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15857_  (.A(\reg_module/_08361_ ),
    .X(\reg_module/_08362_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15858_  (.A(\reg_module/_08362_ ),
    .B(net1825),
    .Y(\reg_module/_08363_ ));
 sky130_fd_sc_hd__buf_8 \reg_module/_15859_  (.A(\reg_module/_07640_ ),
    .X(\reg_module/_08364_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15860_  (.A(\reg_module/_08364_ ),
    .X(\reg_module/_08365_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_15861_  (.A(\reg_module/_08358_ ),
    .Y(\reg_module/_08366_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_15862_  (.A(\reg_module/_08366_ ),
    .X(\reg_module/_08367_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15863_  (.A(\reg_module/_08367_ ),
    .X(\reg_module/_08368_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15864_  (.A(\reg_module/_08368_ ),
    .B(net318),
    .Y(\reg_module/_08369_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15865_  (.A(\reg_module/_08002_ ),
    .B(\reg_module/_08369_ ),
    .Y(\reg_module/_08370_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15866_  (.A(\reg_module/_08365_ ),
    .B(\reg_module/_08370_ ),
    .Y(\reg_module/_08371_ ));
 sky130_fd_sc_hd__buf_8 \reg_module/_15867_  (.A(\reg_module/_07993_ ),
    .X(\reg_module/_08372_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15868_  (.A(\reg_module/_08372_ ),
    .X(\reg_module/_08373_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15869_  (.A1(\reg_module/_08363_ ),
    .A2(\reg_module/_08371_ ),
    .B1(\reg_module/_08373_ ),
    .Y(\reg_module/_00160_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15870_  (.A(\reg_module/_08362_ ),
    .B(net1332),
    .Y(\reg_module/_08374_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15871_  (.A(\reg_module/_08368_ ),
    .B(net317),
    .Y(\reg_module/_08375_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15872_  (.A(\reg_module/_08002_ ),
    .B(\reg_module/_08375_ ),
    .Y(\reg_module/_08376_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15873_  (.A(\reg_module/_08365_ ),
    .B(\reg_module/_08376_ ),
    .Y(\reg_module/_08377_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15874_  (.A1(\reg_module/_08374_ ),
    .A2(\reg_module/_08377_ ),
    .B1(\reg_module/_08373_ ),
    .Y(\reg_module/_00161_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15875_  (.A(\reg_module/_08362_ ),
    .B(net1323),
    .Y(\reg_module/_08378_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15876_  (.A(\reg_module/_08368_ ),
    .B(net316),
    .Y(\reg_module/_08379_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15877_  (.A(\reg_module/_08002_ ),
    .B(\reg_module/_08379_ ),
    .Y(\reg_module/_08380_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15878_  (.A(\reg_module/_08365_ ),
    .B(\reg_module/_08380_ ),
    .Y(\reg_module/_08381_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15879_  (.A1(\reg_module/_08378_ ),
    .A2(\reg_module/_08381_ ),
    .B1(\reg_module/_08373_ ),
    .Y(\reg_module/_00162_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15880_  (.A(\reg_module/_08362_ ),
    .B(net1720),
    .Y(\reg_module/_08382_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15881_  (.A(\reg_module/_08368_ ),
    .B(net315),
    .Y(\reg_module/_08383_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15882_  (.A(\reg_module/_08002_ ),
    .B(\reg_module/_08383_ ),
    .Y(\reg_module/_08384_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15883_  (.A(\reg_module/_08365_ ),
    .B(\reg_module/_08384_ ),
    .Y(\reg_module/_08385_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15884_  (.A1(\reg_module/_08382_ ),
    .A2(\reg_module/_08385_ ),
    .B1(\reg_module/_08373_ ),
    .Y(\reg_module/_00163_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15885_  (.A(\reg_module/_08362_ ),
    .B(net1985),
    .Y(\reg_module/_08386_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15886_  (.A(\reg_module/_07645_ ),
    .X(\reg_module/_08387_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15887_  (.A(\reg_module/_08368_ ),
    .B(\wRegWrData[4] ),
    .Y(\reg_module/_08388_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15888_  (.A(\reg_module/_08387_ ),
    .B(\reg_module/_08388_ ),
    .Y(\reg_module/_08389_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15889_  (.A(\reg_module/_08365_ ),
    .B(\reg_module/_08389_ ),
    .Y(\reg_module/_08390_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15890_  (.A1(\reg_module/_08386_ ),
    .A2(\reg_module/_08390_ ),
    .B1(\reg_module/_08373_ ),
    .Y(\reg_module/_00164_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15891_  (.A(\reg_module/_08362_ ),
    .B(net2045),
    .Y(\reg_module/_08391_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15892_  (.A(\reg_module/_08368_ ),
    .B(net314),
    .Y(\reg_module/_08392_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15893_  (.A(\reg_module/_08387_ ),
    .B(\reg_module/_08392_ ),
    .Y(\reg_module/_08393_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15894_  (.A(\reg_module/_08365_ ),
    .B(\reg_module/_08393_ ),
    .Y(\reg_module/_08394_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15895_  (.A1(\reg_module/_08391_ ),
    .A2(\reg_module/_08394_ ),
    .B1(\reg_module/_08373_ ),
    .Y(\reg_module/_00165_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15896_  (.A(\reg_module/_08361_ ),
    .X(\reg_module/_08395_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15897_  (.A(\reg_module/_08395_ ),
    .B(net1543),
    .Y(\reg_module/_08396_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15898_  (.A(\reg_module/_08364_ ),
    .X(\reg_module/_08397_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15899_  (.A(\reg_module/_08367_ ),
    .X(\reg_module/_08398_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15900_  (.A(\reg_module/_08398_ ),
    .B(\wRegWrData[6] ),
    .Y(\reg_module/_08399_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_15901_  (.A(\reg_module/_08387_ ),
    .B(\reg_module/_08399_ ),
    .Y(\reg_module/_08400_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15902_  (.A(\reg_module/_08397_ ),
    .B(\reg_module/_08400_ ),
    .Y(\reg_module/_08401_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15903_  (.A(\reg_module/_08372_ ),
    .X(\reg_module/_08402_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15904_  (.A1(\reg_module/_08396_ ),
    .A2(\reg_module/_08401_ ),
    .B1(\reg_module/_08402_ ),
    .Y(\reg_module/_00166_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15905_  (.A(\reg_module/_08395_ ),
    .B(net1710),
    .Y(\reg_module/_08403_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15906_  (.A(\reg_module/_08398_ ),
    .B(net313),
    .Y(\reg_module/_08404_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_15907_  (.A(\reg_module/_08387_ ),
    .B(\reg_module/_08404_ ),
    .Y(\reg_module/_08405_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15908_  (.A(\reg_module/_08397_ ),
    .B(\reg_module/_08405_ ),
    .Y(\reg_module/_08406_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15909_  (.A1(\reg_module/_08403_ ),
    .A2(\reg_module/_08406_ ),
    .B1(\reg_module/_08402_ ),
    .Y(\reg_module/_00167_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15910_  (.A(\reg_module/_08395_ ),
    .B(net1675),
    .Y(\reg_module/_08407_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15911_  (.A(\reg_module/_08398_ ),
    .B(\wRegWrData[8] ),
    .Y(\reg_module/_08408_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_15912_  (.A(\reg_module/_08387_ ),
    .B(\reg_module/_08408_ ),
    .Y(\reg_module/_08409_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15913_  (.A(\reg_module/_08397_ ),
    .B(\reg_module/_08409_ ),
    .Y(\reg_module/_08410_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15914_  (.A1(\reg_module/_08407_ ),
    .A2(\reg_module/_08410_ ),
    .B1(\reg_module/_08402_ ),
    .Y(\reg_module/_00168_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15915_  (.A(\reg_module/_08395_ ),
    .B(net1609),
    .Y(\reg_module/_08411_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15916_  (.A(\reg_module/_08398_ ),
    .B(net312),
    .Y(\reg_module/_08412_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_15917_  (.A(\reg_module/_08387_ ),
    .B(\reg_module/_08412_ ),
    .Y(\reg_module/_08413_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15918_  (.A(\reg_module/_08397_ ),
    .B(\reg_module/_08413_ ),
    .Y(\reg_module/_08414_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15919_  (.A1(\reg_module/_08411_ ),
    .A2(\reg_module/_08414_ ),
    .B1(\reg_module/_08402_ ),
    .Y(\reg_module/_00169_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15920_  (.A(\reg_module/_08395_ ),
    .B(net1773),
    .Y(\reg_module/_08415_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15921_  (.A(\reg_module/_07645_ ),
    .X(\reg_module/_08416_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15922_  (.A(\reg_module/_08398_ ),
    .B(net311),
    .Y(\reg_module/_08417_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_15923_  (.A(\reg_module/_08416_ ),
    .B(\reg_module/_08417_ ),
    .Y(\reg_module/_08418_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15924_  (.A(\reg_module/_08397_ ),
    .B(\reg_module/_08418_ ),
    .Y(\reg_module/_08419_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15925_  (.A1(\reg_module/_08415_ ),
    .A2(\reg_module/_08419_ ),
    .B1(\reg_module/_08402_ ),
    .Y(\reg_module/_00170_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15926_  (.A(\reg_module/_08395_ ),
    .B(net1420),
    .Y(\reg_module/_08420_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15927_  (.A(\reg_module/_08398_ ),
    .B(net310),
    .Y(\reg_module/_08421_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_15928_  (.A(\reg_module/_08416_ ),
    .B(\reg_module/_08421_ ),
    .Y(\reg_module/_08422_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15929_  (.A(\reg_module/_08397_ ),
    .B(\reg_module/_08422_ ),
    .Y(\reg_module/_08423_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15930_  (.A1(\reg_module/_08420_ ),
    .A2(\reg_module/_08423_ ),
    .B1(\reg_module/_08402_ ),
    .Y(\reg_module/_00171_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15931_  (.A(\reg_module/_08361_ ),
    .X(\reg_module/_08424_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15932_  (.A(\reg_module/_08424_ ),
    .B(net1861),
    .Y(\reg_module/_08425_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15933_  (.A(\reg_module/_08364_ ),
    .X(\reg_module/_08426_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15934_  (.A(\reg_module/_08367_ ),
    .X(\reg_module/_08427_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15935_  (.A(\reg_module/_08427_ ),
    .B(\wRegWrData[12] ),
    .Y(\reg_module/_08428_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_15936_  (.A(\reg_module/_08416_ ),
    .B(\reg_module/_08428_ ),
    .Y(\reg_module/_08429_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15937_  (.A(\reg_module/_08426_ ),
    .B(\reg_module/_08429_ ),
    .Y(\reg_module/_08430_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15938_  (.A(\reg_module/_08372_ ),
    .X(\reg_module/_08431_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15939_  (.A1(\reg_module/_08425_ ),
    .A2(\reg_module/_08430_ ),
    .B1(\reg_module/_08431_ ),
    .Y(\reg_module/_00172_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15940_  (.A(\reg_module/_08424_ ),
    .B(net1973),
    .Y(\reg_module/_08432_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15941_  (.A(\reg_module/_08427_ ),
    .B(net309),
    .Y(\reg_module/_08433_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_15942_  (.A(\reg_module/_08416_ ),
    .B(\reg_module/_08433_ ),
    .Y(\reg_module/_08434_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15943_  (.A(\reg_module/_08426_ ),
    .B(\reg_module/_08434_ ),
    .Y(\reg_module/_08435_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15944_  (.A1(\reg_module/_08432_ ),
    .A2(\reg_module/_08435_ ),
    .B1(\reg_module/_08431_ ),
    .Y(\reg_module/_00173_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15945_  (.A(\reg_module/_08424_ ),
    .B(net1915),
    .Y(\reg_module/_08436_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15946_  (.A(\reg_module/_08427_ ),
    .B(net308),
    .Y(\reg_module/_08437_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15947_  (.A(\reg_module/_08416_ ),
    .B(\reg_module/_08437_ ),
    .Y(\reg_module/_08438_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15948_  (.A(\reg_module/_08426_ ),
    .B(\reg_module/_08438_ ),
    .Y(\reg_module/_08439_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15949_  (.A1(\reg_module/_08436_ ),
    .A2(\reg_module/_08439_ ),
    .B1(\reg_module/_08431_ ),
    .Y(\reg_module/_00174_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15950_  (.A(\reg_module/_08424_ ),
    .B(net1691),
    .Y(\reg_module/_08440_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15951_  (.A(\reg_module/_08427_ ),
    .B(net306),
    .Y(\reg_module/_08441_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15952_  (.A(\reg_module/_08416_ ),
    .B(\reg_module/_08441_ ),
    .Y(\reg_module/_08442_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15953_  (.A(\reg_module/_08426_ ),
    .B(\reg_module/_08442_ ),
    .Y(\reg_module/_08443_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15954_  (.A1(\reg_module/_08440_ ),
    .A2(\reg_module/_08443_ ),
    .B1(\reg_module/_08431_ ),
    .Y(\reg_module/_00175_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15955_  (.A(\reg_module/_08424_ ),
    .B(net1605),
    .Y(\reg_module/_08444_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15956_  (.A(\reg_module/_07645_ ),
    .X(\reg_module/_08445_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15957_  (.A(\reg_module/_08427_ ),
    .B(\wRegWrData[16] ),
    .Y(\reg_module/_08446_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_15958_  (.A(\reg_module/_08445_ ),
    .B(\reg_module/_08446_ ),
    .Y(\reg_module/_08447_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15959_  (.A(\reg_module/_08426_ ),
    .B(\reg_module/_08447_ ),
    .Y(\reg_module/_08448_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15960_  (.A1(\reg_module/_08444_ ),
    .A2(\reg_module/_08448_ ),
    .B1(\reg_module/_08431_ ),
    .Y(\reg_module/_00176_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15961_  (.A(\reg_module/_08424_ ),
    .B(net1659),
    .Y(\reg_module/_08449_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15962_  (.A(\reg_module/_08427_ ),
    .B(net305),
    .Y(\reg_module/_08450_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15963_  (.A(\reg_module/_08445_ ),
    .B(\reg_module/_08450_ ),
    .Y(\reg_module/_08451_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15964_  (.A(\reg_module/_08426_ ),
    .B(\reg_module/_08451_ ),
    .Y(\reg_module/_08452_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15965_  (.A1(\reg_module/_08449_ ),
    .A2(\reg_module/_08452_ ),
    .B1(\reg_module/_08431_ ),
    .Y(\reg_module/_00177_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15966_  (.A(\reg_module/_08361_ ),
    .X(\reg_module/_08453_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15967_  (.A(\reg_module/_08453_ ),
    .B(net1797),
    .Y(\reg_module/_08454_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15968_  (.A(\reg_module/_08364_ ),
    .X(\reg_module/_08455_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15969_  (.A(\reg_module/_08367_ ),
    .X(\reg_module/_08456_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15970_  (.A(\reg_module/_08456_ ),
    .B(net304),
    .Y(\reg_module/_08457_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15971_  (.A(\reg_module/_08445_ ),
    .B(\reg_module/_08457_ ),
    .Y(\reg_module/_08458_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15972_  (.A(\reg_module/_08455_ ),
    .B(\reg_module/_08458_ ),
    .Y(\reg_module/_08459_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_15973_  (.A(\reg_module/_08372_ ),
    .X(\reg_module/_08460_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15974_  (.A1(\reg_module/_08454_ ),
    .A2(\reg_module/_08459_ ),
    .B1(\reg_module/_08460_ ),
    .Y(\reg_module/_00178_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15975_  (.A(\reg_module/_08453_ ),
    .B(net1600),
    .Y(\reg_module/_08461_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15976_  (.A(\reg_module/_08456_ ),
    .B(net303),
    .Y(\reg_module/_08462_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15977_  (.A(\reg_module/_08445_ ),
    .B(\reg_module/_08462_ ),
    .Y(\reg_module/_08463_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15978_  (.A(\reg_module/_08455_ ),
    .B(\reg_module/_08463_ ),
    .Y(\reg_module/_08464_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15979_  (.A1(\reg_module/_08461_ ),
    .A2(\reg_module/_08464_ ),
    .B1(\reg_module/_08460_ ),
    .Y(\reg_module/_00179_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15980_  (.A(\reg_module/_08453_ ),
    .B(net1656),
    .Y(\reg_module/_08465_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15981_  (.A(\reg_module/_08456_ ),
    .B(net302),
    .Y(\reg_module/_08466_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15982_  (.A(\reg_module/_08445_ ),
    .B(\reg_module/_08466_ ),
    .Y(\reg_module/_08467_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15983_  (.A(\reg_module/_08455_ ),
    .B(\reg_module/_08467_ ),
    .Y(\reg_module/_08468_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15984_  (.A1(\reg_module/_08465_ ),
    .A2(\reg_module/_08468_ ),
    .B1(\reg_module/_08460_ ),
    .Y(\reg_module/_00180_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15985_  (.A(\reg_module/_08453_ ),
    .B(net1528),
    .Y(\reg_module/_08469_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15986_  (.A(\reg_module/_08456_ ),
    .B(net301),
    .Y(\reg_module/_08470_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15987_  (.A(\reg_module/_08445_ ),
    .B(\reg_module/_08470_ ),
    .Y(\reg_module/_08471_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15988_  (.A(\reg_module/_08455_ ),
    .B(\reg_module/_08471_ ),
    .Y(\reg_module/_08472_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15989_  (.A1(\reg_module/_08469_ ),
    .A2(\reg_module/_08472_ ),
    .B1(\reg_module/_08460_ ),
    .Y(\reg_module/_00181_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15990_  (.A(\reg_module/_08453_ ),
    .B(net1541),
    .Y(\reg_module/_08473_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_15991_  (.A(\reg_module/_07645_ ),
    .X(\reg_module/_08474_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15992_  (.A(\reg_module/_08456_ ),
    .B(net300),
    .Y(\reg_module/_08475_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15993_  (.A(\reg_module/_08474_ ),
    .B(\reg_module/_08475_ ),
    .Y(\reg_module/_08476_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15994_  (.A(\reg_module/_08455_ ),
    .B(\reg_module/_08476_ ),
    .Y(\reg_module/_08477_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_15995_  (.A1(\reg_module/_08473_ ),
    .A2(\reg_module/_08477_ ),
    .B1(\reg_module/_08460_ ),
    .Y(\reg_module/_00182_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15996_  (.A(\reg_module/_08453_ ),
    .B(net1672),
    .Y(\reg_module/_08478_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15997_  (.A(\reg_module/_08456_ ),
    .B(net299),
    .Y(\reg_module/_08479_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_15998_  (.A(\reg_module/_08474_ ),
    .B(\reg_module/_08479_ ),
    .Y(\reg_module/_08480_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_15999_  (.A(\reg_module/_08455_ ),
    .B(\reg_module/_08480_ ),
    .Y(\reg_module/_08481_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16000_  (.A1(\reg_module/_08478_ ),
    .A2(\reg_module/_08481_ ),
    .B1(\reg_module/_08460_ ),
    .Y(\reg_module/_00183_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16001_  (.A(\reg_module/_08360_ ),
    .X(\reg_module/_08482_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16002_  (.A(\reg_module/_08482_ ),
    .B(net1436),
    .Y(\reg_module/_08483_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16003_  (.A(\reg_module/_08364_ ),
    .X(\reg_module/_08484_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16004_  (.A(\reg_module/_08366_ ),
    .X(\reg_module/_08485_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16005_  (.A(\reg_module/_08485_ ),
    .B(net298),
    .Y(\reg_module/_08486_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16006_  (.A(\reg_module/_08474_ ),
    .B(\reg_module/_08486_ ),
    .Y(\reg_module/_08487_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16007_  (.A(\reg_module/_08484_ ),
    .B(\reg_module/_08487_ ),
    .Y(\reg_module/_08488_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16008_  (.A(\reg_module/_08372_ ),
    .X(\reg_module/_08489_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16009_  (.A1(\reg_module/_08483_ ),
    .A2(\reg_module/_08488_ ),
    .B1(\reg_module/_08489_ ),
    .Y(\reg_module/_00184_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16010_  (.A(\reg_module/_08482_ ),
    .B(net1310),
    .Y(\reg_module/_08490_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16011_  (.A(\reg_module/_08485_ ),
    .B(net296),
    .Y(\reg_module/_08491_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16012_  (.A(\reg_module/_08474_ ),
    .B(\reg_module/_08491_ ),
    .Y(\reg_module/_08492_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16013_  (.A(\reg_module/_08484_ ),
    .B(\reg_module/_08492_ ),
    .Y(\reg_module/_08493_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16014_  (.A1(\reg_module/_08490_ ),
    .A2(\reg_module/_08493_ ),
    .B1(\reg_module/_08489_ ),
    .Y(\reg_module/_00185_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16015_  (.A(\reg_module/_08482_ ),
    .B(net1412),
    .Y(\reg_module/_08494_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16016_  (.A(\reg_module/_08485_ ),
    .B(net294),
    .Y(\reg_module/_08495_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16017_  (.A(\reg_module/_08474_ ),
    .B(\reg_module/_08495_ ),
    .Y(\reg_module/_08496_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16018_  (.A(\reg_module/_08484_ ),
    .B(\reg_module/_08496_ ),
    .Y(\reg_module/_08497_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16019_  (.A1(\reg_module/_08494_ ),
    .A2(\reg_module/_08497_ ),
    .B1(\reg_module/_08489_ ),
    .Y(\reg_module/_00186_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16020_  (.A(\reg_module/_08482_ ),
    .B(net1297),
    .Y(\reg_module/_08498_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16021_  (.A(\reg_module/_08485_ ),
    .B(net293),
    .Y(\reg_module/_08499_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16022_  (.A(\reg_module/_08474_ ),
    .B(\reg_module/_08499_ ),
    .Y(\reg_module/_08500_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16023_  (.A(\reg_module/_08484_ ),
    .B(\reg_module/_08500_ ),
    .Y(\reg_module/_08501_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16024_  (.A1(\reg_module/_08498_ ),
    .A2(\reg_module/_08501_ ),
    .B1(\reg_module/_08489_ ),
    .Y(\reg_module/_00187_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16025_  (.A(\reg_module/_08482_ ),
    .B(net1257),
    .Y(\reg_module/_08502_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16026_  (.A(\reg_module/_07644_ ),
    .X(\reg_module/_08503_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16027_  (.A(\reg_module/_08485_ ),
    .B(net292),
    .Y(\reg_module/_08504_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16028_  (.A(\reg_module/_08503_ ),
    .B(\reg_module/_08504_ ),
    .Y(\reg_module/_08505_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16029_  (.A(\reg_module/_08484_ ),
    .B(\reg_module/_08505_ ),
    .Y(\reg_module/_08506_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16030_  (.A1(\reg_module/_08502_ ),
    .A2(\reg_module/_08506_ ),
    .B1(\reg_module/_08489_ ),
    .Y(\reg_module/_00188_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16031_  (.A(\reg_module/_08482_ ),
    .B(net1487),
    .Y(\reg_module/_08507_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16032_  (.A(\reg_module/_08485_ ),
    .B(net290),
    .Y(\reg_module/_08508_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16033_  (.A(\reg_module/_08503_ ),
    .B(\reg_module/_08508_ ),
    .Y(\reg_module/_08509_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16034_  (.A(\reg_module/_08484_ ),
    .B(\reg_module/_08509_ ),
    .Y(\reg_module/_08510_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16035_  (.A1(\reg_module/_08507_ ),
    .A2(\reg_module/_08510_ ),
    .B1(\reg_module/_08489_ ),
    .Y(\reg_module/_00189_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16036_  (.A(\reg_module/_08361_ ),
    .B(net1590),
    .Y(\reg_module/_08511_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16037_  (.A(\reg_module/_08364_ ),
    .X(\reg_module/_08512_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16038_  (.A(\reg_module/_08367_ ),
    .B(net289),
    .Y(\reg_module/_08513_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16039_  (.A(\reg_module/_08503_ ),
    .B(\reg_module/_08513_ ),
    .Y(\reg_module/_08514_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16040_  (.A(\reg_module/_08512_ ),
    .B(\reg_module/_08514_ ),
    .Y(\reg_module/_08515_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16041_  (.A(\reg_module/_08372_ ),
    .X(\reg_module/_08516_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16042_  (.A1(\reg_module/_08511_ ),
    .A2(\reg_module/_08515_ ),
    .B1(\reg_module/_08516_ ),
    .Y(\reg_module/_00190_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16043_  (.A(\reg_module/_08361_ ),
    .B(net1592),
    .Y(\reg_module/_08517_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16044_  (.A(\reg_module/_08367_ ),
    .B(net287),
    .Y(\reg_module/_08518_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16045_  (.A(\reg_module/_08503_ ),
    .B(\reg_module/_08518_ ),
    .Y(\reg_module/_08519_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16046_  (.A(\reg_module/_08512_ ),
    .B(\reg_module/_08519_ ),
    .Y(\reg_module/_08520_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16047_  (.A1(\reg_module/_08517_ ),
    .A2(\reg_module/_08520_ ),
    .B1(\reg_module/_08516_ ),
    .Y(\reg_module/_00191_ ));
 sky130_fd_sc_hd__and3_1 \reg_module/_16048_  (.A(\reg_module/_07808_ ),
    .B(net963),
    .C(\reg_module/_07817_ ),
    .X(\reg_module/_08521_ ));
 sky130_fd_sc_hd__nand3_2 \reg_module/_16049_  (.A(\reg_module/_07620_ ),
    .B(\reg_module/_07624_ ),
    .C(\reg_module/_08521_ ),
    .Y(\reg_module/_08522_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_16050_  (.A(\reg_module/_08522_ ),
    .X(\reg_module/_08523_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16051_  (.A(\reg_module/_08523_ ),
    .X(\reg_module/_08524_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16052_  (.A(\reg_module/_08524_ ),
    .B(net1563),
    .Y(\reg_module/_08525_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_16053_  (.A(\reg_module/_07625_ ),
    .X(\reg_module/_08526_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16054_  (.A(\reg_module/_08526_ ),
    .X(\reg_module/_08527_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16055_  (.A(\reg_module/_08527_ ),
    .B(net977),
    .C(\reg_module/_07821_ ),
    .Y(\reg_module/_08528_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16056_  (.A(\reg_module/_08512_ ),
    .B(\reg_module/_08528_ ),
    .Y(\reg_module/_08529_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16057_  (.A1(\reg_module/_08525_ ),
    .A2(\reg_module/_08529_ ),
    .B1(\reg_module/_08516_ ),
    .Y(\reg_module/_00192_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16058_  (.A(\reg_module/_08524_ ),
    .B(net1610),
    .Y(\reg_module/_08530_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16059_  (.A(\reg_module/_08527_ ),
    .B(net977),
    .C(\reg_module/_07826_ ),
    .Y(\reg_module/_08531_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16060_  (.A(\reg_module/_08512_ ),
    .B(\reg_module/_08531_ ),
    .Y(\reg_module/_08532_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16061_  (.A1(\reg_module/_08530_ ),
    .A2(\reg_module/_08532_ ),
    .B1(\reg_module/_08516_ ),
    .Y(\reg_module/_00193_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16062_  (.A(\reg_module/_08524_ ),
    .B(net1601),
    .Y(\reg_module/_08533_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16063_  (.A(\reg_module/_08527_ ),
    .B(net981),
    .C(\reg_module/_07831_ ),
    .Y(\reg_module/_08534_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16064_  (.A(\reg_module/_08512_ ),
    .B(net285),
    .Y(\reg_module/_08535_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16065_  (.A1(\reg_module/_08533_ ),
    .A2(\reg_module/_08535_ ),
    .B1(\reg_module/_08516_ ),
    .Y(\reg_module/_00194_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16066_  (.A(\reg_module/_08524_ ),
    .B(net1891),
    .Y(\reg_module/_08536_ ));
 sky130_fd_sc_hd__nor3_2 \reg_module/_16067_  (.A(\reg_module/_08527_ ),
    .B(net981),
    .C(\reg_module/_07836_ ),
    .Y(\reg_module/_08537_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16068_  (.A(\reg_module/_08512_ ),
    .B(\reg_module/_08537_ ),
    .Y(\reg_module/_08538_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16069_  (.A1(\reg_module/_08536_ ),
    .A2(\reg_module/_08538_ ),
    .B1(\reg_module/_08516_ ),
    .Y(\reg_module/_00195_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16070_  (.A(\reg_module/_08524_ ),
    .B(net1422),
    .Y(\reg_module/_08539_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_16071_  (.A(\reg_module/_08183_ ),
    .X(\reg_module/_08540_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16072_  (.A(\reg_module/_08540_ ),
    .X(\reg_module/_08541_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16073_  (.A(\reg_module/_08527_ ),
    .B(net984),
    .C(\reg_module/_07844_ ),
    .Y(\reg_module/_08542_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16074_  (.A(\reg_module/_08541_ ),
    .B(net284),
    .Y(\reg_module/_08543_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16075_  (.A(\reg_module/_07993_ ),
    .X(\reg_module/_08544_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16076_  (.A(\reg_module/_08544_ ),
    .X(\reg_module/_08545_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16077_  (.A1(\reg_module/_08539_ ),
    .A2(\reg_module/_08543_ ),
    .B1(\reg_module/_08545_ ),
    .Y(\reg_module/_00196_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16078_  (.A(\reg_module/_08524_ ),
    .B(net1296),
    .Y(\reg_module/_08546_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16079_  (.A(\reg_module/_08527_ ),
    .B(net984),
    .C(\reg_module/_07850_ ),
    .Y(\reg_module/_08547_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16080_  (.A(\reg_module/_08541_ ),
    .B(net283),
    .Y(\reg_module/_08548_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16081_  (.A1(\reg_module/_08546_ ),
    .A2(\reg_module/_08548_ ),
    .B1(\reg_module/_08545_ ),
    .Y(\reg_module/_00197_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16082_  (.A(\reg_module/_08523_ ),
    .X(\reg_module/_08549_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16083_  (.A(\reg_module/_08549_ ),
    .B(net1553),
    .Y(\reg_module/_08550_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16084_  (.A(\reg_module/_08526_ ),
    .X(\reg_module/_08551_ ));
 sky130_fd_sc_hd__nor3_2 \reg_module/_16085_  (.A(\reg_module/_08551_ ),
    .B(net982),
    .C(\reg_module/_07858_ ),
    .Y(\reg_module/_08552_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16086_  (.A(\reg_module/_08541_ ),
    .B(\reg_module/_08552_ ),
    .Y(\reg_module/_08553_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16087_  (.A1(\reg_module/_08550_ ),
    .A2(\reg_module/_08553_ ),
    .B1(\reg_module/_08545_ ),
    .Y(\reg_module/_00198_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16088_  (.A(\reg_module/_08549_ ),
    .B(net1751),
    .Y(\reg_module/_08554_ ));
 sky130_fd_sc_hd__nor3_2 \reg_module/_16089_  (.A(\reg_module/_08551_ ),
    .B(net982),
    .C(\reg_module/_07863_ ),
    .Y(\reg_module/_08555_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16090_  (.A(\reg_module/_08541_ ),
    .B(\reg_module/_08555_ ),
    .Y(\reg_module/_08556_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16091_  (.A1(\reg_module/_08554_ ),
    .A2(\reg_module/_08556_ ),
    .B1(\reg_module/_08545_ ),
    .Y(\reg_module/_00199_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16092_  (.A(\reg_module/_08549_ ),
    .B(net1577),
    .Y(\reg_module/_08557_ ));
 sky130_fd_sc_hd__nor3_2 \reg_module/_16093_  (.A(\reg_module/_08551_ ),
    .B(net982),
    .C(\reg_module/_07868_ ),
    .Y(\reg_module/_08558_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16094_  (.A(\reg_module/_08541_ ),
    .B(\reg_module/_08558_ ),
    .Y(\reg_module/_08559_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16095_  (.A1(\reg_module/_08557_ ),
    .A2(\reg_module/_08559_ ),
    .B1(\reg_module/_08545_ ),
    .Y(\reg_module/_00200_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16096_  (.A(\reg_module/_08549_ ),
    .B(net1694),
    .Y(\reg_module/_08560_ ));
 sky130_fd_sc_hd__nor3_2 \reg_module/_16097_  (.A(\reg_module/_08551_ ),
    .B(net983),
    .C(\reg_module/_07873_ ),
    .Y(\reg_module/_08561_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16098_  (.A(\reg_module/_08541_ ),
    .B(\reg_module/_08561_ ),
    .Y(\reg_module/_08562_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16099_  (.A1(\reg_module/_08560_ ),
    .A2(\reg_module/_08562_ ),
    .B1(\reg_module/_08545_ ),
    .Y(\reg_module/_00201_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16100_  (.A(\reg_module/_08549_ ),
    .B(net1955),
    .Y(\reg_module/_08563_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16101_  (.A(\reg_module/_08540_ ),
    .X(\reg_module/_08564_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16102_  (.A(\reg_module/_08551_ ),
    .B(net983),
    .C(\reg_module/_07880_ ),
    .Y(\reg_module/_08565_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16103_  (.A(\reg_module/_08564_ ),
    .B(\reg_module/_08565_ ),
    .Y(\reg_module/_08566_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16104_  (.A(\reg_module/_08544_ ),
    .X(\reg_module/_08567_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16105_  (.A1(\reg_module/_08563_ ),
    .A2(\reg_module/_08566_ ),
    .B1(\reg_module/_08567_ ),
    .Y(\reg_module/_00202_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16106_  (.A(\reg_module/_08549_ ),
    .B(net1637),
    .Y(\reg_module/_08568_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16107_  (.A(\reg_module/_08551_ ),
    .B(net983),
    .C(\reg_module/_07886_ ),
    .Y(\reg_module/_08569_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16108_  (.A(\reg_module/_08564_ ),
    .B(\reg_module/_08569_ ),
    .Y(\reg_module/_08570_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16109_  (.A1(\reg_module/_08568_ ),
    .A2(\reg_module/_08570_ ),
    .B1(\reg_module/_08567_ ),
    .Y(\reg_module/_00203_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16110_  (.A(\reg_module/_08523_ ),
    .X(\reg_module/_08571_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16111_  (.A(\reg_module/_08571_ ),
    .B(net1756),
    .Y(\reg_module/_08572_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16112_  (.A(\reg_module/_07625_ ),
    .X(\reg_module/_08573_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_16113_  (.A(\reg_module/_08573_ ),
    .X(\reg_module/_08574_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16114_  (.A(\reg_module/_08574_ ),
    .B(net988),
    .C(\reg_module/_07894_ ),
    .Y(\reg_module/_08575_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16115_  (.A(\reg_module/_08564_ ),
    .B(\reg_module/_08575_ ),
    .Y(\reg_module/_08576_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16116_  (.A1(\reg_module/_08572_ ),
    .A2(\reg_module/_08576_ ),
    .B1(\reg_module/_08567_ ),
    .Y(\reg_module/_00204_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16117_  (.A(\reg_module/_08571_ ),
    .B(net1863),
    .Y(\reg_module/_08577_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16118_  (.A(\reg_module/_08574_ ),
    .B(net988),
    .C(\reg_module/_07899_ ),
    .Y(\reg_module/_08578_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16119_  (.A(\reg_module/_08564_ ),
    .B(\reg_module/_08578_ ),
    .Y(\reg_module/_08579_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16120_  (.A1(\reg_module/_08577_ ),
    .A2(\reg_module/_08579_ ),
    .B1(\reg_module/_08567_ ),
    .Y(\reg_module/_00205_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16121_  (.A(\reg_module/_08571_ ),
    .B(net1475),
    .Y(\reg_module/_08580_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16122_  (.A(\reg_module/_08574_ ),
    .B(net988),
    .C(\reg_module/_07904_ ),
    .Y(\reg_module/_08581_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16123_  (.A(\reg_module/_08564_ ),
    .B(\reg_module/_08581_ ),
    .Y(\reg_module/_08582_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16124_  (.A1(\reg_module/_08580_ ),
    .A2(\reg_module/_08582_ ),
    .B1(\reg_module/_08567_ ),
    .Y(\reg_module/_00206_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16125_  (.A(\reg_module/_08571_ ),
    .B(net1492),
    .Y(\reg_module/_08583_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16126_  (.A(\reg_module/_08574_ ),
    .B(net988),
    .C(\reg_module/_07909_ ),
    .Y(\reg_module/_08584_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16127_  (.A(\reg_module/_08564_ ),
    .B(\reg_module/_08584_ ),
    .Y(\reg_module/_08585_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16128_  (.A1(\reg_module/_08583_ ),
    .A2(\reg_module/_08585_ ),
    .B1(\reg_module/_08567_ ),
    .Y(\reg_module/_00207_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16129_  (.A(\reg_module/_08571_ ),
    .B(net1442),
    .Y(\reg_module/_08586_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16130_  (.A(\reg_module/_08540_ ),
    .X(\reg_module/_08587_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16131_  (.A(\reg_module/_08574_ ),
    .B(net988),
    .C(\reg_module/_07916_ ),
    .Y(\reg_module/_08588_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16132_  (.A(\reg_module/_08587_ ),
    .B(\reg_module/_08588_ ),
    .Y(\reg_module/_08589_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16133_  (.A(\reg_module/_08544_ ),
    .X(\reg_module/_08590_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16134_  (.A1(\reg_module/_08586_ ),
    .A2(\reg_module/_08589_ ),
    .B1(\reg_module/_08590_ ),
    .Y(\reg_module/_00208_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16135_  (.A(\reg_module/_08571_ ),
    .B(net1452),
    .Y(\reg_module/_08591_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16136_  (.A(\reg_module/_08574_ ),
    .B(net989),
    .C(\reg_module/_07922_ ),
    .Y(\reg_module/_08592_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16137_  (.A(\reg_module/_08587_ ),
    .B(\reg_module/_08592_ ),
    .Y(\reg_module/_08593_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16138_  (.A1(\reg_module/_08591_ ),
    .A2(\reg_module/_08593_ ),
    .B1(\reg_module/_08590_ ),
    .Y(\reg_module/_00209_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16139_  (.A(\reg_module/_08523_ ),
    .X(\reg_module/_08594_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16140_  (.A(\reg_module/_08594_ ),
    .B(net1737),
    .Y(\reg_module/_08595_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16141_  (.A(\reg_module/_08573_ ),
    .X(\reg_module/_08596_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16142_  (.A(\reg_module/_08596_ ),
    .B(net990),
    .C(\reg_module/_07930_ ),
    .Y(\reg_module/_08597_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16143_  (.A(\reg_module/_08587_ ),
    .B(\reg_module/_08597_ ),
    .Y(\reg_module/_08598_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16144_  (.A1(\reg_module/_08595_ ),
    .A2(\reg_module/_08598_ ),
    .B1(\reg_module/_08590_ ),
    .Y(\reg_module/_00210_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16145_  (.A(\reg_module/_08594_ ),
    .B(net1573),
    .Y(\reg_module/_08599_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16146_  (.A(\reg_module/_08596_ ),
    .B(net990),
    .C(\reg_module/_07935_ ),
    .Y(\reg_module/_08600_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16147_  (.A(\reg_module/_08587_ ),
    .B(\reg_module/_08600_ ),
    .Y(\reg_module/_08601_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16148_  (.A1(\reg_module/_08599_ ),
    .A2(\reg_module/_08601_ ),
    .B1(\reg_module/_08590_ ),
    .Y(\reg_module/_00211_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16149_  (.A(\reg_module/_08594_ ),
    .B(net1306),
    .Y(\reg_module/_08602_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16150_  (.A(\reg_module/_08596_ ),
    .B(net986),
    .C(\reg_module/_07940_ ),
    .Y(\reg_module/_08603_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16151_  (.A(\reg_module/_08587_ ),
    .B(net282),
    .Y(\reg_module/_08604_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16152_  (.A1(\reg_module/_08602_ ),
    .A2(\reg_module/_08604_ ),
    .B1(\reg_module/_08590_ ),
    .Y(\reg_module/_00212_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16153_  (.A(\reg_module/_08594_ ),
    .B(net1650),
    .Y(\reg_module/_08605_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16154_  (.A(\reg_module/_08596_ ),
    .B(net986),
    .C(\reg_module/_07945_ ),
    .Y(\reg_module/_08606_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16155_  (.A(\reg_module/_08587_ ),
    .B(net281),
    .Y(\reg_module/_08607_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16156_  (.A1(\reg_module/_08605_ ),
    .A2(\reg_module/_08607_ ),
    .B1(\reg_module/_08590_ ),
    .Y(\reg_module/_00213_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16157_  (.A(\reg_module/_08594_ ),
    .B(net1623),
    .Y(\reg_module/_08608_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16158_  (.A(\reg_module/_08540_ ),
    .X(\reg_module/_08609_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16159_  (.A(\reg_module/_08596_ ),
    .B(net986),
    .C(\reg_module/_07952_ ),
    .Y(\reg_module/_08610_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16160_  (.A(\reg_module/_08609_ ),
    .B(\reg_module/_08610_ ),
    .Y(\reg_module/_08611_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_16161_  (.A(\reg_module/_08544_ ),
    .X(\reg_module/_08612_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16162_  (.A1(\reg_module/_08608_ ),
    .A2(\reg_module/_08611_ ),
    .B1(\reg_module/_08612_ ),
    .Y(\reg_module/_00214_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16163_  (.A(\reg_module/_08594_ ),
    .B(net1772),
    .Y(\reg_module/_08613_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16164_  (.A(\reg_module/_08596_ ),
    .B(net986),
    .C(\reg_module/_07958_ ),
    .Y(\reg_module/_08614_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16165_  (.A(\reg_module/_08609_ ),
    .B(\reg_module/_08614_ ),
    .Y(\reg_module/_08615_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16166_  (.A1(\reg_module/_08613_ ),
    .A2(\reg_module/_08615_ ),
    .B1(\reg_module/_08612_ ),
    .Y(\reg_module/_00215_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16167_  (.A(\reg_module/_08522_ ),
    .X(\reg_module/_08616_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16168_  (.A(\reg_module/_08616_ ),
    .B(net1556),
    .Y(\reg_module/_08617_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16169_  (.A(\reg_module/_08573_ ),
    .X(\reg_module/_08618_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16170_  (.A(\reg_module/_08618_ ),
    .B(net985),
    .C(\reg_module/_07966_ ),
    .Y(\reg_module/_08619_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16171_  (.A(\reg_module/_08609_ ),
    .B(\reg_module/_08619_ ),
    .Y(\reg_module/_08620_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16172_  (.A1(\reg_module/_08617_ ),
    .A2(\reg_module/_08620_ ),
    .B1(\reg_module/_08612_ ),
    .Y(\reg_module/_00216_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16173_  (.A(\reg_module/_08616_ ),
    .B(net1373),
    .Y(\reg_module/_08621_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16174_  (.A(\reg_module/_08618_ ),
    .B(net985),
    .C(\reg_module/_07971_ ),
    .Y(\reg_module/_08622_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16175_  (.A(\reg_module/_08609_ ),
    .B(\reg_module/_08622_ ),
    .Y(\reg_module/_08623_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16176_  (.A1(\reg_module/_08621_ ),
    .A2(\reg_module/_08623_ ),
    .B1(\reg_module/_08612_ ),
    .Y(\reg_module/_00217_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16177_  (.A(\reg_module/_08616_ ),
    .B(net1503),
    .Y(\reg_module/_08624_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16178_  (.A(\reg_module/_08618_ ),
    .B(net979),
    .C(\reg_module/_07976_ ),
    .Y(\reg_module/_08625_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16179_  (.A(\reg_module/_08609_ ),
    .B(\reg_module/_08625_ ),
    .Y(\reg_module/_08626_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16180_  (.A1(\reg_module/_08624_ ),
    .A2(\reg_module/_08626_ ),
    .B1(\reg_module/_08612_ ),
    .Y(\reg_module/_00218_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16181_  (.A(\reg_module/_08616_ ),
    .B(net1666),
    .Y(\reg_module/_08627_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16182_  (.A(\reg_module/_08618_ ),
    .B(net979),
    .C(\reg_module/_07981_ ),
    .Y(\reg_module/_08628_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16183_  (.A(\reg_module/_08609_ ),
    .B(\reg_module/_08628_ ),
    .Y(\reg_module/_08629_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16184_  (.A1(\reg_module/_08627_ ),
    .A2(\reg_module/_08629_ ),
    .B1(\reg_module/_08612_ ),
    .Y(\reg_module/_00219_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16185_  (.A(\reg_module/_08616_ ),
    .B(net1400),
    .Y(\reg_module/_08630_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16186_  (.A(\reg_module/_08540_ ),
    .X(\reg_module/_08631_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16187_  (.A(\reg_module/_08618_ ),
    .B(net976),
    .C(\reg_module/_07989_ ),
    .Y(\reg_module/_08632_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16188_  (.A(\reg_module/_08631_ ),
    .B(\reg_module/_08632_ ),
    .Y(\reg_module/_08633_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_16189_  (.A(\reg_module/_08544_ ),
    .X(\reg_module/_08634_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16190_  (.A1(\reg_module/_08630_ ),
    .A2(\reg_module/_08633_ ),
    .B1(\reg_module/_08634_ ),
    .Y(\reg_module/_00220_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16191_  (.A(\reg_module/_08616_ ),
    .B(net1368),
    .Y(\reg_module/_08635_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16192_  (.A(\reg_module/_08618_ ),
    .B(net977),
    .C(\reg_module/_07997_ ),
    .Y(\reg_module/_08636_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16193_  (.A(\reg_module/_08631_ ),
    .B(\reg_module/_08636_ ),
    .Y(\reg_module/_08637_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16194_  (.A1(\reg_module/_08635_ ),
    .A2(\reg_module/_08637_ ),
    .B1(\reg_module/_08634_ ),
    .Y(\reg_module/_00221_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16195_  (.A(\reg_module/_08523_ ),
    .B(net1385),
    .Y(\reg_module/_08638_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16196_  (.A(\reg_module/_07626_ ),
    .X(\reg_module/_08639_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16197_  (.A(\reg_module/_08639_ ),
    .B(net976),
    .C(\reg_module/_08003_ ),
    .Y(\reg_module/_08640_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16198_  (.A(\reg_module/_08631_ ),
    .B(\reg_module/_08640_ ),
    .Y(\reg_module/_08641_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16199_  (.A1(\reg_module/_08638_ ),
    .A2(\reg_module/_08641_ ),
    .B1(\reg_module/_08634_ ),
    .Y(\reg_module/_00222_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16200_  (.A(\reg_module/_08523_ ),
    .B(net1489),
    .Y(\reg_module/_08642_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_16201_  (.A(\reg_module/_08639_ ),
    .B(net976),
    .C(\reg_module/_08008_ ),
    .Y(\reg_module/_08643_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16202_  (.A(\reg_module/_08631_ ),
    .B(\reg_module/_08643_ ),
    .Y(\reg_module/_08644_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16203_  (.A1(\reg_module/_08642_ ),
    .A2(\reg_module/_08644_ ),
    .B1(\reg_module/_08634_ ),
    .Y(\reg_module/_00223_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16204_  (.A(net978),
    .B(\reg_module/_08012_ ),
    .Y(\reg_module/_08645_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16205_  (.A(\reg_module/_08645_ ),
    .B(net964),
    .Y(\reg_module/_08646_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16206_  (.A(\reg_module/_08646_ ),
    .Y(\reg_module/_08647_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16207_  (.A(\reg_module/_07638_ ),
    .B(\reg_module/_08647_ ),
    .Y(\reg_module/_08648_ ));
 sky130_fd_sc_hd__buf_8 \reg_module/_16208_  (.A(\reg_module/_08648_ ),
    .X(\reg_module/_08649_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16209_  (.A(\reg_module/_08649_ ),
    .X(\reg_module/_08650_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16210_  (.A(\reg_module/_08650_ ),
    .B(\reg_module/_04993_ ),
    .Y(\reg_module/_08651_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16211_  (.A(\reg_module/_08651_ ),
    .Y(\reg_module/_08652_ ));
 sky130_fd_sc_hd__buf_8 \reg_module/_16212_  (.A(\reg_module/_08647_ ),
    .X(\reg_module/_08653_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16213_  (.A(\reg_module/_08653_ ),
    .X(\reg_module/_08654_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16214_  (.A(\reg_module/_08340_ ),
    .B(\reg_module/_07514_ ),
    .C(\reg_module/_08654_ ),
    .Y(\reg_module/_08655_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16215_  (.A(\reg_module/_08655_ ),
    .B(net1032),
    .Y(\reg_module/_08656_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16216_  (.A(\reg_module/_08652_ ),
    .B(\reg_module/_08656_ ),
    .Y(\reg_module/_00224_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16217_  (.A(\reg_module/_08650_ ),
    .B(\reg_module/_05126_ ),
    .Y(\reg_module/_08657_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16218_  (.A(\reg_module/_08657_ ),
    .Y(\reg_module/_08658_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16219_  (.A(\reg_module/_08340_ ),
    .B(\reg_module/_07517_ ),
    .C(\reg_module/_08654_ ),
    .Y(\reg_module/_08659_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16220_  (.A(\reg_module/_08659_ ),
    .B(net1033),
    .Y(\reg_module/_08660_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16221_  (.A(\reg_module/_08658_ ),
    .B(\reg_module/_08660_ ),
    .Y(\reg_module/_00225_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16222_  (.A(\reg_module/_08650_ ),
    .B(\reg_module/_05206_ ),
    .Y(\reg_module/_08661_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16223_  (.A(\reg_module/_08661_ ),
    .Y(\reg_module/_08662_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16224_  (.A(\reg_module/_07639_ ),
    .X(\reg_module/_08663_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_16225_  (.A(\reg_module/_08663_ ),
    .X(\reg_module/_08664_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16226_  (.A(\reg_module/_08664_ ),
    .B(\reg_module/_07520_ ),
    .C(\reg_module/_08654_ ),
    .Y(\reg_module/_08665_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16227_  (.A(\reg_module/_08665_ ),
    .B(net1036),
    .Y(\reg_module/_08666_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16228_  (.A(\reg_module/_08662_ ),
    .B(\reg_module/_08666_ ),
    .Y(\reg_module/_00226_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16229_  (.A(\reg_module/gprf[227] ),
    .Y(\reg_module/_08667_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16230_  (.A(\reg_module/_08650_ ),
    .B(\reg_module/_08667_ ),
    .Y(\reg_module/_08668_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16231_  (.A(\reg_module/_08668_ ),
    .Y(\reg_module/_08669_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16232_  (.A(\reg_module/_08664_ ),
    .B(\reg_module/_07523_ ),
    .C(\reg_module/_08654_ ),
    .Y(\reg_module/_08670_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16233_  (.A(\reg_module/_08670_ ),
    .B(net1035),
    .Y(\reg_module/_08671_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16234_  (.A(\reg_module/_08669_ ),
    .B(\reg_module/_08671_ ),
    .Y(\reg_module/_00227_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16235_  (.A(\reg_module/gprf[228] ),
    .Y(\reg_module/_08672_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16236_  (.A(\reg_module/_08650_ ),
    .B(\reg_module/_08672_ ),
    .Y(\reg_module/_08673_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16237_  (.A(\reg_module/_08673_ ),
    .Y(\reg_module/_08674_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16238_  (.A(\reg_module/_08664_ ),
    .B(\reg_module/_07528_ ),
    .C(\reg_module/_08654_ ),
    .Y(\reg_module/_08675_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16239_  (.A(\reg_module/_08675_ ),
    .B(net1047),
    .Y(\reg_module/_08676_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16240_  (.A(\reg_module/_08674_ ),
    .B(\reg_module/_08676_ ),
    .Y(\reg_module/_00228_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16241_  (.A(\reg_module/gprf[229] ),
    .Y(\reg_module/_08677_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16242_  (.A(\reg_module/_08650_ ),
    .B(\reg_module/_08677_ ),
    .Y(\reg_module/_08678_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16243_  (.A(\reg_module/_08678_ ),
    .Y(\reg_module/_08679_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16244_  (.A(\reg_module/_08664_ ),
    .B(\reg_module/_07531_ ),
    .C(\reg_module/_08654_ ),
    .Y(\reg_module/_08680_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16245_  (.A(\reg_module/_08680_ ),
    .B(net1047),
    .Y(\reg_module/_08681_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16246_  (.A(\reg_module/_08679_ ),
    .B(\reg_module/_08681_ ),
    .Y(\reg_module/_00229_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16247_  (.A(\reg_module/_08649_ ),
    .X(\reg_module/_08682_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16248_  (.A(\reg_module/gprf[230] ),
    .Y(\reg_module/_08683_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16249_  (.A(\reg_module/_08682_ ),
    .B(\reg_module/_08683_ ),
    .Y(\reg_module/_08684_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16250_  (.A(\reg_module/_08684_ ),
    .Y(\reg_module/_08685_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16251_  (.A(\reg_module/_08653_ ),
    .X(\reg_module/_08686_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16252_  (.A(\reg_module/_08664_ ),
    .B(\reg_module/_07535_ ),
    .C(\reg_module/_08686_ ),
    .Y(\reg_module/_08687_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16253_  (.A(\reg_module/_08687_ ),
    .B(net1051),
    .Y(\reg_module/_08688_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16254_  (.A(\reg_module/_08685_ ),
    .B(\reg_module/_08688_ ),
    .Y(\reg_module/_00230_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16255_  (.A(net2157),
    .Y(\reg_module/_08689_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16256_  (.A(\reg_module/_08682_ ),
    .B(\reg_module/_08689_ ),
    .Y(\reg_module/_08690_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16257_  (.A(\reg_module/_08690_ ),
    .Y(\reg_module/_08691_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16258_  (.A(\reg_module/_08664_ ),
    .B(\reg_module/_07538_ ),
    .C(\reg_module/_08686_ ),
    .Y(\reg_module/_08692_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16259_  (.A(\reg_module/_08692_ ),
    .B(net1050),
    .Y(\reg_module/_08693_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16260_  (.A(\reg_module/_08691_ ),
    .B(\reg_module/_08693_ ),
    .Y(\reg_module/_00231_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16261_  (.A(net2220),
    .Y(\reg_module/_08694_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16262_  (.A(\reg_module/_08682_ ),
    .B(\reg_module/_08694_ ),
    .Y(\reg_module/_08695_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16263_  (.A(\reg_module/_08695_ ),
    .Y(\reg_module/_08696_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16264_  (.A(\reg_module/_08663_ ),
    .X(\reg_module/_08697_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16265_  (.A(\reg_module/_08697_ ),
    .B(\reg_module/_07541_ ),
    .C(\reg_module/_08686_ ),
    .Y(\reg_module/_08698_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16266_  (.A(\reg_module/_08698_ ),
    .B(net1048),
    .Y(\reg_module/_08699_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16267_  (.A(\reg_module/_08696_ ),
    .B(\reg_module/_08699_ ),
    .Y(\reg_module/_00232_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16268_  (.A(net2219),
    .Y(\reg_module/_08700_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16269_  (.A(\reg_module/_08682_ ),
    .B(\reg_module/_08700_ ),
    .Y(\reg_module/_08701_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16270_  (.A(\reg_module/_08701_ ),
    .Y(\reg_module/_08702_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16271_  (.A(\reg_module/_08697_ ),
    .B(\reg_module/_07544_ ),
    .C(\reg_module/_08686_ ),
    .Y(\reg_module/_08703_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16272_  (.A(\reg_module/_08703_ ),
    .B(net1049),
    .Y(\reg_module/_08704_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16273_  (.A(\reg_module/_08702_ ),
    .B(\reg_module/_08704_ ),
    .Y(\reg_module/_00233_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16274_  (.A(\reg_module/gprf[234] ),
    .Y(\reg_module/_08705_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16275_  (.A(\reg_module/_08682_ ),
    .B(\reg_module/_08705_ ),
    .Y(\reg_module/_08706_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16276_  (.A(\reg_module/_08706_ ),
    .Y(\reg_module/_08707_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16277_  (.A(\reg_module/_08697_ ),
    .B(\reg_module/_07548_ ),
    .C(\reg_module/_08686_ ),
    .Y(\reg_module/_08708_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16278_  (.A(\reg_module/_08708_ ),
    .B(net1049),
    .Y(\reg_module/_08709_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16279_  (.A(\reg_module/_08707_ ),
    .B(\reg_module/_08709_ ),
    .Y(\reg_module/_00234_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16280_  (.A(\reg_module/gprf[235] ),
    .Y(\reg_module/_08710_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16281_  (.A(\reg_module/_08682_ ),
    .B(\reg_module/_08710_ ),
    .Y(\reg_module/_08711_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16282_  (.A(\reg_module/_08711_ ),
    .Y(\reg_module/_08712_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16283_  (.A(\reg_module/_08697_ ),
    .B(\reg_module/_07551_ ),
    .C(\reg_module/_08686_ ),
    .Y(\reg_module/_08713_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16284_  (.A(\reg_module/_08713_ ),
    .B(net1049),
    .Y(\reg_module/_08714_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16285_  (.A(\reg_module/_08712_ ),
    .B(\reg_module/_08714_ ),
    .Y(\reg_module/_00235_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16286_  (.A(\reg_module/_08649_ ),
    .X(\reg_module/_08715_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16287_  (.A(\reg_module/gprf[236] ),
    .Y(\reg_module/_08716_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16288_  (.A(\reg_module/_08715_ ),
    .B(\reg_module/_08716_ ),
    .Y(\reg_module/_08717_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16289_  (.A(\reg_module/_08717_ ),
    .Y(\reg_module/_08718_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_16290_  (.A(\reg_module/_08653_ ),
    .X(\reg_module/_08719_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16291_  (.A(\reg_module/_08697_ ),
    .B(\reg_module/_07555_ ),
    .C(\reg_module/_08719_ ),
    .Y(\reg_module/_08720_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16292_  (.A(\reg_module/_08720_ ),
    .B(net1063),
    .Y(\reg_module/_08721_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16293_  (.A(\reg_module/_08718_ ),
    .B(\reg_module/_08721_ ),
    .Y(\reg_module/_00236_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16294_  (.A(net2216),
    .Y(\reg_module/_08722_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16295_  (.A(\reg_module/_08715_ ),
    .B(\reg_module/_08722_ ),
    .Y(\reg_module/_08723_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16296_  (.A(\reg_module/_08723_ ),
    .Y(\reg_module/_08724_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16297_  (.A(\reg_module/_08697_ ),
    .B(\reg_module/_07558_ ),
    .C(\reg_module/_08719_ ),
    .Y(\reg_module/_08725_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16298_  (.A(\reg_module/_08725_ ),
    .B(net1063),
    .Y(\reg_module/_08726_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16299_  (.A(\reg_module/_08724_ ),
    .B(\reg_module/_08726_ ),
    .Y(\reg_module/_00237_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16300_  (.A(net2210),
    .Y(\reg_module/_08727_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16301_  (.A(\reg_module/_08715_ ),
    .B(\reg_module/_08727_ ),
    .Y(\reg_module/_08728_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16302_  (.A(\reg_module/_08728_ ),
    .Y(\reg_module/_08729_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_16303_  (.A(\reg_module/_08663_ ),
    .X(\reg_module/_08730_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16304_  (.A(\reg_module/_08730_ ),
    .B(\reg_module/_07561_ ),
    .C(\reg_module/_08719_ ),
    .Y(\reg_module/_08731_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16305_  (.A(\reg_module/_08731_ ),
    .B(net1063),
    .Y(\reg_module/_08732_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16306_  (.A(\reg_module/_08729_ ),
    .B(\reg_module/_08732_ ),
    .Y(\reg_module/_00238_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16307_  (.A(\reg_module/gprf[239] ),
    .Y(\reg_module/_08733_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16308_  (.A(\reg_module/_08715_ ),
    .B(\reg_module/_08733_ ),
    .Y(\reg_module/_08734_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16309_  (.A(\reg_module/_08734_ ),
    .Y(\reg_module/_08735_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16310_  (.A(\reg_module/_08730_ ),
    .B(\reg_module/_07564_ ),
    .C(\reg_module/_08719_ ),
    .Y(\reg_module/_08736_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16311_  (.A(\reg_module/_08736_ ),
    .B(net1063),
    .Y(\reg_module/_08737_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16312_  (.A(\reg_module/_08735_ ),
    .B(\reg_module/_08737_ ),
    .Y(\reg_module/_00239_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16313_  (.A(net2215),
    .Y(\reg_module/_08738_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16314_  (.A(\reg_module/_08715_ ),
    .B(\reg_module/_08738_ ),
    .Y(\reg_module/_08739_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16315_  (.A(\reg_module/_08739_ ),
    .Y(\reg_module/_08740_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16316_  (.A(\reg_module/_08730_ ),
    .B(\reg_module/_07568_ ),
    .C(\reg_module/_08719_ ),
    .Y(\reg_module/_08741_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16317_  (.A(\reg_module/_08741_ ),
    .B(net1055),
    .Y(\reg_module/_08742_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16318_  (.A(\reg_module/_08740_ ),
    .B(\reg_module/_08742_ ),
    .Y(\reg_module/_00240_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16319_  (.A(net2224),
    .Y(\reg_module/_08743_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16320_  (.A(\reg_module/_08715_ ),
    .B(\reg_module/_08743_ ),
    .Y(\reg_module/_08744_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16321_  (.A(\reg_module/_08744_ ),
    .Y(\reg_module/_08745_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16322_  (.A(\reg_module/_08730_ ),
    .B(\reg_module/_07571_ ),
    .C(\reg_module/_08719_ ),
    .Y(\reg_module/_08746_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16323_  (.A(\reg_module/_08746_ ),
    .B(net1055),
    .Y(\reg_module/_08747_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16324_  (.A(\reg_module/_08745_ ),
    .B(\reg_module/_08747_ ),
    .Y(\reg_module/_00241_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16325_  (.A(\reg_module/_08649_ ),
    .X(\reg_module/_08748_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16326_  (.A(\reg_module/gprf[242] ),
    .Y(\reg_module/_08749_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16327_  (.A(\reg_module/_08748_ ),
    .B(\reg_module/_08749_ ),
    .Y(\reg_module/_08750_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16328_  (.A(\reg_module/_08750_ ),
    .Y(\reg_module/_08751_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16329_  (.A(\reg_module/_08653_ ),
    .X(\reg_module/_08752_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16330_  (.A(\reg_module/_08730_ ),
    .B(\reg_module/_07575_ ),
    .C(\reg_module/_08752_ ),
    .Y(\reg_module/_08753_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16331_  (.A(\reg_module/_08753_ ),
    .B(net1040),
    .Y(\reg_module/_08754_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16332_  (.A(\reg_module/_08751_ ),
    .B(\reg_module/_08754_ ),
    .Y(\reg_module/_00242_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16333_  (.A(net2162),
    .Y(\reg_module/_08755_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16334_  (.A(\reg_module/_08748_ ),
    .B(\reg_module/_08755_ ),
    .Y(\reg_module/_08756_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16335_  (.A(\reg_module/_08756_ ),
    .Y(\reg_module/_08757_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16336_  (.A(\reg_module/_08730_ ),
    .B(\reg_module/_07578_ ),
    .C(\reg_module/_08752_ ),
    .Y(\reg_module/_08758_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16337_  (.A(\reg_module/_08758_ ),
    .B(net1040),
    .Y(\reg_module/_08759_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16338_  (.A(\reg_module/_08757_ ),
    .B(\reg_module/_08759_ ),
    .Y(\reg_module/_00243_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16339_  (.A(\reg_module/gprf[244] ),
    .Y(\reg_module/_08760_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16340_  (.A(\reg_module/_08748_ ),
    .B(\reg_module/_08760_ ),
    .Y(\reg_module/_08761_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16341_  (.A(\reg_module/_08761_ ),
    .Y(\reg_module/_08762_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16342_  (.A(\reg_module/_08663_ ),
    .X(\reg_module/_08763_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16343_  (.A(\reg_module/_08763_ ),
    .B(\reg_module/_07581_ ),
    .C(\reg_module/_08752_ ),
    .Y(\reg_module/_08764_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16344_  (.A(\reg_module/_08764_ ),
    .B(net1040),
    .Y(\reg_module/_08765_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16345_  (.A(\reg_module/_08762_ ),
    .B(\reg_module/_08765_ ),
    .Y(\reg_module/_00244_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16346_  (.A(net2150),
    .Y(\reg_module/_08766_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16347_  (.A(\reg_module/_08748_ ),
    .B(\reg_module/_08766_ ),
    .Y(\reg_module/_08767_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16348_  (.A(\reg_module/_08767_ ),
    .Y(\reg_module/_08768_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16349_  (.A(\reg_module/_08763_ ),
    .B(\reg_module/_07584_ ),
    .C(\reg_module/_08752_ ),
    .Y(\reg_module/_08769_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16350_  (.A(\reg_module/_08769_ ),
    .B(net1040),
    .Y(\reg_module/_08770_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16351_  (.A(\reg_module/_08768_ ),
    .B(\reg_module/_08770_ ),
    .Y(\reg_module/_00245_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16352_  (.A(net2201),
    .Y(\reg_module/_08771_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16353_  (.A(\reg_module/_08748_ ),
    .B(\reg_module/_08771_ ),
    .Y(\reg_module/_08772_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16354_  (.A(\reg_module/_08772_ ),
    .Y(\reg_module/_08773_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16355_  (.A(\reg_module/_08763_ ),
    .B(\reg_module/_07588_ ),
    .C(\reg_module/_08752_ ),
    .Y(\reg_module/_08774_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16356_  (.A(\reg_module/_08774_ ),
    .B(net1040),
    .Y(\reg_module/_08775_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16357_  (.A(\reg_module/_08773_ ),
    .B(\reg_module/_08775_ ),
    .Y(\reg_module/_00246_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16358_  (.A(net2196),
    .Y(\reg_module/_08776_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16359_  (.A(\reg_module/_08748_ ),
    .B(\reg_module/_08776_ ),
    .Y(\reg_module/_08777_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16360_  (.A(\reg_module/_08777_ ),
    .Y(\reg_module/_08778_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16361_  (.A(\reg_module/_08763_ ),
    .B(\reg_module/_07591_ ),
    .C(\reg_module/_08752_ ),
    .Y(\reg_module/_08779_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16362_  (.A(\reg_module/_08779_ ),
    .B(net1038),
    .Y(\reg_module/_08780_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16363_  (.A(\reg_module/_08778_ ),
    .B(\reg_module/_08780_ ),
    .Y(\reg_module/_00247_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16364_  (.A(\reg_module/_08648_ ),
    .X(\reg_module/_08781_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16365_  (.A(net2185),
    .Y(\reg_module/_08782_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16366_  (.A(\reg_module/_08781_ ),
    .B(\reg_module/_08782_ ),
    .Y(\reg_module/_08783_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16367_  (.A(\reg_module/_08783_ ),
    .Y(\reg_module/_08784_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16368_  (.A(\reg_module/_08647_ ),
    .X(\reg_module/_08785_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16369_  (.A(\reg_module/_08763_ ),
    .B(\reg_module/_07595_ ),
    .C(\reg_module/_08785_ ),
    .Y(\reg_module/_08786_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16370_  (.A(\reg_module/_08786_ ),
    .B(net1006),
    .Y(\reg_module/_08787_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16371_  (.A(\reg_module/_08784_ ),
    .B(\reg_module/_08787_ ),
    .Y(\reg_module/_00248_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16372_  (.A(net2166),
    .Y(\reg_module/_08788_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16373_  (.A(\reg_module/_08781_ ),
    .B(\reg_module/_08788_ ),
    .Y(\reg_module/_08789_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16374_  (.A(\reg_module/_08789_ ),
    .Y(\reg_module/_08790_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16375_  (.A(\reg_module/_08763_ ),
    .B(\reg_module/_07598_ ),
    .C(\reg_module/_08785_ ),
    .Y(\reg_module/_08791_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16376_  (.A(\reg_module/_08791_ ),
    .B(net1006),
    .Y(\reg_module/_08792_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16377_  (.A(\reg_module/_08790_ ),
    .B(\reg_module/_08792_ ),
    .Y(\reg_module/_00249_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16378_  (.A(net2183),
    .Y(\reg_module/_08793_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16379_  (.A(\reg_module/_08781_ ),
    .B(\reg_module/_08793_ ),
    .Y(\reg_module/_08794_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16380_  (.A(\reg_module/_08794_ ),
    .Y(\reg_module/_08795_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16381_  (.A(\reg_module/_08663_ ),
    .X(\reg_module/_08796_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16382_  (.A(\reg_module/_08796_ ),
    .B(\reg_module/_07601_ ),
    .C(\reg_module/_08785_ ),
    .Y(\reg_module/_08797_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16383_  (.A(\reg_module/_08797_ ),
    .B(net1005),
    .Y(\reg_module/_08798_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16384_  (.A(\reg_module/_08795_ ),
    .B(\reg_module/_08798_ ),
    .Y(\reg_module/_00250_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16385_  (.A(net2171),
    .Y(\reg_module/_08799_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16386_  (.A(\reg_module/_08781_ ),
    .B(\reg_module/_08799_ ),
    .Y(\reg_module/_08800_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16387_  (.A(\reg_module/_08800_ ),
    .Y(\reg_module/_08801_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16388_  (.A(\reg_module/_08796_ ),
    .B(\reg_module/_07604_ ),
    .C(\reg_module/_08785_ ),
    .Y(\reg_module/_08802_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16389_  (.A(\reg_module/_08802_ ),
    .B(net1005),
    .Y(\reg_module/_08803_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16390_  (.A(\reg_module/_08801_ ),
    .B(\reg_module/_08803_ ),
    .Y(\reg_module/_00251_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16391_  (.A(\reg_module/gprf[252] ),
    .Y(\reg_module/_08804_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16392_  (.A(\reg_module/_08781_ ),
    .B(\reg_module/_08804_ ),
    .Y(\reg_module/_08805_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16393_  (.A(\reg_module/_08805_ ),
    .Y(\reg_module/_08806_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16394_  (.A(\reg_module/_08796_ ),
    .B(\reg_module/_07607_ ),
    .C(\reg_module/_08785_ ),
    .Y(\reg_module/_08807_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16395_  (.A(\reg_module/_08807_ ),
    .B(net1009),
    .Y(\reg_module/_08808_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16396_  (.A(\reg_module/_08806_ ),
    .B(\reg_module/_08808_ ),
    .Y(\reg_module/_00252_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16397_  (.A(net2172),
    .Y(\reg_module/_08809_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16398_  (.A(\reg_module/_08781_ ),
    .B(\reg_module/_08809_ ),
    .Y(\reg_module/_08810_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16399_  (.A(\reg_module/_08810_ ),
    .Y(\reg_module/_08811_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16400_  (.A(\reg_module/_08796_ ),
    .B(\reg_module/_07610_ ),
    .C(\reg_module/_08785_ ),
    .Y(\reg_module/_08812_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16401_  (.A(\reg_module/_08812_ ),
    .B(net1009),
    .Y(\reg_module/_08813_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16402_  (.A(\reg_module/_08811_ ),
    .B(\reg_module/_08813_ ),
    .Y(\reg_module/_00253_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16403_  (.A(net2154),
    .Y(\reg_module/_08814_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16404_  (.A(\reg_module/_08649_ ),
    .B(\reg_module/_08814_ ),
    .Y(\reg_module/_08815_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16405_  (.A(\reg_module/_08815_ ),
    .Y(\reg_module/_08816_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16406_  (.A(\reg_module/_08796_ ),
    .B(\reg_module/_07613_ ),
    .C(\reg_module/_08653_ ),
    .Y(\reg_module/_08817_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16407_  (.A(\reg_module/_08817_ ),
    .B(net1010),
    .Y(\reg_module/_08818_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16408_  (.A(\reg_module/_08816_ ),
    .B(\reg_module/_08818_ ),
    .Y(\reg_module/_00254_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16409_  (.A(net2225),
    .Y(\reg_module/_08819_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16410_  (.A(\reg_module/_08649_ ),
    .B(\reg_module/_08819_ ),
    .Y(\reg_module/_08820_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16411_  (.A(\reg_module/_08820_ ),
    .Y(\reg_module/_08821_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16412_  (.A(\reg_module/_08796_ ),
    .B(\reg_module/_07616_ ),
    .C(\reg_module/_08653_ ),
    .Y(\reg_module/_08822_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16413_  (.A(\reg_module/_08822_ ),
    .B(net1010),
    .Y(\reg_module/_08823_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16414_  (.A(\reg_module/_08821_ ),
    .B(\reg_module/_08823_ ),
    .Y(\reg_module/_00255_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16415_  (.A(\reg_module/_07508_ ),
    .Y(\reg_module/_08824_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16416_  (.A(\reg_module/_07623_ ),
    .X(\reg_module/_08825_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_16417_  (.A(net963),
    .B(\reg_module/_07499_ ),
    .Y(\reg_module/_08826_ ));
 sky130_fd_sc_hd__nand3_2 \reg_module/_16418_  (.A(\reg_module/_08824_ ),
    .B(\reg_module/_08825_ ),
    .C(\reg_module/_08826_ ),
    .Y(\reg_module/_08827_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16419_  (.A(\reg_module/_08827_ ),
    .X(\reg_module/_08828_ ));
 sky130_fd_sc_hd__inv_6 \reg_module/_16420_  (.A(\reg_module/_08828_ ),
    .Y(\reg_module/_08829_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16421_  (.A(\reg_module/_08827_ ),
    .X(\reg_module/_08830_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16422_  (.A(net2188),
    .Y(\reg_module/_08831_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16423_  (.A(\reg_module/_08830_ ),
    .B(\reg_module/_08831_ ),
    .Y(\reg_module/_08832_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16424_  (.A(\reg_module/_08832_ ),
    .B(net1038),
    .Y(\reg_module/_08833_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16425_  (.A1(\reg_module/_08829_ ),
    .A2(\reg_module/_07514_ ),
    .B1(\reg_module/_08833_ ),
    .Y(\reg_module/_00256_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16426_  (.A(\reg_module/_08828_ ),
    .X(\reg_module/_08834_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16427_  (.A(\reg_module/_08834_ ),
    .B(net1822),
    .Y(\reg_module/_08835_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16428_  (.A(\reg_module/_08826_ ),
    .Y(\reg_module/_08836_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16429_  (.A(\reg_module/_08836_ ),
    .X(\reg_module/_08837_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16430_  (.A(\reg_module/_08837_ ),
    .X(\reg_module/_08838_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16431_  (.A(\reg_module/_07516_ ),
    .B(\reg_module/_08838_ ),
    .Y(\reg_module/_08839_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16432_  (.A(\reg_module/_08631_ ),
    .B(\reg_module/_08839_ ),
    .Y(\reg_module/_08840_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16433_  (.A1(\reg_module/_08835_ ),
    .A2(\reg_module/_08840_ ),
    .B1(\reg_module/_08634_ ),
    .Y(\reg_module/_00257_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16434_  (.A(\reg_module/_08834_ ),
    .B(net1578),
    .Y(\reg_module/_08841_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16435_  (.A(\reg_module/_07519_ ),
    .B(\reg_module/_08838_ ),
    .Y(\reg_module/_08842_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16436_  (.A(\reg_module/_08631_ ),
    .B(\reg_module/_08842_ ),
    .Y(\reg_module/_08843_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16437_  (.A1(\reg_module/_08841_ ),
    .A2(\reg_module/_08843_ ),
    .B1(\reg_module/_08634_ ),
    .Y(\reg_module/_00258_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16438_  (.A(net2169),
    .Y(\reg_module/_08844_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16439_  (.A(\reg_module/_08830_ ),
    .B(\reg_module/_08844_ ),
    .Y(\reg_module/_08845_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16440_  (.A(\reg_module/_08845_ ),
    .B(net1042),
    .Y(\reg_module/_08846_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16441_  (.A1(\reg_module/_08829_ ),
    .A2(\reg_module/_07523_ ),
    .B1(\reg_module/_08846_ ),
    .Y(\reg_module/_00259_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16442_  (.A(\reg_module/_08834_ ),
    .B(net1471),
    .Y(\reg_module/_08847_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16443_  (.A(\reg_module/_08540_ ),
    .X(\reg_module/_08848_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16444_  (.A(\reg_module/_07527_ ),
    .B(\reg_module/_08838_ ),
    .Y(\reg_module/_08849_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16445_  (.A(\reg_module/_08848_ ),
    .B(\reg_module/_08849_ ),
    .Y(\reg_module/_08850_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16446_  (.A(\reg_module/_08544_ ),
    .X(\reg_module/_08851_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16447_  (.A1(\reg_module/_08847_ ),
    .A2(\reg_module/_08850_ ),
    .B1(\reg_module/_08851_ ),
    .Y(\reg_module/_00260_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16448_  (.A(\reg_module/_08834_ ),
    .B(net1464),
    .Y(\reg_module/_08852_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16449_  (.A(\reg_module/_07530_ ),
    .B(\reg_module/_08838_ ),
    .Y(\reg_module/_08853_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16450_  (.A(\reg_module/_08848_ ),
    .B(\reg_module/_08853_ ),
    .Y(\reg_module/_08854_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16451_  (.A1(\reg_module/_08852_ ),
    .A2(\reg_module/_08854_ ),
    .B1(\reg_module/_08851_ ),
    .Y(\reg_module/_00261_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16452_  (.A(\reg_module/_08834_ ),
    .B(net1494),
    .Y(\reg_module/_08855_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16453_  (.A(\reg_module/_07534_ ),
    .B(\reg_module/_08838_ ),
    .Y(\reg_module/_08856_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16454_  (.A(\reg_module/_08848_ ),
    .B(\reg_module/_08856_ ),
    .Y(\reg_module/_08857_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16455_  (.A1(\reg_module/_08855_ ),
    .A2(\reg_module/_08857_ ),
    .B1(\reg_module/_08851_ ),
    .Y(\reg_module/_00262_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16456_  (.A(\reg_module/_08834_ ),
    .B(net1747),
    .Y(\reg_module/_08858_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16457_  (.A(\reg_module/_07537_ ),
    .B(\reg_module/_08838_ ),
    .Y(\reg_module/_08859_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16458_  (.A(\reg_module/_08848_ ),
    .B(\reg_module/_08859_ ),
    .Y(\reg_module/_08860_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16459_  (.A1(\reg_module/_08858_ ),
    .A2(\reg_module/_08860_ ),
    .B1(\reg_module/_08851_ ),
    .Y(\reg_module/_00263_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_16460_  (.A(\reg_module/_08828_ ),
    .X(\reg_module/_08861_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16461_  (.A(\reg_module/_08861_ ),
    .B(net1607),
    .Y(\reg_module/_08862_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_16462_  (.A(\reg_module/_08837_ ),
    .X(\reg_module/_08863_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16463_  (.A(\reg_module/_07540_ ),
    .B(\reg_module/_08863_ ),
    .Y(\reg_module/_08864_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16464_  (.A(\reg_module/_08848_ ),
    .B(\reg_module/_08864_ ),
    .Y(\reg_module/_08865_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16465_  (.A1(\reg_module/_08862_ ),
    .A2(\reg_module/_08865_ ),
    .B1(\reg_module/_08851_ ),
    .Y(\reg_module/_00264_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16466_  (.A(\reg_module/_08861_ ),
    .B(net1829),
    .Y(\reg_module/_08866_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16467_  (.A(\reg_module/_07543_ ),
    .B(\reg_module/_08863_ ),
    .Y(\reg_module/_08867_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16468_  (.A(\reg_module/_08848_ ),
    .B(\reg_module/_08867_ ),
    .Y(\reg_module/_08868_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16469_  (.A1(\reg_module/_08866_ ),
    .A2(\reg_module/_08868_ ),
    .B1(\reg_module/_08851_ ),
    .Y(\reg_module/_00265_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16470_  (.A(\reg_module/gprf[266] ),
    .Y(\reg_module/_08869_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16471_  (.A(\reg_module/_08830_ ),
    .B(\reg_module/_08869_ ),
    .Y(\reg_module/_08870_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16472_  (.A(\reg_module/_08870_ ),
    .B(net1066),
    .Y(\reg_module/_08871_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16473_  (.A1(\reg_module/_08829_ ),
    .A2(\reg_module/_07548_ ),
    .B1(\reg_module/_08871_ ),
    .Y(\reg_module/_00266_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16474_  (.A(\reg_module/_08861_ ),
    .B(net2114),
    .Y(\reg_module/_08872_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16475_  (.A(\reg_module/_08183_ ),
    .X(\reg_module/_08873_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16476_  (.A(\reg_module/_08873_ ),
    .X(\reg_module/_08874_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_16477_  (.A(\reg_module/_07550_ ),
    .B(\reg_module/_08863_ ),
    .Y(\reg_module/_08875_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16478_  (.A(\reg_module/_08874_ ),
    .B(\reg_module/_08875_ ),
    .Y(\reg_module/_08876_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_16479_  (.A(\reg_module/_07993_ ),
    .X(\reg_module/_08877_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16480_  (.A(\reg_module/_08877_ ),
    .X(\reg_module/_08878_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16481_  (.A1(\reg_module/_08872_ ),
    .A2(\reg_module/_08876_ ),
    .B1(\reg_module/_08878_ ),
    .Y(\reg_module/_00267_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16482_  (.A(\reg_module/_08861_ ),
    .B(net1534),
    .Y(\reg_module/_08879_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16483_  (.A(\reg_module/_07554_ ),
    .B(\reg_module/_08863_ ),
    .Y(\reg_module/_08880_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16484_  (.A(\reg_module/_08874_ ),
    .B(\reg_module/_08880_ ),
    .Y(\reg_module/_08881_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16485_  (.A1(\reg_module/_08879_ ),
    .A2(\reg_module/_08881_ ),
    .B1(\reg_module/_08878_ ),
    .Y(\reg_module/_00268_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16486_  (.A(net2222),
    .Y(\reg_module/_08882_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16487_  (.A(\reg_module/_08830_ ),
    .B(\reg_module/_08882_ ),
    .Y(\reg_module/_08883_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16488_  (.A(\reg_module/_08883_ ),
    .B(net1066),
    .Y(\reg_module/_08884_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16489_  (.A1(\reg_module/_08829_ ),
    .A2(\reg_module/_07558_ ),
    .B1(\reg_module/_08884_ ),
    .Y(\reg_module/_00269_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16490_  (.A(\reg_module/_08861_ ),
    .B(net1550),
    .Y(\reg_module/_08885_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16491_  (.A(\reg_module/_07560_ ),
    .B(\reg_module/_08863_ ),
    .Y(\reg_module/_08886_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16492_  (.A(\reg_module/_08874_ ),
    .B(\reg_module/_08886_ ),
    .Y(\reg_module/_08887_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16493_  (.A1(\reg_module/_08885_ ),
    .A2(\reg_module/_08887_ ),
    .B1(\reg_module/_08878_ ),
    .Y(\reg_module/_00270_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16494_  (.A(\reg_module/_08861_ ),
    .B(net1387),
    .Y(\reg_module/_08888_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16495_  (.A(\reg_module/_07563_ ),
    .B(\reg_module/_08863_ ),
    .Y(\reg_module/_08889_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16496_  (.A(\reg_module/_08874_ ),
    .B(\reg_module/_08889_ ),
    .Y(\reg_module/_08890_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16497_  (.A1(\reg_module/_08888_ ),
    .A2(\reg_module/_08890_ ),
    .B1(\reg_module/_08878_ ),
    .Y(\reg_module/_00271_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16498_  (.A(\reg_module/_08828_ ),
    .X(\reg_module/_08891_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16499_  (.A(\reg_module/_08891_ ),
    .B(net1498),
    .Y(\reg_module/_08892_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_16500_  (.A(\reg_module/_08837_ ),
    .X(\reg_module/_08893_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16501_  (.A(\reg_module/_07567_ ),
    .B(\reg_module/_08893_ ),
    .Y(\reg_module/_08894_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16502_  (.A(\reg_module/_08874_ ),
    .B(\reg_module/_08894_ ),
    .Y(\reg_module/_08895_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16503_  (.A1(\reg_module/_08892_ ),
    .A2(\reg_module/_08895_ ),
    .B1(\reg_module/_08878_ ),
    .Y(\reg_module/_00272_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16504_  (.A(\reg_module/_08891_ ),
    .B(net1645),
    .Y(\reg_module/_08896_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16505_  (.A(\reg_module/_07570_ ),
    .B(\reg_module/_08893_ ),
    .Y(\reg_module/_08897_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16506_  (.A(\reg_module/_08874_ ),
    .B(\reg_module/_08897_ ),
    .Y(\reg_module/_08898_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16507_  (.A1(\reg_module/_08896_ ),
    .A2(\reg_module/_08898_ ),
    .B1(\reg_module/_08878_ ),
    .Y(\reg_module/_00273_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16508_  (.A(net2167),
    .Y(\reg_module/_08899_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16509_  (.A(\reg_module/_08828_ ),
    .B(\reg_module/_08899_ ),
    .Y(\reg_module/_08900_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16510_  (.A(\reg_module/_08900_ ),
    .B(net1060),
    .Y(\reg_module/_08901_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16511_  (.A1(\reg_module/_08829_ ),
    .A2(\reg_module/_07575_ ),
    .B1(\reg_module/_08901_ ),
    .Y(\reg_module/_00274_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16512_  (.A(\reg_module/_08891_ ),
    .B(net2158),
    .Y(\reg_module/_08902_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16513_  (.A(\reg_module/_08873_ ),
    .X(\reg_module/_08903_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_16514_  (.A(\reg_module/_07577_ ),
    .B(\reg_module/_08893_ ),
    .Y(\reg_module/_08904_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16515_  (.A(\reg_module/_08903_ ),
    .B(\reg_module/_08904_ ),
    .Y(\reg_module/_08905_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16516_  (.A(\reg_module/_08877_ ),
    .X(\reg_module/_08906_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16517_  (.A1(\reg_module/_08902_ ),
    .A2(\reg_module/_08905_ ),
    .B1(\reg_module/_08906_ ),
    .Y(\reg_module/_00275_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16518_  (.A(\reg_module/_08891_ ),
    .B(net1937),
    .Y(\reg_module/_08907_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16519_  (.A(\reg_module/_07580_ ),
    .B(\reg_module/_08893_ ),
    .Y(\reg_module/_08908_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16520_  (.A(\reg_module/_08903_ ),
    .B(\reg_module/_08908_ ),
    .Y(\reg_module/_08909_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16521_  (.A1(\reg_module/_08907_ ),
    .A2(\reg_module/_08909_ ),
    .B1(\reg_module/_08906_ ),
    .Y(\reg_module/_00276_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16522_  (.A(\reg_module/_08891_ ),
    .B(net1889),
    .Y(\reg_module/_08910_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16523_  (.A(\reg_module/_07583_ ),
    .B(\reg_module/_08893_ ),
    .Y(\reg_module/_08911_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16524_  (.A(\reg_module/_08903_ ),
    .B(\reg_module/_08911_ ),
    .Y(\reg_module/_08912_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16525_  (.A1(\reg_module/_08910_ ),
    .A2(\reg_module/_08912_ ),
    .B1(\reg_module/_08906_ ),
    .Y(\reg_module/_00277_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16526_  (.A(\reg_module/_08891_ ),
    .B(net1324),
    .Y(\reg_module/_08913_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16527_  (.A(\reg_module/_07587_ ),
    .B(\reg_module/_08893_ ),
    .Y(\reg_module/_08914_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16528_  (.A(\reg_module/_08903_ ),
    .B(\reg_module/_08914_ ),
    .Y(\reg_module/_08915_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16529_  (.A1(\reg_module/_08913_ ),
    .A2(\reg_module/_08915_ ),
    .B1(\reg_module/_08906_ ),
    .Y(\reg_module/_00278_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16530_  (.A(net2207),
    .Y(\reg_module/_08916_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16531_  (.A(\reg_module/_08828_ ),
    .B(\reg_module/_08916_ ),
    .Y(\reg_module/_08917_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16532_  (.A(\reg_module/_08917_ ),
    .B(net1026),
    .Y(\reg_module/_08918_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16533_  (.A1(\reg_module/_08829_ ),
    .A2(\reg_module/_07591_ ),
    .B1(\reg_module/_08918_ ),
    .Y(\reg_module/_00279_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16534_  (.A(\reg_module/_08827_ ),
    .X(\reg_module/_08919_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16535_  (.A(\reg_module/_08919_ ),
    .B(net1265),
    .Y(\reg_module/_08920_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16536_  (.A(\reg_module/_08837_ ),
    .X(\reg_module/_08921_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16537_  (.A(\reg_module/_07594_ ),
    .B(\reg_module/_08921_ ),
    .Y(\reg_module/_08922_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16538_  (.A(\reg_module/_08903_ ),
    .B(\reg_module/_08922_ ),
    .Y(\reg_module/_08923_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16539_  (.A1(\reg_module/_08920_ ),
    .A2(\reg_module/_08923_ ),
    .B1(\reg_module/_08906_ ),
    .Y(\reg_module/_00280_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16540_  (.A(\reg_module/_08919_ ),
    .B(net1611),
    .Y(\reg_module/_08924_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16541_  (.A(\reg_module/_07597_ ),
    .B(\reg_module/_08921_ ),
    .Y(\reg_module/_08925_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16542_  (.A(\reg_module/_08903_ ),
    .B(\reg_module/_08925_ ),
    .Y(\reg_module/_08926_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16543_  (.A1(\reg_module/_08924_ ),
    .A2(\reg_module/_08926_ ),
    .B1(\reg_module/_08906_ ),
    .Y(\reg_module/_00281_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16544_  (.A(\reg_module/_08919_ ),
    .B(net1940),
    .Y(\reg_module/_08927_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16545_  (.A(\reg_module/_08873_ ),
    .X(\reg_module/_08928_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16546_  (.A(\reg_module/_07600_ ),
    .B(\reg_module/_08921_ ),
    .Y(\reg_module/_08929_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16547_  (.A(\reg_module/_08928_ ),
    .B(\reg_module/_08929_ ),
    .Y(\reg_module/_08930_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16548_  (.A(\reg_module/_08877_ ),
    .X(\reg_module/_08931_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16549_  (.A1(\reg_module/_08927_ ),
    .A2(\reg_module/_08930_ ),
    .B1(\reg_module/_08931_ ),
    .Y(\reg_module/_00282_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16550_  (.A(\reg_module/_08919_ ),
    .B(net1895),
    .Y(\reg_module/_08932_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16551_  (.A(\reg_module/_07603_ ),
    .B(\reg_module/_08921_ ),
    .Y(\reg_module/_08933_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16552_  (.A(\reg_module/_08928_ ),
    .B(\reg_module/_08933_ ),
    .Y(\reg_module/_08934_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16553_  (.A1(\reg_module/_08932_ ),
    .A2(\reg_module/_08934_ ),
    .B1(\reg_module/_08931_ ),
    .Y(\reg_module/_00283_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16554_  (.A(\reg_module/_08919_ ),
    .B(net1746),
    .Y(\reg_module/_08935_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16555_  (.A(\reg_module/_07606_ ),
    .B(\reg_module/_08921_ ),
    .Y(\reg_module/_08936_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16556_  (.A(\reg_module/_08928_ ),
    .B(\reg_module/_08936_ ),
    .Y(\reg_module/_08937_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16557_  (.A1(\reg_module/_08935_ ),
    .A2(\reg_module/_08937_ ),
    .B1(\reg_module/_08931_ ),
    .Y(\reg_module/_00284_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16558_  (.A(\reg_module/_08919_ ),
    .B(net1510),
    .Y(\reg_module/_08938_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16559_  (.A(\reg_module/_07609_ ),
    .B(\reg_module/_08921_ ),
    .Y(\reg_module/_08939_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16560_  (.A(\reg_module/_08928_ ),
    .B(\reg_module/_08939_ ),
    .Y(\reg_module/_08940_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16561_  (.A1(\reg_module/_08938_ ),
    .A2(\reg_module/_08940_ ),
    .B1(\reg_module/_08931_ ),
    .Y(\reg_module/_00285_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16562_  (.A(\reg_module/_08830_ ),
    .B(net1688),
    .Y(\reg_module/_08941_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16563_  (.A(\reg_module/_07612_ ),
    .B(\reg_module/_08837_ ),
    .Y(\reg_module/_08942_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16564_  (.A(\reg_module/_08928_ ),
    .B(\reg_module/_08942_ ),
    .Y(\reg_module/_08943_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16565_  (.A1(\reg_module/_08941_ ),
    .A2(\reg_module/_08943_ ),
    .B1(\reg_module/_08931_ ),
    .Y(\reg_module/_00286_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16566_  (.A(\reg_module/_08830_ ),
    .B(net1507),
    .Y(\reg_module/_08944_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16567_  (.A(\reg_module/_07615_ ),
    .B(\reg_module/_08837_ ),
    .Y(\reg_module/_08945_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16568_  (.A(\reg_module/_08928_ ),
    .B(\reg_module/_08945_ ),
    .Y(\reg_module/_08946_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16569_  (.A1(\reg_module/_08944_ ),
    .A2(\reg_module/_08946_ ),
    .B1(\reg_module/_08931_ ),
    .Y(\reg_module/_00287_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16570_  (.A(net963),
    .B(\reg_module/_07629_ ),
    .Y(\reg_module/_08947_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16571_  (.A(\reg_module/_07620_ ),
    .B(\reg_module/_07624_ ),
    .C(\reg_module/_08947_ ),
    .Y(\reg_module/_08948_ ));
 sky130_fd_sc_hd__buf_8 \reg_module/_16572_  (.A(\reg_module/_08948_ ),
    .X(\reg_module/_08949_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16573_  (.A(\reg_module/_08949_ ),
    .X(\reg_module/_08950_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16574_  (.A(\reg_module/_08950_ ),
    .B(net1390),
    .Y(\reg_module/_08951_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16575_  (.A(\reg_module/_07644_ ),
    .Y(\reg_module/_08952_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_16576_  (.A(\reg_module/_08952_ ),
    .X(\reg_module/_08953_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16577_  (.A(\reg_module/_08953_ ),
    .X(\reg_module/_08954_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16578_  (.A(\reg_module/_08954_ ),
    .X(\reg_module/_08955_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16579_  (.A(\reg_module/_07650_ ),
    .B(\reg_module/_08955_ ),
    .Y(\reg_module/_08956_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_16580_  (.A(\reg_module/_07639_ ),
    .X(\reg_module/_08957_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_16581_  (.A(\reg_module/_08957_ ),
    .X(\reg_module/_08958_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16582_  (.A(\reg_module/_08956_ ),
    .B(\reg_module/_08958_ ),
    .Y(\reg_module/_08959_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16583_  (.A(\reg_module/_08877_ ),
    .X(\reg_module/_08960_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16584_  (.A1(\reg_module/_08951_ ),
    .A2(\reg_module/_08959_ ),
    .B1(\reg_module/_08960_ ),
    .Y(\reg_module/_00288_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16585_  (.A(\reg_module/_08950_ ),
    .B(net1378),
    .Y(\reg_module/_08961_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16586_  (.A(\reg_module/_07658_ ),
    .B(\reg_module/_08955_ ),
    .Y(\reg_module/_08962_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16587_  (.A(\reg_module/_08962_ ),
    .B(\reg_module/_08958_ ),
    .Y(\reg_module/_08963_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16588_  (.A1(\reg_module/_08961_ ),
    .A2(\reg_module/_08963_ ),
    .B1(\reg_module/_08960_ ),
    .Y(\reg_module/_00289_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16589_  (.A(\reg_module/_08950_ ),
    .B(net1739),
    .Y(\reg_module/_08964_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16590_  (.A(\reg_module/_07664_ ),
    .B(\reg_module/_08955_ ),
    .Y(\reg_module/_08965_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16591_  (.A(\reg_module/_08965_ ),
    .B(\reg_module/_08958_ ),
    .Y(\reg_module/_08966_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16592_  (.A1(\reg_module/_08964_ ),
    .A2(\reg_module/_08966_ ),
    .B1(\reg_module/_08960_ ),
    .Y(\reg_module/_00290_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16593_  (.A(\reg_module/_08950_ ),
    .B(net1234),
    .Y(\reg_module/_08967_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16594_  (.A(\reg_module/_07668_ ),
    .B(\reg_module/_08955_ ),
    .Y(\reg_module/_08968_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16595_  (.A(\reg_module/_08968_ ),
    .B(\reg_module/_08958_ ),
    .Y(\reg_module/_08969_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16596_  (.A1(\reg_module/_08967_ ),
    .A2(\reg_module/_08969_ ),
    .B1(\reg_module/_08960_ ),
    .Y(\reg_module/_00291_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16597_  (.A(\reg_module/_08950_ ),
    .B(net1529),
    .Y(\reg_module/_08970_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16598_  (.A(\reg_module/_07672_ ),
    .B(\reg_module/_08955_ ),
    .Y(\reg_module/_08971_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16599_  (.A(\reg_module/_08957_ ),
    .X(\reg_module/_08972_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16600_  (.A(\reg_module/_08971_ ),
    .B(\reg_module/_08972_ ),
    .Y(\reg_module/_08973_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16601_  (.A1(\reg_module/_08970_ ),
    .A2(\reg_module/_08973_ ),
    .B1(\reg_module/_08960_ ),
    .Y(\reg_module/_00292_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16602_  (.A(\reg_module/_08950_ ),
    .B(net1612),
    .Y(\reg_module/_08974_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16603_  (.A(\reg_module/_07676_ ),
    .B(\reg_module/_08955_ ),
    .Y(\reg_module/_08975_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16604_  (.A(\reg_module/_08975_ ),
    .B(\reg_module/_08972_ ),
    .Y(\reg_module/_08976_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16605_  (.A1(\reg_module/_08974_ ),
    .A2(\reg_module/_08976_ ),
    .B1(\reg_module/_08960_ ),
    .Y(\reg_module/_00293_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16606_  (.A(\reg_module/_08949_ ),
    .X(\reg_module/_08977_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16607_  (.A(\reg_module/_08977_ ),
    .B(net1621),
    .Y(\reg_module/_08978_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16608_  (.A(\reg_module/_08954_ ),
    .X(\reg_module/_08979_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16609_  (.A(\reg_module/_07683_ ),
    .B(\reg_module/_08979_ ),
    .Y(\reg_module/_08980_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16610_  (.A(\reg_module/_08980_ ),
    .B(\reg_module/_08972_ ),
    .Y(\reg_module/_08981_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16611_  (.A(\reg_module/_08877_ ),
    .X(\reg_module/_08982_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16612_  (.A1(\reg_module/_08978_ ),
    .A2(\reg_module/_08981_ ),
    .B1(\reg_module/_08982_ ),
    .Y(\reg_module/_00294_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16613_  (.A(\reg_module/_08977_ ),
    .B(net1337),
    .Y(\reg_module/_08983_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16614_  (.A(\reg_module/_07688_ ),
    .B(\reg_module/_08979_ ),
    .Y(\reg_module/_08984_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16615_  (.A(\reg_module/_08984_ ),
    .B(\reg_module/_08972_ ),
    .Y(\reg_module/_08985_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16616_  (.A1(\reg_module/_08983_ ),
    .A2(\reg_module/_08985_ ),
    .B1(\reg_module/_08982_ ),
    .Y(\reg_module/_00295_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16617_  (.A(\reg_module/_08977_ ),
    .B(net1260),
    .Y(\reg_module/_08986_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16618_  (.A(\reg_module/_07693_ ),
    .B(\reg_module/_08979_ ),
    .Y(\reg_module/_08987_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16619_  (.A(\reg_module/_08987_ ),
    .B(\reg_module/_08972_ ),
    .Y(\reg_module/_08988_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16620_  (.A1(\reg_module/_08986_ ),
    .A2(\reg_module/_08988_ ),
    .B1(\reg_module/_08982_ ),
    .Y(\reg_module/_00296_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16621_  (.A(\reg_module/_08977_ ),
    .B(net1278),
    .Y(\reg_module/_08989_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16622_  (.A(\reg_module/_07697_ ),
    .B(\reg_module/_08979_ ),
    .Y(\reg_module/_08990_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16623_  (.A(\reg_module/_08990_ ),
    .B(\reg_module/_08972_ ),
    .Y(\reg_module/_08991_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16624_  (.A1(\reg_module/_08989_ ),
    .A2(\reg_module/_08991_ ),
    .B1(\reg_module/_08982_ ),
    .Y(\reg_module/_00297_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16625_  (.A(\reg_module/_08977_ ),
    .B(net1292),
    .Y(\reg_module/_08992_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16626_  (.A(\reg_module/_07701_ ),
    .B(\reg_module/_08979_ ),
    .Y(\reg_module/_08993_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16627_  (.A(\reg_module/_07639_ ),
    .X(\reg_module/_08994_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16628_  (.A(\reg_module/_08994_ ),
    .X(\reg_module/_08995_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16629_  (.A(\reg_module/_08993_ ),
    .B(\reg_module/_08995_ ),
    .Y(\reg_module/_08996_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16630_  (.A1(\reg_module/_08992_ ),
    .A2(\reg_module/_08996_ ),
    .B1(\reg_module/_08982_ ),
    .Y(\reg_module/_00298_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16631_  (.A(\reg_module/_08977_ ),
    .B(net1467),
    .Y(\reg_module/_08997_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16632_  (.A(\reg_module/_07705_ ),
    .B(\reg_module/_08979_ ),
    .Y(\reg_module/_08998_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16633_  (.A(\reg_module/_08998_ ),
    .B(\reg_module/_08995_ ),
    .Y(\reg_module/_08999_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16634_  (.A1(\reg_module/_08997_ ),
    .A2(\reg_module/_08999_ ),
    .B1(\reg_module/_08982_ ),
    .Y(\reg_module/_00299_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16635_  (.A(\reg_module/_08949_ ),
    .X(\reg_module/_09000_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16636_  (.A(\reg_module/_09000_ ),
    .B(net1429),
    .Y(\reg_module/_09001_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16637_  (.A(\reg_module/_08954_ ),
    .X(\reg_module/_09002_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16638_  (.A(\reg_module/_07712_ ),
    .B(\reg_module/_09002_ ),
    .Y(\reg_module/_09003_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16639_  (.A(\reg_module/_09003_ ),
    .B(\reg_module/_08995_ ),
    .Y(\reg_module/_09004_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16640_  (.A(\reg_module/_08877_ ),
    .X(\reg_module/_09005_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16641_  (.A1(\reg_module/_09001_ ),
    .A2(\reg_module/_09004_ ),
    .B1(\reg_module/_09005_ ),
    .Y(\reg_module/_00300_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16642_  (.A(\reg_module/_09000_ ),
    .B(net1847),
    .Y(\reg_module/_09006_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16643_  (.A(\reg_module/_07717_ ),
    .B(\reg_module/_09002_ ),
    .Y(\reg_module/_09007_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16644_  (.A(\reg_module/_09007_ ),
    .B(\reg_module/_08995_ ),
    .Y(\reg_module/_09008_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16645_  (.A1(\reg_module/_09006_ ),
    .A2(\reg_module/_09008_ ),
    .B1(\reg_module/_09005_ ),
    .Y(\reg_module/_00301_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16646_  (.A(\reg_module/_09000_ ),
    .B(net1670),
    .Y(\reg_module/_09009_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16647_  (.A(\reg_module/_07722_ ),
    .B(\reg_module/_09002_ ),
    .Y(\reg_module/_09010_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16648_  (.A(\reg_module/_09010_ ),
    .B(\reg_module/_08995_ ),
    .Y(\reg_module/_09011_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16649_  (.A1(\reg_module/_09009_ ),
    .A2(\reg_module/_09011_ ),
    .B1(\reg_module/_09005_ ),
    .Y(\reg_module/_00302_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16650_  (.A(\reg_module/_09000_ ),
    .B(net1500),
    .Y(\reg_module/_09012_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16651_  (.A(\reg_module/_07726_ ),
    .B(\reg_module/_09002_ ),
    .Y(\reg_module/_09013_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16652_  (.A(\reg_module/_09013_ ),
    .B(\reg_module/_08995_ ),
    .Y(\reg_module/_09014_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16653_  (.A1(\reg_module/_09012_ ),
    .A2(\reg_module/_09014_ ),
    .B1(\reg_module/_09005_ ),
    .Y(\reg_module/_00303_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16654_  (.A(\reg_module/_09000_ ),
    .B(net1380),
    .Y(\reg_module/_09015_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16655_  (.A(\reg_module/_07730_ ),
    .B(\reg_module/_09002_ ),
    .Y(\reg_module/_09016_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16656_  (.A(\reg_module/_08994_ ),
    .X(\reg_module/_09017_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16657_  (.A(\reg_module/_09016_ ),
    .B(\reg_module/_09017_ ),
    .Y(\reg_module/_09018_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16658_  (.A1(\reg_module/_09015_ ),
    .A2(\reg_module/_09018_ ),
    .B1(\reg_module/_09005_ ),
    .Y(\reg_module/_00304_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16659_  (.A(\reg_module/_09000_ ),
    .B(net1239),
    .Y(\reg_module/_09019_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16660_  (.A(\reg_module/_07734_ ),
    .B(\reg_module/_09002_ ),
    .Y(\reg_module/_09020_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16661_  (.A(\reg_module/_09020_ ),
    .B(\reg_module/_09017_ ),
    .Y(\reg_module/_09021_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16662_  (.A1(\reg_module/_09019_ ),
    .A2(\reg_module/_09021_ ),
    .B1(\reg_module/_09005_ ),
    .Y(\reg_module/_00305_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16663_  (.A(\reg_module/_08949_ ),
    .X(\reg_module/_09022_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16664_  (.A(\reg_module/_09022_ ),
    .B(net1884),
    .Y(\reg_module/_09023_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16665_  (.A(\reg_module/_08954_ ),
    .X(\reg_module/_09024_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16666_  (.A(\reg_module/_07741_ ),
    .B(\reg_module/_09024_ ),
    .Y(\reg_module/_09025_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16667_  (.A(\reg_module/_09025_ ),
    .B(\reg_module/_09017_ ),
    .Y(\reg_module/_09026_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16668_  (.A(\reg_module/_07993_ ),
    .X(\reg_module/_09027_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16669_  (.A(\reg_module/_09027_ ),
    .X(\reg_module/_09028_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16670_  (.A1(\reg_module/_09023_ ),
    .A2(\reg_module/_09026_ ),
    .B1(\reg_module/_09028_ ),
    .Y(\reg_module/_00306_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16671_  (.A(\reg_module/_09022_ ),
    .B(net1671),
    .Y(\reg_module/_09029_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16672_  (.A(\reg_module/_07746_ ),
    .B(\reg_module/_09024_ ),
    .Y(\reg_module/_09030_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16673_  (.A(\reg_module/_09030_ ),
    .B(\reg_module/_09017_ ),
    .Y(\reg_module/_09031_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16674_  (.A1(\reg_module/_09029_ ),
    .A2(\reg_module/_09031_ ),
    .B1(\reg_module/_09028_ ),
    .Y(\reg_module/_00307_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16675_  (.A(\reg_module/_09022_ ),
    .B(net1283),
    .Y(\reg_module/_09032_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16676_  (.A(\reg_module/_07751_ ),
    .B(\reg_module/_09024_ ),
    .Y(\reg_module/_09033_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16677_  (.A(\reg_module/_09033_ ),
    .B(\reg_module/_09017_ ),
    .Y(\reg_module/_09034_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16678_  (.A1(\reg_module/_09032_ ),
    .A2(\reg_module/_09034_ ),
    .B1(\reg_module/_09028_ ),
    .Y(\reg_module/_00308_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16679_  (.A(\reg_module/_09022_ ),
    .B(net1327),
    .Y(\reg_module/_09035_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16680_  (.A(\reg_module/_07755_ ),
    .B(\reg_module/_09024_ ),
    .Y(\reg_module/_09036_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16681_  (.A(\reg_module/_09036_ ),
    .B(\reg_module/_09017_ ),
    .Y(\reg_module/_09037_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16682_  (.A1(\reg_module/_09035_ ),
    .A2(\reg_module/_09037_ ),
    .B1(\reg_module/_09028_ ),
    .Y(\reg_module/_00309_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16683_  (.A(\reg_module/_09022_ ),
    .B(net1367),
    .Y(\reg_module/_09038_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16684_  (.A(\reg_module/_07759_ ),
    .B(\reg_module/_09024_ ),
    .Y(\reg_module/_09039_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16685_  (.A(\reg_module/_08994_ ),
    .X(\reg_module/_09040_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16686_  (.A(\reg_module/_09039_ ),
    .B(\reg_module/_09040_ ),
    .Y(\reg_module/_09041_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16687_  (.A1(\reg_module/_09038_ ),
    .A2(\reg_module/_09041_ ),
    .B1(\reg_module/_09028_ ),
    .Y(\reg_module/_00310_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16688_  (.A(\reg_module/_09022_ ),
    .B(net1778),
    .Y(\reg_module/_09042_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16689_  (.A(\reg_module/_07763_ ),
    .B(\reg_module/_09024_ ),
    .Y(\reg_module/_09043_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16690_  (.A(\reg_module/_09043_ ),
    .B(\reg_module/_09040_ ),
    .Y(\reg_module/_09044_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16691_  (.A1(\reg_module/_09042_ ),
    .A2(\reg_module/_09044_ ),
    .B1(\reg_module/_09028_ ),
    .Y(\reg_module/_00311_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16692_  (.A(\reg_module/_08948_ ),
    .X(\reg_module/_09045_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16693_  (.A(\reg_module/_09045_ ),
    .B(net1806),
    .Y(\reg_module/_09046_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_16694_  (.A(\reg_module/_08952_ ),
    .X(\reg_module/_09047_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16695_  (.A(\reg_module/_09047_ ),
    .X(\reg_module/_09048_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16696_  (.A(\reg_module/_07771_ ),
    .B(\reg_module/_09048_ ),
    .Y(\reg_module/_09049_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16697_  (.A(\reg_module/_09049_ ),
    .B(\reg_module/_09040_ ),
    .Y(\reg_module/_09050_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16698_  (.A(\reg_module/_09027_ ),
    .X(\reg_module/_09051_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16699_  (.A1(\reg_module/_09046_ ),
    .A2(\reg_module/_09050_ ),
    .B1(\reg_module/_09051_ ),
    .Y(\reg_module/_00312_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16700_  (.A(\reg_module/_09045_ ),
    .B(net1741),
    .Y(\reg_module/_09052_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16701_  (.A(\reg_module/_07777_ ),
    .B(\reg_module/_09048_ ),
    .Y(\reg_module/_09053_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16702_  (.A(\reg_module/_09053_ ),
    .B(\reg_module/_09040_ ),
    .Y(\reg_module/_09054_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16703_  (.A1(\reg_module/_09052_ ),
    .A2(\reg_module/_09054_ ),
    .B1(\reg_module/_09051_ ),
    .Y(\reg_module/_00313_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16704_  (.A(\reg_module/_09045_ ),
    .B(net1275),
    .Y(\reg_module/_09055_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16705_  (.A(\reg_module/_07783_ ),
    .B(\reg_module/_09048_ ),
    .Y(\reg_module/_09056_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16706_  (.A(\reg_module/_09056_ ),
    .B(\reg_module/_09040_ ),
    .Y(\reg_module/_09057_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16707_  (.A1(\reg_module/_09055_ ),
    .A2(\reg_module/_09057_ ),
    .B1(\reg_module/_09051_ ),
    .Y(\reg_module/_00314_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16708_  (.A(\reg_module/_09045_ ),
    .B(net1555),
    .Y(\reg_module/_09058_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16709_  (.A(\reg_module/_07787_ ),
    .B(\reg_module/_09048_ ),
    .Y(\reg_module/_09059_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16710_  (.A(\reg_module/_09059_ ),
    .B(\reg_module/_09040_ ),
    .Y(\reg_module/_09060_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16711_  (.A1(\reg_module/_09058_ ),
    .A2(\reg_module/_09060_ ),
    .B1(\reg_module/_09051_ ),
    .Y(\reg_module/_00315_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16712_  (.A(\reg_module/_09045_ ),
    .B(net1496),
    .Y(\reg_module/_09061_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16713_  (.A(\reg_module/_07791_ ),
    .B(\reg_module/_09048_ ),
    .Y(\reg_module/_09062_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16714_  (.A(\reg_module/_08994_ ),
    .X(\reg_module/_09063_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16715_  (.A(\reg_module/_09062_ ),
    .B(\reg_module/_09063_ ),
    .Y(\reg_module/_09064_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16716_  (.A1(\reg_module/_09061_ ),
    .A2(\reg_module/_09064_ ),
    .B1(\reg_module/_09051_ ),
    .Y(\reg_module/_00316_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16717_  (.A(\reg_module/_09045_ ),
    .B(net1277),
    .Y(\reg_module/_09065_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16718_  (.A(\reg_module/_07795_ ),
    .B(\reg_module/_09048_ ),
    .Y(\reg_module/_09066_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16719_  (.A(\reg_module/_09066_ ),
    .B(\reg_module/_09063_ ),
    .Y(\reg_module/_09067_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16720_  (.A1(\reg_module/_09065_ ),
    .A2(\reg_module/_09067_ ),
    .B1(\reg_module/_09051_ ),
    .Y(\reg_module/_00317_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16721_  (.A(\reg_module/_08949_ ),
    .B(net1916),
    .Y(\reg_module/_09068_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16722_  (.A(\reg_module/_09047_ ),
    .X(\reg_module/_09069_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16723_  (.A(\reg_module/_07800_ ),
    .B(\reg_module/_09069_ ),
    .Y(\reg_module/_09070_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16724_  (.A(\reg_module/_09070_ ),
    .B(\reg_module/_09063_ ),
    .Y(\reg_module/_09071_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16725_  (.A(\reg_module/_09027_ ),
    .X(\reg_module/_09072_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16726_  (.A1(\reg_module/_09068_ ),
    .A2(\reg_module/_09071_ ),
    .B1(\reg_module/_09072_ ),
    .Y(\reg_module/_00318_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16727_  (.A(\reg_module/_08949_ ),
    .B(net1692),
    .Y(\reg_module/_09073_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16728_  (.A(\reg_module/_07805_ ),
    .B(\reg_module/_09069_ ),
    .Y(\reg_module/_09074_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16729_  (.A(\reg_module/_09074_ ),
    .B(\reg_module/_09063_ ),
    .Y(\reg_module/_09075_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16730_  (.A1(\reg_module/_09073_ ),
    .A2(\reg_module/_09075_ ),
    .B1(\reg_module/_09072_ ),
    .Y(\reg_module/_00319_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16731_  (.A(net965),
    .B(\reg_module/_07809_ ),
    .Y(\reg_module/_09076_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16732_  (.A(\reg_module/_07619_ ),
    .B(\reg_module/_08825_ ),
    .C(\reg_module/_09076_ ),
    .Y(\reg_module/_09077_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_16733_  (.A(\reg_module/_09077_ ),
    .X(\reg_module/_09078_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16734_  (.A(\reg_module/_09078_ ),
    .X(\reg_module/_09079_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16735_  (.A(\reg_module/_09079_ ),
    .B(net1450),
    .Y(\reg_module/_09080_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16736_  (.A(\reg_module/_07822_ ),
    .B(\reg_module/_09069_ ),
    .Y(\reg_module/_09081_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16737_  (.A(\reg_module/_09081_ ),
    .B(\reg_module/_09063_ ),
    .Y(\reg_module/_09082_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16738_  (.A1(\reg_module/_09080_ ),
    .A2(\reg_module/_09082_ ),
    .B1(\reg_module/_09072_ ),
    .Y(\reg_module/_00320_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16739_  (.A(\reg_module/_09079_ ),
    .B(net1350),
    .Y(\reg_module/_09083_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16740_  (.A(\reg_module/_07827_ ),
    .B(\reg_module/_09069_ ),
    .Y(\reg_module/_09084_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16741_  (.A(\reg_module/_09084_ ),
    .B(\reg_module/_09063_ ),
    .Y(\reg_module/_09085_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16742_  (.A1(\reg_module/_09083_ ),
    .A2(\reg_module/_09085_ ),
    .B1(\reg_module/_09072_ ),
    .Y(\reg_module/_00321_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16743_  (.A(\reg_module/_09079_ ),
    .B(net1481),
    .Y(\reg_module/_09086_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16744_  (.A(\reg_module/_07832_ ),
    .B(\reg_module/_09069_ ),
    .Y(\reg_module/_09087_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16745_  (.A(\reg_module/_08994_ ),
    .X(\reg_module/_09088_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16746_  (.A(\reg_module/_09087_ ),
    .B(\reg_module/_09088_ ),
    .Y(\reg_module/_09089_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16747_  (.A1(\reg_module/_09086_ ),
    .A2(\reg_module/_09089_ ),
    .B1(\reg_module/_09072_ ),
    .Y(\reg_module/_00322_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16748_  (.A(\reg_module/_09079_ ),
    .B(net1377),
    .Y(\reg_module/_09090_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16749_  (.A(\reg_module/_07837_ ),
    .B(\reg_module/_09069_ ),
    .Y(\reg_module/_09091_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16750_  (.A(\reg_module/_09091_ ),
    .B(\reg_module/_09088_ ),
    .Y(\reg_module/_09092_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16751_  (.A1(\reg_module/_09090_ ),
    .A2(\reg_module/_09092_ ),
    .B1(\reg_module/_09072_ ),
    .Y(\reg_module/_00323_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16752_  (.A(\reg_module/_09079_ ),
    .B(net1526),
    .Y(\reg_module/_09093_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16753_  (.A(\reg_module/_09047_ ),
    .X(\reg_module/_09094_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16754_  (.A(\reg_module/_07845_ ),
    .B(\reg_module/_09094_ ),
    .Y(\reg_module/_09095_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16755_  (.A(\reg_module/_09095_ ),
    .B(\reg_module/_09088_ ),
    .Y(\reg_module/_09096_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16756_  (.A(\reg_module/_09027_ ),
    .X(\reg_module/_09097_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16757_  (.A1(\reg_module/_09093_ ),
    .A2(\reg_module/_09096_ ),
    .B1(\reg_module/_09097_ ),
    .Y(\reg_module/_00324_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16758_  (.A(\reg_module/_09079_ ),
    .B(net1552),
    .Y(\reg_module/_09098_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16759_  (.A(\reg_module/_07851_ ),
    .B(\reg_module/_09094_ ),
    .Y(\reg_module/_09099_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16760_  (.A(\reg_module/_09099_ ),
    .B(\reg_module/_09088_ ),
    .Y(\reg_module/_09100_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16761_  (.A1(\reg_module/_09098_ ),
    .A2(\reg_module/_09100_ ),
    .B1(\reg_module/_09097_ ),
    .Y(\reg_module/_00325_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16762_  (.A(\reg_module/_09078_ ),
    .X(\reg_module/_09101_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16763_  (.A(\reg_module/_09101_ ),
    .B(net1527),
    .Y(\reg_module/_09102_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16764_  (.A(\reg_module/_07859_ ),
    .B(\reg_module/_09094_ ),
    .Y(\reg_module/_09103_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16765_  (.A(\reg_module/_09103_ ),
    .B(\reg_module/_09088_ ),
    .Y(\reg_module/_09104_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16766_  (.A1(\reg_module/_09102_ ),
    .A2(\reg_module/_09104_ ),
    .B1(\reg_module/_09097_ ),
    .Y(\reg_module/_00326_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16767_  (.A(\reg_module/_09101_ ),
    .B(net1604),
    .Y(\reg_module/_09105_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16768_  (.A(\reg_module/_07864_ ),
    .B(\reg_module/_09094_ ),
    .Y(\reg_module/_09106_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16769_  (.A(\reg_module/_09106_ ),
    .B(\reg_module/_09088_ ),
    .Y(\reg_module/_09107_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16770_  (.A1(\reg_module/_09105_ ),
    .A2(\reg_module/_09107_ ),
    .B1(\reg_module/_09097_ ),
    .Y(\reg_module/_00327_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16771_  (.A(\reg_module/_09101_ ),
    .B(net1424),
    .Y(\reg_module/_09108_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16772_  (.A(\reg_module/_07869_ ),
    .B(\reg_module/_09094_ ),
    .Y(\reg_module/_09109_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16773_  (.A(\reg_module/_08994_ ),
    .X(\reg_module/_09110_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16774_  (.A(\reg_module/_09109_ ),
    .B(\reg_module/_09110_ ),
    .Y(\reg_module/_09111_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16775_  (.A1(\reg_module/_09108_ ),
    .A2(\reg_module/_09111_ ),
    .B1(\reg_module/_09097_ ),
    .Y(\reg_module/_00328_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16776_  (.A(\reg_module/_09101_ ),
    .B(net1406),
    .Y(\reg_module/_09112_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16777_  (.A(\reg_module/_07874_ ),
    .B(\reg_module/_09094_ ),
    .Y(\reg_module/_09113_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16778_  (.A(\reg_module/_09113_ ),
    .B(\reg_module/_09110_ ),
    .Y(\reg_module/_09114_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16779_  (.A1(\reg_module/_09112_ ),
    .A2(\reg_module/_09114_ ),
    .B1(\reg_module/_09097_ ),
    .Y(\reg_module/_00329_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16780_  (.A(\reg_module/_09101_ ),
    .B(net1473),
    .Y(\reg_module/_09115_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16781_  (.A(\reg_module/_09047_ ),
    .X(\reg_module/_09116_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16782_  (.A(\reg_module/_07881_ ),
    .B(\reg_module/_09116_ ),
    .Y(\reg_module/_09117_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16783_  (.A(\reg_module/_09117_ ),
    .B(\reg_module/_09110_ ),
    .Y(\reg_module/_09118_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16784_  (.A(\reg_module/_09027_ ),
    .X(\reg_module/_09119_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16785_  (.A1(\reg_module/_09115_ ),
    .A2(\reg_module/_09118_ ),
    .B1(\reg_module/_09119_ ),
    .Y(\reg_module/_00330_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16786_  (.A(\reg_module/_09101_ ),
    .B(net1356),
    .Y(\reg_module/_09120_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16787_  (.A(\reg_module/_07887_ ),
    .B(\reg_module/_09116_ ),
    .Y(\reg_module/_09121_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16788_  (.A(\reg_module/_09121_ ),
    .B(\reg_module/_09110_ ),
    .Y(\reg_module/_09122_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16789_  (.A1(\reg_module/_09120_ ),
    .A2(\reg_module/_09122_ ),
    .B1(\reg_module/_09119_ ),
    .Y(\reg_module/_00331_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16790_  (.A(\reg_module/_09078_ ),
    .X(\reg_module/_09123_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16791_  (.A(\reg_module/_09123_ ),
    .B(net1549),
    .Y(\reg_module/_09124_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16792_  (.A(\reg_module/_07895_ ),
    .B(\reg_module/_09116_ ),
    .Y(\reg_module/_09125_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16793_  (.A(\reg_module/_09125_ ),
    .B(\reg_module/_09110_ ),
    .Y(\reg_module/_09126_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16794_  (.A1(\reg_module/_09124_ ),
    .A2(\reg_module/_09126_ ),
    .B1(\reg_module/_09119_ ),
    .Y(\reg_module/_00332_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16795_  (.A(\reg_module/_09123_ ),
    .B(net1501),
    .Y(\reg_module/_09127_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16796_  (.A(\reg_module/_07900_ ),
    .B(\reg_module/_09116_ ),
    .Y(\reg_module/_09128_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16797_  (.A(\reg_module/_09128_ ),
    .B(\reg_module/_09110_ ),
    .Y(\reg_module/_09129_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16798_  (.A1(\reg_module/_09127_ ),
    .A2(\reg_module/_09129_ ),
    .B1(\reg_module/_09119_ ),
    .Y(\reg_module/_00333_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16799_  (.A(\reg_module/_09123_ ),
    .B(net1295),
    .Y(\reg_module/_09130_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16800_  (.A(\reg_module/_07905_ ),
    .B(\reg_module/_09116_ ),
    .Y(\reg_module/_09131_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16801_  (.A(\reg_module/_07639_ ),
    .X(\reg_module/_09132_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16802_  (.A(\reg_module/_09132_ ),
    .X(\reg_module/_09133_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16803_  (.A(\reg_module/_09131_ ),
    .B(\reg_module/_09133_ ),
    .Y(\reg_module/_09134_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16804_  (.A1(\reg_module/_09130_ ),
    .A2(\reg_module/_09134_ ),
    .B1(\reg_module/_09119_ ),
    .Y(\reg_module/_00334_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16805_  (.A(\reg_module/_09123_ ),
    .B(net1491),
    .Y(\reg_module/_09135_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16806_  (.A(\reg_module/_07910_ ),
    .B(\reg_module/_09116_ ),
    .Y(\reg_module/_09136_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16807_  (.A(\reg_module/_09136_ ),
    .B(\reg_module/_09133_ ),
    .Y(\reg_module/_09137_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16808_  (.A1(\reg_module/_09135_ ),
    .A2(\reg_module/_09137_ ),
    .B1(\reg_module/_09119_ ),
    .Y(\reg_module/_00335_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16809_  (.A(\reg_module/_09123_ ),
    .B(net1813),
    .Y(\reg_module/_09138_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16810_  (.A(\reg_module/_09047_ ),
    .X(\reg_module/_09139_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16811_  (.A(\reg_module/_07917_ ),
    .B(\reg_module/_09139_ ),
    .Y(\reg_module/_09140_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16812_  (.A(\reg_module/_09140_ ),
    .B(\reg_module/_09133_ ),
    .Y(\reg_module/_09141_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16813_  (.A(\reg_module/_09027_ ),
    .X(\reg_module/_09142_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16814_  (.A1(\reg_module/_09138_ ),
    .A2(\reg_module/_09141_ ),
    .B1(\reg_module/_09142_ ),
    .Y(\reg_module/_00336_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16815_  (.A(\reg_module/_09123_ ),
    .B(net1465),
    .Y(\reg_module/_09143_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16816_  (.A(\reg_module/_07923_ ),
    .B(\reg_module/_09139_ ),
    .Y(\reg_module/_09144_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16817_  (.A(\reg_module/_09144_ ),
    .B(\reg_module/_09133_ ),
    .Y(\reg_module/_09145_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16818_  (.A1(\reg_module/_09143_ ),
    .A2(\reg_module/_09145_ ),
    .B1(\reg_module/_09142_ ),
    .Y(\reg_module/_00337_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16819_  (.A(\reg_module/_09078_ ),
    .X(\reg_module/_09146_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16820_  (.A(\reg_module/_09146_ ),
    .B(net1321),
    .Y(\reg_module/_09147_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16821_  (.A(\reg_module/_07931_ ),
    .B(\reg_module/_09139_ ),
    .Y(\reg_module/_09148_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16822_  (.A(\reg_module/_09148_ ),
    .B(\reg_module/_09133_ ),
    .Y(\reg_module/_09149_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16823_  (.A1(\reg_module/_09147_ ),
    .A2(\reg_module/_09149_ ),
    .B1(\reg_module/_09142_ ),
    .Y(\reg_module/_00338_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16824_  (.A(\reg_module/_09146_ ),
    .B(net1551),
    .Y(\reg_module/_09150_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16825_  (.A(\reg_module/_07936_ ),
    .B(\reg_module/_09139_ ),
    .Y(\reg_module/_09151_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16826_  (.A(\reg_module/_09151_ ),
    .B(\reg_module/_09133_ ),
    .Y(\reg_module/_09152_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16827_  (.A1(\reg_module/_09150_ ),
    .A2(\reg_module/_09152_ ),
    .B1(\reg_module/_09142_ ),
    .Y(\reg_module/_00339_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16828_  (.A(\reg_module/_09146_ ),
    .B(net1430),
    .Y(\reg_module/_09153_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16829_  (.A(\reg_module/_07941_ ),
    .B(\reg_module/_09139_ ),
    .Y(\reg_module/_09154_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16830_  (.A(\reg_module/_09132_ ),
    .X(\reg_module/_09155_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16831_  (.A(\reg_module/_09154_ ),
    .B(\reg_module/_09155_ ),
    .Y(\reg_module/_09156_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16832_  (.A1(\reg_module/_09153_ ),
    .A2(\reg_module/_09156_ ),
    .B1(\reg_module/_09142_ ),
    .Y(\reg_module/_00340_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16833_  (.A(\reg_module/_09146_ ),
    .B(net1472),
    .Y(\reg_module/_09157_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16834_  (.A(\reg_module/_07946_ ),
    .B(\reg_module/_09139_ ),
    .Y(\reg_module/_09158_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16835_  (.A(\reg_module/_09158_ ),
    .B(\reg_module/_09155_ ),
    .Y(\reg_module/_09159_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16836_  (.A1(\reg_module/_09157_ ),
    .A2(\reg_module/_09159_ ),
    .B1(\reg_module/_09142_ ),
    .Y(\reg_module/_00341_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16837_  (.A(\reg_module/_09146_ ),
    .B(net1518),
    .Y(\reg_module/_09160_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16838_  (.A(\reg_module/_09047_ ),
    .X(\reg_module/_09161_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16839_  (.A(\reg_module/_07953_ ),
    .B(\reg_module/_09161_ ),
    .Y(\reg_module/_09162_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16840_  (.A(\reg_module/_09162_ ),
    .B(\reg_module/_09155_ ),
    .Y(\reg_module/_09163_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_16841_  (.A(\reg_module/_07993_ ),
    .X(\reg_module/_09164_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16842_  (.A(\reg_module/_09164_ ),
    .X(\reg_module/_09165_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16843_  (.A1(\reg_module/_09160_ ),
    .A2(\reg_module/_09163_ ),
    .B1(\reg_module/_09165_ ),
    .Y(\reg_module/_00342_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16844_  (.A(\reg_module/_09146_ ),
    .B(net1399),
    .Y(\reg_module/_09166_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16845_  (.A(\reg_module/_07959_ ),
    .B(\reg_module/_09161_ ),
    .Y(\reg_module/_09167_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16846_  (.A(\reg_module/_09167_ ),
    .B(\reg_module/_09155_ ),
    .Y(\reg_module/_09168_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16847_  (.A1(\reg_module/_09166_ ),
    .A2(\reg_module/_09168_ ),
    .B1(\reg_module/_09165_ ),
    .Y(\reg_module/_00343_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16848_  (.A(\reg_module/_09077_ ),
    .X(\reg_module/_09169_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16849_  (.A(\reg_module/_09169_ ),
    .B(net1353),
    .Y(\reg_module/_09170_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16850_  (.A(\reg_module/_07967_ ),
    .B(\reg_module/_09161_ ),
    .Y(\reg_module/_09171_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16851_  (.A(\reg_module/_09171_ ),
    .B(\reg_module/_09155_ ),
    .Y(\reg_module/_09172_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16852_  (.A1(\reg_module/_09170_ ),
    .A2(\reg_module/_09172_ ),
    .B1(\reg_module/_09165_ ),
    .Y(\reg_module/_00344_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16853_  (.A(\reg_module/_09169_ ),
    .B(net1307),
    .Y(\reg_module/_09173_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16854_  (.A(\reg_module/_07972_ ),
    .B(\reg_module/_09161_ ),
    .Y(\reg_module/_09174_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16855_  (.A(\reg_module/_09174_ ),
    .B(\reg_module/_09155_ ),
    .Y(\reg_module/_09175_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16856_  (.A1(\reg_module/_09173_ ),
    .A2(\reg_module/_09175_ ),
    .B1(\reg_module/_09165_ ),
    .Y(\reg_module/_00345_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16857_  (.A(\reg_module/_09169_ ),
    .B(net1524),
    .Y(\reg_module/_09176_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16858_  (.A(\reg_module/_07977_ ),
    .B(\reg_module/_09161_ ),
    .Y(\reg_module/_09177_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16859_  (.A(\reg_module/_09132_ ),
    .X(\reg_module/_09178_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16860_  (.A(\reg_module/_09177_ ),
    .B(\reg_module/_09178_ ),
    .Y(\reg_module/_09179_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16861_  (.A1(\reg_module/_09176_ ),
    .A2(\reg_module/_09179_ ),
    .B1(\reg_module/_09165_ ),
    .Y(\reg_module/_00346_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16862_  (.A(\reg_module/_09169_ ),
    .B(net1444),
    .Y(\reg_module/_09180_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16863_  (.A(\reg_module/_07982_ ),
    .B(\reg_module/_09161_ ),
    .Y(\reg_module/_09181_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16864_  (.A(\reg_module/_09181_ ),
    .B(\reg_module/_09178_ ),
    .Y(\reg_module/_09182_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16865_  (.A1(\reg_module/_09180_ ),
    .A2(\reg_module/_09182_ ),
    .B1(\reg_module/_09165_ ),
    .Y(\reg_module/_00347_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16866_  (.A(\reg_module/_09169_ ),
    .B(net1329),
    .Y(\reg_module/_09183_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_16867_  (.A(\reg_module/_08952_ ),
    .X(\reg_module/_09184_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16868_  (.A(\reg_module/_09184_ ),
    .X(\reg_module/_09185_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16869_  (.A(\reg_module/_07990_ ),
    .B(\reg_module/_09185_ ),
    .Y(\reg_module/_09186_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16870_  (.A(\reg_module/_09186_ ),
    .B(\reg_module/_09178_ ),
    .Y(\reg_module/_09187_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16871_  (.A(\reg_module/_09164_ ),
    .X(\reg_module/_09188_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16872_  (.A1(\reg_module/_09183_ ),
    .A2(\reg_module/_09187_ ),
    .B1(\reg_module/_09188_ ),
    .Y(\reg_module/_00348_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16873_  (.A(\reg_module/_09169_ ),
    .B(net1708),
    .Y(\reg_module/_09189_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16874_  (.A(\reg_module/_07998_ ),
    .B(\reg_module/_09185_ ),
    .Y(\reg_module/_09190_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16875_  (.A(\reg_module/_09190_ ),
    .B(\reg_module/_09178_ ),
    .Y(\reg_module/_09191_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16876_  (.A1(\reg_module/_09189_ ),
    .A2(\reg_module/_09191_ ),
    .B1(\reg_module/_09188_ ),
    .Y(\reg_module/_00349_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16877_  (.A(\reg_module/_09078_ ),
    .B(net1506),
    .Y(\reg_module/_09192_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16878_  (.A(\reg_module/_08004_ ),
    .B(\reg_module/_09185_ ),
    .Y(\reg_module/_09193_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16879_  (.A(\reg_module/_09193_ ),
    .B(\reg_module/_09178_ ),
    .Y(\reg_module/_09194_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16880_  (.A1(\reg_module/_09192_ ),
    .A2(\reg_module/_09194_ ),
    .B1(\reg_module/_09188_ ),
    .Y(\reg_module/_00350_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16881_  (.A(\reg_module/_09078_ ),
    .B(net1391),
    .Y(\reg_module/_09195_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16882_  (.A(\reg_module/_08009_ ),
    .B(\reg_module/_09185_ ),
    .Y(\reg_module/_09196_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16883_  (.A(\reg_module/_09196_ ),
    .B(\reg_module/_09178_ ),
    .Y(\reg_module/_09197_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16884_  (.A1(\reg_module/_09195_ ),
    .A2(\reg_module/_09197_ ),
    .B1(\reg_module/_09188_ ),
    .Y(\reg_module/_00351_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16885_  (.A(\reg_module/_08013_ ),
    .B(\reg_module/_07625_ ),
    .Y(\reg_module/_09198_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_16886_  (.A(\reg_module/_09198_ ),
    .Y(\reg_module/_09199_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_16887_  (.A(\reg_module/_07619_ ),
    .B(\reg_module/_08825_ ),
    .C(\reg_module/_09199_ ),
    .Y(\reg_module/_09200_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16888_  (.A(\reg_module/_09200_ ),
    .X(\reg_module/_09201_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16889_  (.A(\reg_module/_09201_ ),
    .X(\reg_module/_09202_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16890_  (.A(\reg_module/_09202_ ),
    .B(net1715),
    .Y(\reg_module/_09203_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_16891_  (.A(\reg_module/_08873_ ),
    .X(\reg_module/_09204_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16892_  (.A(\reg_module/_08953_ ),
    .X(\reg_module/_09205_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16893_  (.A(\reg_module/_08022_ ),
    .B(\reg_module/_09205_ ),
    .Y(\reg_module/_09206_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16894_  (.A(\reg_module/_09204_ ),
    .B(\reg_module/_09206_ ),
    .Y(\reg_module/_09207_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16895_  (.A1(\reg_module/_09203_ ),
    .A2(\reg_module/_09207_ ),
    .B1(\reg_module/_09188_ ),
    .Y(\reg_module/_00352_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16896_  (.A(\reg_module/_09202_ ),
    .B(net1227),
    .Y(\reg_module/_09208_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16897_  (.A(\reg_module/_08027_ ),
    .B(\reg_module/_09205_ ),
    .Y(\reg_module/_09209_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16898_  (.A(\reg_module/_09204_ ),
    .B(\reg_module/_09209_ ),
    .Y(\reg_module/_09210_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16899_  (.A1(\reg_module/_09208_ ),
    .A2(\reg_module/_09210_ ),
    .B1(\reg_module/_09188_ ),
    .Y(\reg_module/_00353_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16900_  (.A(\reg_module/_09202_ ),
    .B(net1841),
    .Y(\reg_module/_09211_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16901_  (.A(\reg_module/_08034_ ),
    .B(\reg_module/_09205_ ),
    .Y(\reg_module/_09212_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16902_  (.A(\reg_module/_09204_ ),
    .B(\reg_module/_09212_ ),
    .Y(\reg_module/_09213_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16903_  (.A(\reg_module/_09164_ ),
    .X(\reg_module/_09214_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16904_  (.A1(\reg_module/_09211_ ),
    .A2(\reg_module/_09213_ ),
    .B1(\reg_module/_09214_ ),
    .Y(\reg_module/_00354_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16905_  (.A(\reg_module/_09202_ ),
    .B(net2065),
    .Y(\reg_module/_09215_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16906_  (.A(\reg_module/_08039_ ),
    .B(\reg_module/_09205_ ),
    .Y(\reg_module/_09216_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16907_  (.A(\reg_module/_09204_ ),
    .B(\reg_module/_09216_ ),
    .Y(\reg_module/_09217_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16908_  (.A1(\reg_module/_09215_ ),
    .A2(\reg_module/_09217_ ),
    .B1(\reg_module/_09214_ ),
    .Y(\reg_module/_00355_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16909_  (.A(\reg_module/_09202_ ),
    .B(net1410),
    .Y(\reg_module/_09218_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16910_  (.A(\reg_module/_08043_ ),
    .B(\reg_module/_09205_ ),
    .Y(\reg_module/_09219_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16911_  (.A(\reg_module/_09204_ ),
    .B(\reg_module/_09219_ ),
    .Y(\reg_module/_09220_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16912_  (.A1(\reg_module/_09218_ ),
    .A2(\reg_module/_09220_ ),
    .B1(\reg_module/_09214_ ),
    .Y(\reg_module/_00356_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16913_  (.A(\reg_module/_09202_ ),
    .B(net1683),
    .Y(\reg_module/_09221_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16914_  (.A(\reg_module/_08047_ ),
    .B(\reg_module/_09205_ ),
    .Y(\reg_module/_09222_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16915_  (.A(\reg_module/_09204_ ),
    .B(\reg_module/_09222_ ),
    .Y(\reg_module/_09223_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16916_  (.A1(\reg_module/_09221_ ),
    .A2(\reg_module/_09223_ ),
    .B1(\reg_module/_09214_ ),
    .Y(\reg_module/_00357_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16917_  (.A(\reg_module/_09201_ ),
    .X(\reg_module/_09224_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16918_  (.A(\reg_module/_09224_ ),
    .B(net1514),
    .Y(\reg_module/_09225_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16919_  (.A(\reg_module/_08873_ ),
    .X(\reg_module/_09226_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_16920_  (.A(\reg_module/_08953_ ),
    .X(\reg_module/_09227_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16921_  (.A(\reg_module/_08053_ ),
    .B(\reg_module/_09227_ ),
    .Y(\reg_module/_09228_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16922_  (.A(\reg_module/_09226_ ),
    .B(\reg_module/_09228_ ),
    .Y(\reg_module/_09229_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16923_  (.A1(\reg_module/_09225_ ),
    .A2(\reg_module/_09229_ ),
    .B1(\reg_module/_09214_ ),
    .Y(\reg_module/_00358_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16924_  (.A(\reg_module/_09224_ ),
    .B(net1447),
    .Y(\reg_module/_09230_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16925_  (.A(\reg_module/_08057_ ),
    .B(\reg_module/_09227_ ),
    .Y(\reg_module/_09231_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16926_  (.A(\reg_module/_09226_ ),
    .B(\reg_module/_09231_ ),
    .Y(\reg_module/_09232_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16927_  (.A1(\reg_module/_09230_ ),
    .A2(\reg_module/_09232_ ),
    .B1(\reg_module/_09214_ ),
    .Y(\reg_module/_00359_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16928_  (.A(\reg_module/_09224_ ),
    .B(net1900),
    .Y(\reg_module/_09233_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16929_  (.A(\reg_module/_08062_ ),
    .B(\reg_module/_09227_ ),
    .Y(\reg_module/_09234_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16930_  (.A(\reg_module/_09226_ ),
    .B(\reg_module/_09234_ ),
    .Y(\reg_module/_09235_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16931_  (.A(\reg_module/_09164_ ),
    .X(\reg_module/_09236_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16932_  (.A1(\reg_module/_09233_ ),
    .A2(\reg_module/_09235_ ),
    .B1(\reg_module/_09236_ ),
    .Y(\reg_module/_00360_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16933_  (.A(\reg_module/_09224_ ),
    .B(net1736),
    .Y(\reg_module/_09237_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16934_  (.A(\reg_module/_08068_ ),
    .B(\reg_module/_09227_ ),
    .Y(\reg_module/_09238_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16935_  (.A(\reg_module/_09226_ ),
    .B(\reg_module/_09238_ ),
    .Y(\reg_module/_09239_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16936_  (.A1(\reg_module/_09237_ ),
    .A2(\reg_module/_09239_ ),
    .B1(\reg_module/_09236_ ),
    .Y(\reg_module/_00361_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16937_  (.A(\reg_module/_09224_ ),
    .B(net1661),
    .Y(\reg_module/_09240_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16938_  (.A(\reg_module/_08072_ ),
    .B(\reg_module/_09227_ ),
    .Y(\reg_module/_09241_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16939_  (.A(\reg_module/_09226_ ),
    .B(\reg_module/_09241_ ),
    .Y(\reg_module/_09242_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16940_  (.A1(\reg_module/_09240_ ),
    .A2(\reg_module/_09242_ ),
    .B1(\reg_module/_09236_ ),
    .Y(\reg_module/_00362_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16941_  (.A(\reg_module/_09224_ ),
    .B(net1744),
    .Y(\reg_module/_09243_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16942_  (.A(\reg_module/_08076_ ),
    .B(\reg_module/_09227_ ),
    .Y(\reg_module/_09244_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16943_  (.A(\reg_module/_09226_ ),
    .B(\reg_module/_09244_ ),
    .Y(\reg_module/_09245_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16944_  (.A1(\reg_module/_09243_ ),
    .A2(\reg_module/_09245_ ),
    .B1(\reg_module/_09236_ ),
    .Y(\reg_module/_00363_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16945_  (.A(\reg_module/_09201_ ),
    .X(\reg_module/_09246_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16946_  (.A(\reg_module/_09246_ ),
    .B(net1532),
    .Y(\reg_module/_09247_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16947_  (.A(\reg_module/_08873_ ),
    .X(\reg_module/_09248_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_16948_  (.A(\reg_module/_08953_ ),
    .X(\reg_module/_09249_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16949_  (.A(\reg_module/_08082_ ),
    .B(\reg_module/_09249_ ),
    .Y(\reg_module/_09250_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16950_  (.A(\reg_module/_09248_ ),
    .B(\reg_module/_09250_ ),
    .Y(\reg_module/_09251_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16951_  (.A1(\reg_module/_09247_ ),
    .A2(\reg_module/_09251_ ),
    .B1(\reg_module/_09236_ ),
    .Y(\reg_module/_00364_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16952_  (.A(\reg_module/_09246_ ),
    .B(net1333),
    .Y(\reg_module/_09252_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16953_  (.A(\reg_module/_08086_ ),
    .B(\reg_module/_09249_ ),
    .Y(\reg_module/_09253_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16954_  (.A(\reg_module/_09248_ ),
    .B(\reg_module/_09253_ ),
    .Y(\reg_module/_09254_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16955_  (.A1(\reg_module/_09252_ ),
    .A2(\reg_module/_09254_ ),
    .B1(\reg_module/_09236_ ),
    .Y(\reg_module/_00365_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16956_  (.A(\reg_module/_09246_ ),
    .B(net1351),
    .Y(\reg_module/_09255_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16957_  (.A(\reg_module/_08091_ ),
    .B(\reg_module/_09249_ ),
    .Y(\reg_module/_09256_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16958_  (.A(\reg_module/_09248_ ),
    .B(\reg_module/_09256_ ),
    .Y(\reg_module/_09257_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_16959_  (.A(\reg_module/_09164_ ),
    .X(\reg_module/_09258_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16960_  (.A1(\reg_module/_09255_ ),
    .A2(\reg_module/_09257_ ),
    .B1(\reg_module/_09258_ ),
    .Y(\reg_module/_00366_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16961_  (.A(\reg_module/_09246_ ),
    .B(net1781),
    .Y(\reg_module/_09259_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16962_  (.A(\reg_module/_08096_ ),
    .B(\reg_module/_09249_ ),
    .Y(\reg_module/_09260_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16963_  (.A(\reg_module/_09248_ ),
    .B(\reg_module/_09260_ ),
    .Y(\reg_module/_09261_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16964_  (.A1(\reg_module/_09259_ ),
    .A2(\reg_module/_09261_ ),
    .B1(\reg_module/_09258_ ),
    .Y(\reg_module/_00367_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16965_  (.A(\reg_module/_09246_ ),
    .B(net2131),
    .Y(\reg_module/_09262_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16966_  (.A(\reg_module/_08101_ ),
    .B(\reg_module/_09249_ ),
    .Y(\reg_module/_09263_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16967_  (.A(\reg_module/_09248_ ),
    .B(\reg_module/_09263_ ),
    .Y(\reg_module/_09264_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16968_  (.A1(\reg_module/_09262_ ),
    .A2(\reg_module/_09264_ ),
    .B1(\reg_module/_09258_ ),
    .Y(\reg_module/_00368_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16969_  (.A(\reg_module/_09246_ ),
    .B(net2063),
    .Y(\reg_module/_09265_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16970_  (.A(\reg_module/_08105_ ),
    .B(\reg_module/_09249_ ),
    .Y(\reg_module/_09266_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16971_  (.A(\reg_module/_09248_ ),
    .B(\reg_module/_09266_ ),
    .Y(\reg_module/_09267_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16972_  (.A1(\reg_module/_09265_ ),
    .A2(\reg_module/_09267_ ),
    .B1(\reg_module/_09258_ ),
    .Y(\reg_module/_00369_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16973_  (.A(\reg_module/_09201_ ),
    .X(\reg_module/_09268_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16974_  (.A(\reg_module/_09268_ ),
    .B(net2040),
    .Y(\reg_module/_09269_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_16975_  (.A(\reg_module/_08183_ ),
    .X(\reg_module/_09270_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_16976_  (.A(\reg_module/_09270_ ),
    .X(\reg_module/_09271_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_16977_  (.A(\reg_module/_08953_ ),
    .X(\reg_module/_09272_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16978_  (.A(\reg_module/_08111_ ),
    .B(\reg_module/_09272_ ),
    .Y(\reg_module/_09273_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16979_  (.A(\reg_module/_09271_ ),
    .B(\reg_module/_09273_ ),
    .Y(\reg_module/_09274_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16980_  (.A1(\reg_module/_09269_ ),
    .A2(\reg_module/_09274_ ),
    .B1(\reg_module/_09258_ ),
    .Y(\reg_module/_00370_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16981_  (.A(\reg_module/_09268_ ),
    .B(net1871),
    .Y(\reg_module/_09275_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16982_  (.A(\reg_module/_08115_ ),
    .B(\reg_module/_09272_ ),
    .Y(\reg_module/_09276_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16983_  (.A(\reg_module/_09271_ ),
    .B(\reg_module/_09276_ ),
    .Y(\reg_module/_09277_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16984_  (.A1(\reg_module/_09275_ ),
    .A2(\reg_module/_09277_ ),
    .B1(\reg_module/_09258_ ),
    .Y(\reg_module/_00371_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16985_  (.A(\reg_module/_09268_ ),
    .B(net1598),
    .Y(\reg_module/_09278_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16986_  (.A(\reg_module/_08120_ ),
    .B(\reg_module/_09272_ ),
    .Y(\reg_module/_09279_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16987_  (.A(\reg_module/_09271_ ),
    .B(\reg_module/_09279_ ),
    .Y(\reg_module/_09280_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_16988_  (.A(\reg_module/_09164_ ),
    .X(\reg_module/_09281_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16989_  (.A1(\reg_module/_09278_ ),
    .A2(\reg_module/_09280_ ),
    .B1(\reg_module/_09281_ ),
    .Y(\reg_module/_00372_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16990_  (.A(\reg_module/_09268_ ),
    .B(net1537),
    .Y(\reg_module/_09282_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16991_  (.A(\reg_module/_08125_ ),
    .B(\reg_module/_09272_ ),
    .Y(\reg_module/_09283_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16992_  (.A(\reg_module/_09271_ ),
    .B(\reg_module/_09283_ ),
    .Y(\reg_module/_09284_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16993_  (.A1(\reg_module/_09282_ ),
    .A2(\reg_module/_09284_ ),
    .B1(\reg_module/_09281_ ),
    .Y(\reg_module/_00373_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16994_  (.A(\reg_module/_09268_ ),
    .B(net1365),
    .Y(\reg_module/_09285_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16995_  (.A(\reg_module/_08130_ ),
    .B(\reg_module/_09272_ ),
    .Y(\reg_module/_09286_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16996_  (.A(\reg_module/_09271_ ),
    .B(\reg_module/_09286_ ),
    .Y(\reg_module/_09287_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_16997_  (.A1(\reg_module/_09285_ ),
    .A2(\reg_module/_09287_ ),
    .B1(\reg_module/_09281_ ),
    .Y(\reg_module/_00374_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_16998_  (.A(\reg_module/_09268_ ),
    .B(net1314),
    .Y(\reg_module/_09288_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_16999_  (.A(\reg_module/_08134_ ),
    .B(\reg_module/_09272_ ),
    .Y(\reg_module/_09289_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17000_  (.A(\reg_module/_09271_ ),
    .B(\reg_module/_09289_ ),
    .Y(\reg_module/_09290_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17001_  (.A1(\reg_module/_09288_ ),
    .A2(\reg_module/_09290_ ),
    .B1(\reg_module/_09281_ ),
    .Y(\reg_module/_00375_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17002_  (.A(\reg_module/_09200_ ),
    .X(\reg_module/_09291_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17003_  (.A(\reg_module/_09291_ ),
    .B(net1620),
    .Y(\reg_module/_09292_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17004_  (.A(\reg_module/_09270_ ),
    .X(\reg_module/_09293_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17005_  (.A(\reg_module/_08953_ ),
    .X(\reg_module/_09294_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17006_  (.A(\reg_module/_08140_ ),
    .B(\reg_module/_09294_ ),
    .Y(\reg_module/_09295_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17007_  (.A(\reg_module/_09293_ ),
    .B(\reg_module/_09295_ ),
    .Y(\reg_module/_09296_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17008_  (.A1(\reg_module/_09292_ ),
    .A2(\reg_module/_09296_ ),
    .B1(\reg_module/_09281_ ),
    .Y(\reg_module/_00376_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17009_  (.A(\reg_module/_09291_ ),
    .B(net1259),
    .Y(\reg_module/_09297_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17010_  (.A(\reg_module/_08144_ ),
    .B(\reg_module/_09294_ ),
    .Y(\reg_module/_09298_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17011_  (.A(\reg_module/_09293_ ),
    .B(\reg_module/_09298_ ),
    .Y(\reg_module/_09299_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17012_  (.A1(\reg_module/_09297_ ),
    .A2(\reg_module/_09299_ ),
    .B1(\reg_module/_09281_ ),
    .Y(\reg_module/_00377_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17013_  (.A(\reg_module/_09291_ ),
    .B(net1319),
    .Y(\reg_module/_09300_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17014_  (.A(\reg_module/_08149_ ),
    .B(\reg_module/_09294_ ),
    .Y(\reg_module/_09301_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17015_  (.A(\reg_module/_09293_ ),
    .B(\reg_module/_09301_ ),
    .Y(\reg_module/_09302_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17016_  (.A(\reg_module/_07653_ ),
    .X(\reg_module/_09303_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_17017_  (.A(\reg_module/_09303_ ),
    .X(\reg_module/_09304_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17018_  (.A(\reg_module/_09304_ ),
    .X(\reg_module/_09305_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17019_  (.A1(\reg_module/_09300_ ),
    .A2(\reg_module/_09302_ ),
    .B1(\reg_module/_09305_ ),
    .Y(\reg_module/_00378_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17020_  (.A(\reg_module/_09291_ ),
    .B(net1238),
    .Y(\reg_module/_09306_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17021_  (.A(\reg_module/_08154_ ),
    .B(\reg_module/_09294_ ),
    .Y(\reg_module/_09307_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17022_  (.A(\reg_module/_09293_ ),
    .B(\reg_module/_09307_ ),
    .Y(\reg_module/_09308_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17023_  (.A1(\reg_module/_09306_ ),
    .A2(\reg_module/_09308_ ),
    .B1(\reg_module/_09305_ ),
    .Y(\reg_module/_00379_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17024_  (.A(\reg_module/_09291_ ),
    .B(net1328),
    .Y(\reg_module/_09309_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17025_  (.A(\reg_module/_08158_ ),
    .B(\reg_module/_09294_ ),
    .Y(\reg_module/_09310_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17026_  (.A(\reg_module/_09293_ ),
    .B(\reg_module/_09310_ ),
    .Y(\reg_module/_09311_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17027_  (.A1(\reg_module/_09309_ ),
    .A2(\reg_module/_09311_ ),
    .B1(\reg_module/_09305_ ),
    .Y(\reg_module/_00380_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17028_  (.A(\reg_module/_09291_ ),
    .B(net1262),
    .Y(\reg_module/_09312_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17029_  (.A(\reg_module/_08162_ ),
    .B(\reg_module/_09294_ ),
    .Y(\reg_module/_09313_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17030_  (.A(\reg_module/_09293_ ),
    .B(\reg_module/_09313_ ),
    .Y(\reg_module/_09314_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17031_  (.A1(\reg_module/_09312_ ),
    .A2(\reg_module/_09314_ ),
    .B1(\reg_module/_09305_ ),
    .Y(\reg_module/_00381_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17032_  (.A(\reg_module/_09201_ ),
    .B(net1230),
    .Y(\reg_module/_09315_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17033_  (.A(\reg_module/_09270_ ),
    .X(\reg_module/_09316_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17034_  (.A(\reg_module/_08166_ ),
    .B(\reg_module/_08954_ ),
    .Y(\reg_module/_09317_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17035_  (.A(\reg_module/_09316_ ),
    .B(\reg_module/_09317_ ),
    .Y(\reg_module/_09318_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17036_  (.A1(\reg_module/_09315_ ),
    .A2(\reg_module/_09318_ ),
    .B1(\reg_module/_09305_ ),
    .Y(\reg_module/_00382_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17037_  (.A(\reg_module/_09201_ ),
    .B(net1815),
    .Y(\reg_module/_09319_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17038_  (.A(\reg_module/_08170_ ),
    .B(\reg_module/_08954_ ),
    .Y(\reg_module/_09320_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17039_  (.A(\reg_module/_09316_ ),
    .B(\reg_module/_09320_ ),
    .Y(\reg_module/_09321_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17040_  (.A1(\reg_module/_09319_ ),
    .A2(\reg_module/_09321_ ),
    .B1(\reg_module/_09305_ ),
    .Y(\reg_module/_00383_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17041_  (.A(\reg_module/_08174_ ),
    .B(\reg_module/_07506_ ),
    .Y(\reg_module/_09322_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17042_  (.A(\reg_module/_09322_ ),
    .Y(\reg_module/_09323_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17043_  (.A(\reg_module/_07638_ ),
    .B(\reg_module/_09323_ ),
    .Y(\reg_module/_09324_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17044_  (.A(\reg_module/_09324_ ),
    .X(\reg_module/_09325_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17045_  (.A(\reg_module/_09325_ ),
    .X(\reg_module/_09326_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17046_  (.A(\reg_module/gprf[384] ),
    .Y(\reg_module/_09327_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17047_  (.A(\reg_module/_09326_ ),
    .B(\reg_module/_09327_ ),
    .Y(\reg_module/_09328_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17048_  (.A(\reg_module/_09328_ ),
    .Y(\reg_module/_09329_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17049_  (.A(\reg_module/_08663_ ),
    .X(\reg_module/_09330_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17050_  (.A(\reg_module/_09323_ ),
    .X(\reg_module/_09331_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17051_  (.A(\reg_module/_09331_ ),
    .X(\reg_module/_09332_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17052_  (.A(\reg_module/_09330_ ),
    .B(\reg_module/_07514_ ),
    .C(\reg_module/_09332_ ),
    .Y(\reg_module/_09333_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17053_  (.A(\reg_module/_09333_ ),
    .B(net1032),
    .Y(\reg_module/_09334_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17054_  (.A(\reg_module/_09329_ ),
    .B(\reg_module/_09334_ ),
    .Y(\reg_module/_00384_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17055_  (.A(\reg_module/gprf[385] ),
    .Y(\reg_module/_09335_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17056_  (.A(\reg_module/_09326_ ),
    .B(\reg_module/_09335_ ),
    .Y(\reg_module/_09336_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17057_  (.A(\reg_module/_09336_ ),
    .Y(\reg_module/_09337_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17058_  (.A(\reg_module/_09330_ ),
    .B(\reg_module/_07517_ ),
    .C(\reg_module/_09332_ ),
    .Y(\reg_module/_09338_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17059_  (.A(\reg_module/_09338_ ),
    .B(net1032),
    .Y(\reg_module/_09339_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17060_  (.A(\reg_module/_09337_ ),
    .B(\reg_module/_09339_ ),
    .Y(\reg_module/_00385_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17061_  (.A(\reg_module/gprf[386] ),
    .Y(\reg_module/_09340_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17062_  (.A(\reg_module/_09326_ ),
    .B(\reg_module/_09340_ ),
    .Y(\reg_module/_09341_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17063_  (.A(\reg_module/_09341_ ),
    .Y(\reg_module/_09342_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17064_  (.A(\reg_module/_09330_ ),
    .B(\reg_module/_07520_ ),
    .C(\reg_module/_09332_ ),
    .Y(\reg_module/_09343_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17065_  (.A(\reg_module/_09343_ ),
    .B(net1036),
    .Y(\reg_module/_09344_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17066_  (.A(\reg_module/_09342_ ),
    .B(\reg_module/_09344_ ),
    .Y(\reg_module/_00386_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17067_  (.A(\reg_module/gprf[387] ),
    .Y(\reg_module/_09345_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17068_  (.A(\reg_module/_09326_ ),
    .B(\reg_module/_09345_ ),
    .Y(\reg_module/_09346_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17069_  (.A(\reg_module/_09346_ ),
    .Y(\reg_module/_09347_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17070_  (.A(\reg_module/_09330_ ),
    .B(\reg_module/_07522_ ),
    .C(\reg_module/_09332_ ),
    .Y(\reg_module/_09348_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17071_  (.A(\reg_module/_09348_ ),
    .B(net1035),
    .Y(\reg_module/_09349_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17072_  (.A(\reg_module/_09347_ ),
    .B(\reg_module/_09349_ ),
    .Y(\reg_module/_00387_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17073_  (.A(\reg_module/gprf[388] ),
    .Y(\reg_module/_09350_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17074_  (.A(\reg_module/_09326_ ),
    .B(\reg_module/_09350_ ),
    .Y(\reg_module/_09351_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17075_  (.A(\reg_module/_09351_ ),
    .Y(\reg_module/_09352_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17076_  (.A(\reg_module/_09330_ ),
    .B(\reg_module/_07528_ ),
    .C(\reg_module/_09332_ ),
    .Y(\reg_module/_09353_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17077_  (.A(\reg_module/_09353_ ),
    .B(net1035),
    .Y(\reg_module/_09354_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17078_  (.A(\reg_module/_09352_ ),
    .B(\reg_module/_09354_ ),
    .Y(\reg_module/_00388_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17079_  (.A(\reg_module/gprf[389] ),
    .Y(\reg_module/_09355_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17080_  (.A(\reg_module/_09326_ ),
    .B(\reg_module/_09355_ ),
    .Y(\reg_module/_09356_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17081_  (.A(\reg_module/_09356_ ),
    .Y(\reg_module/_09357_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17082_  (.A(\reg_module/_09330_ ),
    .B(\reg_module/_07531_ ),
    .C(\reg_module/_09332_ ),
    .Y(\reg_module/_09358_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17083_  (.A(\reg_module/_09358_ ),
    .B(net1035),
    .Y(\reg_module/_09359_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17084_  (.A(\reg_module/_09357_ ),
    .B(\reg_module/_09359_ ),
    .Y(\reg_module/_00389_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17085_  (.A(\reg_module/_09325_ ),
    .X(\reg_module/_09360_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17086_  (.A(net2164),
    .Y(\reg_module/_09361_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17087_  (.A(\reg_module/_09360_ ),
    .B(\reg_module/_09361_ ),
    .Y(\reg_module/_09362_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17088_  (.A(\reg_module/_09362_ ),
    .Y(\reg_module/_09363_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17089_  (.A(\reg_module/_08957_ ),
    .X(\reg_module/_09364_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17090_  (.A(\reg_module/_09331_ ),
    .X(\reg_module/_09365_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17091_  (.A(\reg_module/_09364_ ),
    .B(\reg_module/_07535_ ),
    .C(\reg_module/_09365_ ),
    .Y(\reg_module/_09366_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17092_  (.A(\reg_module/_09366_ ),
    .B(net1042),
    .Y(\reg_module/_09367_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17093_  (.A(\reg_module/_09363_ ),
    .B(\reg_module/_09367_ ),
    .Y(\reg_module/_00390_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17094_  (.A(net2176),
    .Y(\reg_module/_09368_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17095_  (.A(\reg_module/_09360_ ),
    .B(\reg_module/_09368_ ),
    .Y(\reg_module/_09369_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17096_  (.A(\reg_module/_09369_ ),
    .Y(\reg_module/_09370_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17097_  (.A(\reg_module/_09364_ ),
    .B(\reg_module/_07538_ ),
    .C(\reg_module/_09365_ ),
    .Y(\reg_module/_09371_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17098_  (.A(\reg_module/_09371_ ),
    .B(net1042),
    .Y(\reg_module/_09372_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17099_  (.A(\reg_module/_09370_ ),
    .B(\reg_module/_09372_ ),
    .Y(\reg_module/_00391_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17100_  (.A(net2160),
    .Y(\reg_module/_09373_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17101_  (.A(\reg_module/_09360_ ),
    .B(\reg_module/_09373_ ),
    .Y(\reg_module/_09374_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17102_  (.A(\reg_module/_09374_ ),
    .Y(\reg_module/_09375_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17103_  (.A(\reg_module/_09364_ ),
    .B(\reg_module/_07541_ ),
    .C(\reg_module/_09365_ ),
    .Y(\reg_module/_09376_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17104_  (.A(\reg_module/_09376_ ),
    .B(net1042),
    .Y(\reg_module/_09377_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17105_  (.A(\reg_module/_09375_ ),
    .B(\reg_module/_09377_ ),
    .Y(\reg_module/_00392_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17106_  (.A(net2168),
    .Y(\reg_module/_09378_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17107_  (.A(\reg_module/_09360_ ),
    .B(\reg_module/_09378_ ),
    .Y(\reg_module/_09379_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17108_  (.A(\reg_module/_09379_ ),
    .Y(\reg_module/_09380_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17109_  (.A(\reg_module/_09364_ ),
    .B(\reg_module/_07544_ ),
    .C(\reg_module/_09365_ ),
    .Y(\reg_module/_09381_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17110_  (.A(\reg_module/_09381_ ),
    .B(net1043),
    .Y(\reg_module/_09382_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17111_  (.A(\reg_module/_09380_ ),
    .B(\reg_module/_09382_ ),
    .Y(\reg_module/_00393_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17112_  (.A(net2161),
    .Y(\reg_module/_09383_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17113_  (.A(\reg_module/_09360_ ),
    .B(\reg_module/_09383_ ),
    .Y(\reg_module/_09384_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17114_  (.A(\reg_module/_09384_ ),
    .Y(\reg_module/_09385_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17115_  (.A(\reg_module/_09364_ ),
    .B(\reg_module/_07547_ ),
    .C(\reg_module/_09365_ ),
    .Y(\reg_module/_09386_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17116_  (.A(\reg_module/_09386_ ),
    .B(net1044),
    .Y(\reg_module/_09387_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17117_  (.A(\reg_module/_09385_ ),
    .B(\reg_module/_09387_ ),
    .Y(\reg_module/_00394_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17118_  (.A(net2200),
    .Y(\reg_module/_09388_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17119_  (.A(\reg_module/_09360_ ),
    .B(\reg_module/_09388_ ),
    .Y(\reg_module/_09389_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17120_  (.A(\reg_module/_09389_ ),
    .Y(\reg_module/_09390_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17121_  (.A(\reg_module/_09364_ ),
    .B(\reg_module/_07551_ ),
    .C(\reg_module/_09365_ ),
    .Y(\reg_module/_09391_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17122_  (.A(\reg_module/_09391_ ),
    .B(net1044),
    .Y(\reg_module/_09392_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17123_  (.A(\reg_module/_09390_ ),
    .B(\reg_module/_09392_ ),
    .Y(\reg_module/_00395_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17124_  (.A(\reg_module/_09325_ ),
    .X(\reg_module/_09393_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17125_  (.A(\reg_module/gprf[396] ),
    .Y(\reg_module/_09394_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17126_  (.A(\reg_module/_09393_ ),
    .B(\reg_module/_09394_ ),
    .Y(\reg_module/_09395_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17127_  (.A(\reg_module/_09395_ ),
    .Y(\reg_module/_09396_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17128_  (.A(\reg_module/_08957_ ),
    .X(\reg_module/_09397_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17129_  (.A(\reg_module/_09331_ ),
    .X(\reg_module/_09398_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17130_  (.A(\reg_module/_09397_ ),
    .B(\reg_module/_07555_ ),
    .C(\reg_module/_09398_ ),
    .Y(\reg_module/_09399_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17131_  (.A(\reg_module/_09399_ ),
    .B(net1059),
    .Y(\reg_module/_09400_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17132_  (.A(\reg_module/_09396_ ),
    .B(\reg_module/_09400_ ),
    .Y(\reg_module/_00396_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17133_  (.A(net2199),
    .Y(\reg_module/_09401_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17134_  (.A(\reg_module/_09393_ ),
    .B(\reg_module/_09401_ ),
    .Y(\reg_module/_09402_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17135_  (.A(\reg_module/_09402_ ),
    .Y(\reg_module/_09403_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17136_  (.A(\reg_module/_09397_ ),
    .B(\reg_module/_07557_ ),
    .C(\reg_module/_09398_ ),
    .Y(\reg_module/_09404_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17137_  (.A(\reg_module/_09404_ ),
    .B(net1059),
    .Y(\reg_module/_09405_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17138_  (.A(\reg_module/_09403_ ),
    .B(\reg_module/_09405_ ),
    .Y(\reg_module/_00397_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17139_  (.A(net2156),
    .Y(\reg_module/_09406_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17140_  (.A(\reg_module/_09393_ ),
    .B(\reg_module/_09406_ ),
    .Y(\reg_module/_09407_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17141_  (.A(\reg_module/_09407_ ),
    .Y(\reg_module/_09408_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17142_  (.A(\reg_module/_09397_ ),
    .B(\reg_module/_07561_ ),
    .C(\reg_module/_09398_ ),
    .Y(\reg_module/_09409_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17143_  (.A(\reg_module/_09409_ ),
    .B(net1059),
    .Y(\reg_module/_09410_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17144_  (.A(\reg_module/_09408_ ),
    .B(\reg_module/_09410_ ),
    .Y(\reg_module/_00398_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17145_  (.A(net2159),
    .Y(\reg_module/_09411_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17146_  (.A(\reg_module/_09393_ ),
    .B(\reg_module/_09411_ ),
    .Y(\reg_module/_09412_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17147_  (.A(\reg_module/_09412_ ),
    .Y(\reg_module/_09413_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17148_  (.A(\reg_module/_09397_ ),
    .B(\reg_module/_07564_ ),
    .C(\reg_module/_09398_ ),
    .Y(\reg_module/_09414_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17149_  (.A(\reg_module/_09414_ ),
    .B(net1059),
    .Y(\reg_module/_09415_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17150_  (.A(\reg_module/_09413_ ),
    .B(\reg_module/_09415_ ),
    .Y(\reg_module/_00399_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17151_  (.A(net2190),
    .Y(\reg_module/_09416_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17152_  (.A(\reg_module/_09393_ ),
    .B(\reg_module/_09416_ ),
    .Y(\reg_module/_09417_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17153_  (.A(\reg_module/_09417_ ),
    .Y(\reg_module/_09418_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17154_  (.A(\reg_module/_09397_ ),
    .B(\reg_module/_07568_ ),
    .C(\reg_module/_09398_ ),
    .Y(\reg_module/_09419_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17155_  (.A(\reg_module/_09419_ ),
    .B(net1059),
    .Y(\reg_module/_09420_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17156_  (.A(\reg_module/_09418_ ),
    .B(\reg_module/_09420_ ),
    .Y(\reg_module/_00400_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17157_  (.A(\reg_module/gprf[401] ),
    .Y(\reg_module/_09421_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17158_  (.A(\reg_module/_09393_ ),
    .B(\reg_module/_09421_ ),
    .Y(\reg_module/_09422_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17159_  (.A(\reg_module/_09422_ ),
    .Y(\reg_module/_09423_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17160_  (.A(\reg_module/_09397_ ),
    .B(\reg_module/_07571_ ),
    .C(\reg_module/_09398_ ),
    .Y(\reg_module/_09424_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17161_  (.A(\reg_module/_09424_ ),
    .B(net1060),
    .Y(\reg_module/_09425_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17162_  (.A(\reg_module/_09423_ ),
    .B(\reg_module/_09425_ ),
    .Y(\reg_module/_00401_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17163_  (.A(\reg_module/_09325_ ),
    .X(\reg_module/_09426_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17164_  (.A(\reg_module/gprf[402] ),
    .Y(\reg_module/_09427_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17165_  (.A(\reg_module/_09426_ ),
    .B(\reg_module/_09427_ ),
    .Y(\reg_module/_09428_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17166_  (.A(\reg_module/_09428_ ),
    .Y(\reg_module/_09429_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17167_  (.A(\reg_module/_08957_ ),
    .X(\reg_module/_09430_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_17168_  (.A(\reg_module/_09331_ ),
    .X(\reg_module/_09431_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17169_  (.A(\reg_module/_09430_ ),
    .B(\reg_module/_07574_ ),
    .C(\reg_module/_09431_ ),
    .Y(\reg_module/_09432_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17170_  (.A(\reg_module/_09432_ ),
    .B(net1024),
    .Y(\reg_module/_09433_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17171_  (.A(\reg_module/_09429_ ),
    .B(\reg_module/_09433_ ),
    .Y(\reg_module/_00402_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17172_  (.A(\reg_module/gprf[403] ),
    .Y(\reg_module/_09434_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17173_  (.A(\reg_module/_09426_ ),
    .B(\reg_module/_09434_ ),
    .Y(\reg_module/_09435_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17174_  (.A(\reg_module/_09435_ ),
    .Y(\reg_module/_09436_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17175_  (.A(\reg_module/_09430_ ),
    .B(\reg_module/_07578_ ),
    .C(\reg_module/_09431_ ),
    .Y(\reg_module/_09437_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17176_  (.A(\reg_module/_09437_ ),
    .B(net1024),
    .Y(\reg_module/_09438_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17177_  (.A(\reg_module/_09436_ ),
    .B(\reg_module/_09438_ ),
    .Y(\reg_module/_00403_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17178_  (.A(net2186),
    .Y(\reg_module/_09439_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17179_  (.A(\reg_module/_09426_ ),
    .B(\reg_module/_09439_ ),
    .Y(\reg_module/_09440_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17180_  (.A(\reg_module/_09440_ ),
    .Y(\reg_module/_09441_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17181_  (.A(\reg_module/_09430_ ),
    .B(\reg_module/_07581_ ),
    .C(\reg_module/_09431_ ),
    .Y(\reg_module/_09442_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17182_  (.A(\reg_module/_09442_ ),
    .B(net1025),
    .Y(\reg_module/_09443_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17183_  (.A(\reg_module/_09441_ ),
    .B(\reg_module/_09443_ ),
    .Y(\reg_module/_00404_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17184_  (.A(net2177),
    .Y(\reg_module/_09444_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17185_  (.A(\reg_module/_09426_ ),
    .B(\reg_module/_09444_ ),
    .Y(\reg_module/_09445_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17186_  (.A(\reg_module/_09445_ ),
    .Y(\reg_module/_09446_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17187_  (.A(\reg_module/_09430_ ),
    .B(\reg_module/_07584_ ),
    .C(\reg_module/_09431_ ),
    .Y(\reg_module/_09447_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17188_  (.A(\reg_module/_09447_ ),
    .B(net1025),
    .Y(\reg_module/_09448_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17189_  (.A(\reg_module/_09446_ ),
    .B(\reg_module/_09448_ ),
    .Y(\reg_module/_00405_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17190_  (.A(net2202),
    .Y(\reg_module/_09449_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17191_  (.A(\reg_module/_09426_ ),
    .B(\reg_module/_09449_ ),
    .Y(\reg_module/_09450_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17192_  (.A(\reg_module/_09450_ ),
    .Y(\reg_module/_09451_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17193_  (.A(\reg_module/_09430_ ),
    .B(\reg_module/_07588_ ),
    .C(\reg_module/_09431_ ),
    .Y(\reg_module/_09452_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17194_  (.A(\reg_module/_09452_ ),
    .B(net1025),
    .Y(\reg_module/_09453_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17195_  (.A(\reg_module/_09451_ ),
    .B(\reg_module/_09453_ ),
    .Y(\reg_module/_00406_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17196_  (.A(net2197),
    .Y(\reg_module/_09454_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17197_  (.A(\reg_module/_09426_ ),
    .B(\reg_module/_09454_ ),
    .Y(\reg_module/_09455_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17198_  (.A(\reg_module/_09455_ ),
    .Y(\reg_module/_09456_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17199_  (.A(\reg_module/_09430_ ),
    .B(\reg_module/_07590_ ),
    .C(\reg_module/_09431_ ),
    .Y(\reg_module/_09457_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17200_  (.A(\reg_module/_09457_ ),
    .B(net1025),
    .Y(\reg_module/_09458_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17201_  (.A(\reg_module/_09456_ ),
    .B(\reg_module/_09458_ ),
    .Y(\reg_module/_00407_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17202_  (.A(\reg_module/_09324_ ),
    .X(\reg_module/_09459_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17203_  (.A(\reg_module/gprf[408] ),
    .Y(\reg_module/_09460_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17204_  (.A(\reg_module/_09459_ ),
    .B(\reg_module/_09460_ ),
    .Y(\reg_module/_09461_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17205_  (.A(\reg_module/_09461_ ),
    .Y(\reg_module/_09462_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17206_  (.A(\reg_module/_08957_ ),
    .X(\reg_module/_09463_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17207_  (.A(\reg_module/_09323_ ),
    .X(\reg_module/_09464_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17208_  (.A(\reg_module/_09463_ ),
    .B(\reg_module/_07595_ ),
    .C(\reg_module/_09464_ ),
    .Y(\reg_module/_09465_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17209_  (.A(\reg_module/_09465_ ),
    .B(net1007),
    .Y(\reg_module/_09466_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17210_  (.A(\reg_module/_09462_ ),
    .B(\reg_module/_09466_ ),
    .Y(\reg_module/_00408_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17211_  (.A(\reg_module/gprf[409] ),
    .Y(\reg_module/_09467_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17212_  (.A(\reg_module/_09459_ ),
    .B(\reg_module/_09467_ ),
    .Y(\reg_module/_09468_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17213_  (.A(\reg_module/_09468_ ),
    .Y(\reg_module/_09469_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17214_  (.A(\reg_module/_09463_ ),
    .B(\reg_module/_07598_ ),
    .C(\reg_module/_09464_ ),
    .Y(\reg_module/_09470_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17215_  (.A(\reg_module/_09470_ ),
    .B(net1007),
    .Y(\reg_module/_09471_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17216_  (.A(\reg_module/_09469_ ),
    .B(\reg_module/_09471_ ),
    .Y(\reg_module/_00409_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17217_  (.A(\reg_module/gprf[410] ),
    .Y(\reg_module/_09472_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17218_  (.A(\reg_module/_09459_ ),
    .B(\reg_module/_09472_ ),
    .Y(\reg_module/_09473_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17219_  (.A(\reg_module/_09473_ ),
    .Y(\reg_module/_09474_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17220_  (.A(\reg_module/_09463_ ),
    .B(\reg_module/_07601_ ),
    .C(\reg_module/_09464_ ),
    .Y(\reg_module/_09475_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17221_  (.A(\reg_module/_09475_ ),
    .B(net1005),
    .Y(\reg_module/_09476_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17222_  (.A(\reg_module/_09474_ ),
    .B(\reg_module/_09476_ ),
    .Y(\reg_module/_00410_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17223_  (.A(net2213),
    .Y(\reg_module/_09477_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17224_  (.A(\reg_module/_09459_ ),
    .B(\reg_module/_09477_ ),
    .Y(\reg_module/_09478_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17225_  (.A(\reg_module/_09478_ ),
    .Y(\reg_module/_09479_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17226_  (.A(\reg_module/_09463_ ),
    .B(\reg_module/_07604_ ),
    .C(\reg_module/_09464_ ),
    .Y(\reg_module/_09480_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17227_  (.A(\reg_module/_09480_ ),
    .B(net1004),
    .Y(\reg_module/_09481_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17228_  (.A(\reg_module/_09479_ ),
    .B(\reg_module/_09481_ ),
    .Y(\reg_module/_00411_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17229_  (.A(net2180),
    .Y(\reg_module/_09482_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17230_  (.A(\reg_module/_09459_ ),
    .B(\reg_module/_09482_ ),
    .Y(\reg_module/_09483_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17231_  (.A(\reg_module/_09483_ ),
    .Y(\reg_module/_09484_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17232_  (.A(\reg_module/_09463_ ),
    .B(\reg_module/_07607_ ),
    .C(\reg_module/_09464_ ),
    .Y(\reg_module/_09485_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17233_  (.A(\reg_module/_09485_ ),
    .B(net1004),
    .Y(\reg_module/_09486_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17234_  (.A(\reg_module/_09484_ ),
    .B(\reg_module/_09486_ ),
    .Y(\reg_module/_00412_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17235_  (.A(\reg_module/gprf[413] ),
    .Y(\reg_module/_09487_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17236_  (.A(\reg_module/_09459_ ),
    .B(\reg_module/_09487_ ),
    .Y(\reg_module/_09488_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17237_  (.A(\reg_module/_09488_ ),
    .Y(\reg_module/_09489_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17238_  (.A(\reg_module/_09463_ ),
    .B(\reg_module/_07610_ ),
    .C(\reg_module/_09464_ ),
    .Y(\reg_module/_09490_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17239_  (.A(\reg_module/_09490_ ),
    .B(net1004),
    .Y(\reg_module/_09491_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17240_  (.A(\reg_module/_09489_ ),
    .B(\reg_module/_09491_ ),
    .Y(\reg_module/_00413_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17241_  (.A(net2212),
    .Y(\reg_module/_09492_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17242_  (.A(\reg_module/_09325_ ),
    .B(\reg_module/_09492_ ),
    .Y(\reg_module/_09493_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17243_  (.A(\reg_module/_09493_ ),
    .Y(\reg_module/_09494_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17244_  (.A(\reg_module/_08958_ ),
    .B(\reg_module/_07613_ ),
    .C(\reg_module/_09331_ ),
    .Y(\reg_module/_09495_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17245_  (.A(\reg_module/_09495_ ),
    .B(net1010),
    .Y(\reg_module/_09496_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17246_  (.A(\reg_module/_09494_ ),
    .B(\reg_module/_09496_ ),
    .Y(\reg_module/_00414_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17247_  (.A(\reg_module/gprf[415] ),
    .Y(\reg_module/_09497_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17248_  (.A(\reg_module/_09325_ ),
    .B(\reg_module/_09497_ ),
    .Y(\reg_module/_09498_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17249_  (.A(\reg_module/_09498_ ),
    .Y(\reg_module/_09499_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17250_  (.A(\reg_module/_08958_ ),
    .B(\reg_module/_07616_ ),
    .C(\reg_module/_09331_ ),
    .Y(\reg_module/_09500_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17251_  (.A(\reg_module/_09500_ ),
    .B(net1011),
    .Y(\reg_module/_09501_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17252_  (.A(\reg_module/_09499_ ),
    .B(\reg_module/_09501_ ),
    .Y(\reg_module/_00415_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17253_  (.A(net963),
    .B(\reg_module/_08358_ ),
    .Y(\reg_module/_09502_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17254_  (.A(\reg_module/_07619_ ),
    .B(\reg_module/_08825_ ),
    .C(\reg_module/_09502_ ),
    .Y(\reg_module/_09503_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_17255_  (.A(\reg_module/_09503_ ),
    .X(\reg_module/_09504_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17256_  (.A(\reg_module/_09504_ ),
    .X(\reg_module/_09505_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17257_  (.A(\reg_module/_09505_ ),
    .B(net1396),
    .Y(\reg_module/_09506_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17258_  (.A(\reg_module/_08369_ ),
    .B(\reg_module/_09185_ ),
    .Y(\reg_module/_09507_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17259_  (.A(\reg_module/_09132_ ),
    .X(\reg_module/_09508_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17260_  (.A(\reg_module/_09507_ ),
    .B(\reg_module/_09508_ ),
    .Y(\reg_module/_09509_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17261_  (.A(\reg_module/_09304_ ),
    .X(\reg_module/_09510_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17262_  (.A1(\reg_module/_09506_ ),
    .A2(\reg_module/_09509_ ),
    .B1(\reg_module/_09510_ ),
    .Y(\reg_module/_00416_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17263_  (.A(\reg_module/_09505_ ),
    .B(net1658),
    .Y(\reg_module/_09511_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17264_  (.A(\reg_module/_08375_ ),
    .B(\reg_module/_09185_ ),
    .Y(\reg_module/_09512_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17265_  (.A(\reg_module/_09512_ ),
    .B(\reg_module/_09508_ ),
    .Y(\reg_module/_09513_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17266_  (.A1(\reg_module/_09511_ ),
    .A2(\reg_module/_09513_ ),
    .B1(\reg_module/_09510_ ),
    .Y(\reg_module/_00417_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17267_  (.A(\reg_module/_09505_ ),
    .B(net1754),
    .Y(\reg_module/_09514_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17268_  (.A(\reg_module/_09184_ ),
    .X(\reg_module/_09515_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17269_  (.A(\reg_module/_08379_ ),
    .B(\reg_module/_09515_ ),
    .Y(\reg_module/_09516_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17270_  (.A(\reg_module/_09516_ ),
    .B(\reg_module/_09508_ ),
    .Y(\reg_module/_09517_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17271_  (.A1(\reg_module/_09514_ ),
    .A2(\reg_module/_09517_ ),
    .B1(\reg_module/_09510_ ),
    .Y(\reg_module/_00418_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17272_  (.A(\reg_module/_09505_ ),
    .B(net1699),
    .Y(\reg_module/_09518_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17273_  (.A(\reg_module/_08383_ ),
    .B(\reg_module/_09515_ ),
    .Y(\reg_module/_09519_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17274_  (.A(\reg_module/_09519_ ),
    .B(\reg_module/_09508_ ),
    .Y(\reg_module/_09520_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17275_  (.A1(\reg_module/_09518_ ),
    .A2(\reg_module/_09520_ ),
    .B1(\reg_module/_09510_ ),
    .Y(\reg_module/_00419_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17276_  (.A(\reg_module/_09505_ ),
    .B(net1613),
    .Y(\reg_module/_09521_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17277_  (.A(\reg_module/_08388_ ),
    .B(\reg_module/_09515_ ),
    .Y(\reg_module/_09522_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17278_  (.A(\reg_module/_09522_ ),
    .B(\reg_module/_09508_ ),
    .Y(\reg_module/_09523_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17279_  (.A1(\reg_module/_09521_ ),
    .A2(\reg_module/_09523_ ),
    .B1(\reg_module/_09510_ ),
    .Y(\reg_module/_00420_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17280_  (.A(\reg_module/_09505_ ),
    .B(net1903),
    .Y(\reg_module/_09524_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17281_  (.A(\reg_module/_08392_ ),
    .B(\reg_module/_09515_ ),
    .Y(\reg_module/_09525_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17282_  (.A(\reg_module/_09525_ ),
    .B(\reg_module/_09508_ ),
    .Y(\reg_module/_09526_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17283_  (.A1(\reg_module/_09524_ ),
    .A2(\reg_module/_09526_ ),
    .B1(\reg_module/_09510_ ),
    .Y(\reg_module/_00421_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17284_  (.A(\reg_module/_09504_ ),
    .X(\reg_module/_09527_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17285_  (.A(\reg_module/_09527_ ),
    .B(net1657),
    .Y(\reg_module/_09528_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17286_  (.A(\reg_module/_08399_ ),
    .B(\reg_module/_09515_ ),
    .Y(\reg_module/_09529_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17287_  (.A(\reg_module/_09132_ ),
    .X(\reg_module/_09530_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17288_  (.A(\reg_module/_09529_ ),
    .B(\reg_module/_09530_ ),
    .Y(\reg_module/_09531_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17289_  (.A(\reg_module/_09304_ ),
    .X(\reg_module/_09532_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17290_  (.A1(\reg_module/_09528_ ),
    .A2(\reg_module/_09531_ ),
    .B1(\reg_module/_09532_ ),
    .Y(\reg_module/_00422_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17291_  (.A(\reg_module/_09527_ ),
    .B(net1517),
    .Y(\reg_module/_09533_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17292_  (.A(\reg_module/_08404_ ),
    .B(\reg_module/_09515_ ),
    .Y(\reg_module/_09534_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17293_  (.A(\reg_module/_09534_ ),
    .B(\reg_module/_09530_ ),
    .Y(\reg_module/_09535_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17294_  (.A1(\reg_module/_09533_ ),
    .A2(\reg_module/_09535_ ),
    .B1(\reg_module/_09532_ ),
    .Y(\reg_module/_00423_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17295_  (.A(\reg_module/_09527_ ),
    .B(net1674),
    .Y(\reg_module/_09536_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17296_  (.A(\reg_module/_09184_ ),
    .X(\reg_module/_09537_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17297_  (.A(\reg_module/_08408_ ),
    .B(\reg_module/_09537_ ),
    .Y(\reg_module/_09538_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17298_  (.A(\reg_module/_09538_ ),
    .B(\reg_module/_09530_ ),
    .Y(\reg_module/_09539_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17299_  (.A1(\reg_module/_09536_ ),
    .A2(\reg_module/_09539_ ),
    .B1(\reg_module/_09532_ ),
    .Y(\reg_module/_00424_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17300_  (.A(\reg_module/_09527_ ),
    .B(net1290),
    .Y(\reg_module/_09540_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17301_  (.A(\reg_module/_08412_ ),
    .B(\reg_module/_09537_ ),
    .Y(\reg_module/_09541_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17302_  (.A(\reg_module/_09541_ ),
    .B(\reg_module/_09530_ ),
    .Y(\reg_module/_09542_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17303_  (.A1(\reg_module/_09540_ ),
    .A2(\reg_module/_09542_ ),
    .B1(\reg_module/_09532_ ),
    .Y(\reg_module/_00425_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17304_  (.A(\reg_module/_09527_ ),
    .B(net1245),
    .Y(\reg_module/_09543_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17305_  (.A(\reg_module/_08417_ ),
    .B(\reg_module/_09537_ ),
    .Y(\reg_module/_09544_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17306_  (.A(\reg_module/_09544_ ),
    .B(\reg_module/_09530_ ),
    .Y(\reg_module/_09545_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17307_  (.A1(\reg_module/_09543_ ),
    .A2(\reg_module/_09545_ ),
    .B1(\reg_module/_09532_ ),
    .Y(\reg_module/_00426_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17308_  (.A(\reg_module/_09527_ ),
    .B(net1783),
    .Y(\reg_module/_09546_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17309_  (.A(\reg_module/_08421_ ),
    .B(\reg_module/_09537_ ),
    .Y(\reg_module/_09547_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17310_  (.A(\reg_module/_09547_ ),
    .B(\reg_module/_09530_ ),
    .Y(\reg_module/_09548_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17311_  (.A1(\reg_module/_09546_ ),
    .A2(\reg_module/_09548_ ),
    .B1(\reg_module/_09532_ ),
    .Y(\reg_module/_00427_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17312_  (.A(\reg_module/_09504_ ),
    .X(\reg_module/_09549_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17313_  (.A(\reg_module/_09549_ ),
    .B(net1345),
    .Y(\reg_module/_09550_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17314_  (.A(\reg_module/_08428_ ),
    .B(\reg_module/_09537_ ),
    .Y(\reg_module/_09551_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17315_  (.A(\reg_module/_09132_ ),
    .X(\reg_module/_09552_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17316_  (.A(\reg_module/_09551_ ),
    .B(\reg_module/_09552_ ),
    .Y(\reg_module/_09553_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17317_  (.A(\reg_module/_09304_ ),
    .X(\reg_module/_09554_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17318_  (.A1(\reg_module/_09550_ ),
    .A2(\reg_module/_09553_ ),
    .B1(\reg_module/_09554_ ),
    .Y(\reg_module/_00428_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17319_  (.A(\reg_module/_09549_ ),
    .B(net1229),
    .Y(\reg_module/_09555_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17320_  (.A(\reg_module/_08433_ ),
    .B(\reg_module/_09537_ ),
    .Y(\reg_module/_09556_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17321_  (.A(\reg_module/_09556_ ),
    .B(\reg_module/_09552_ ),
    .Y(\reg_module/_09557_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17322_  (.A1(\reg_module/_09555_ ),
    .A2(\reg_module/_09557_ ),
    .B1(\reg_module/_09554_ ),
    .Y(\reg_module/_00429_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17323_  (.A(\reg_module/_09549_ ),
    .B(net1285),
    .Y(\reg_module/_09558_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17324_  (.A(\reg_module/_09184_ ),
    .X(\reg_module/_09559_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17325_  (.A(\reg_module/_08437_ ),
    .B(\reg_module/_09559_ ),
    .Y(\reg_module/_09560_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17326_  (.A(\reg_module/_09560_ ),
    .B(\reg_module/_09552_ ),
    .Y(\reg_module/_09561_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17327_  (.A1(\reg_module/_09558_ ),
    .A2(\reg_module/_09561_ ),
    .B1(\reg_module/_09554_ ),
    .Y(\reg_module/_00430_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17328_  (.A(\reg_module/_09549_ ),
    .B(net1279),
    .Y(\reg_module/_09562_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17329_  (.A(\reg_module/_08441_ ),
    .B(\reg_module/_09559_ ),
    .Y(\reg_module/_09563_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17330_  (.A(\reg_module/_09563_ ),
    .B(\reg_module/_09552_ ),
    .Y(\reg_module/_09564_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17331_  (.A1(\reg_module/_09562_ ),
    .A2(\reg_module/_09564_ ),
    .B1(\reg_module/_09554_ ),
    .Y(\reg_module/_00431_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17332_  (.A(\reg_module/_09549_ ),
    .B(net1359),
    .Y(\reg_module/_09565_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17333_  (.A(\reg_module/_08446_ ),
    .B(\reg_module/_09559_ ),
    .Y(\reg_module/_09566_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17334_  (.A(\reg_module/_09566_ ),
    .B(\reg_module/_09552_ ),
    .Y(\reg_module/_09567_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17335_  (.A1(\reg_module/_09565_ ),
    .A2(\reg_module/_09567_ ),
    .B1(\reg_module/_09554_ ),
    .Y(\reg_module/_00432_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17336_  (.A(\reg_module/_09549_ ),
    .B(net1363),
    .Y(\reg_module/_09568_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17337_  (.A(\reg_module/_08450_ ),
    .B(\reg_module/_09559_ ),
    .Y(\reg_module/_09569_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17338_  (.A(\reg_module/_09569_ ),
    .B(\reg_module/_09552_ ),
    .Y(\reg_module/_09570_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17339_  (.A1(\reg_module/_09568_ ),
    .A2(\reg_module/_09570_ ),
    .B1(\reg_module/_09554_ ),
    .Y(\reg_module/_00433_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17340_  (.A(\reg_module/_09504_ ),
    .X(\reg_module/_09571_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17341_  (.A(\reg_module/_09571_ ),
    .B(net2089),
    .Y(\reg_module/_09572_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17342_  (.A(\reg_module/_08457_ ),
    .B(\reg_module/_09559_ ),
    .Y(\reg_module/_09573_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17343_  (.A(\reg_module/_07640_ ),
    .X(\reg_module/_09574_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17344_  (.A(\reg_module/_09573_ ),
    .B(\reg_module/_09574_ ),
    .Y(\reg_module/_09575_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17345_  (.A(\reg_module/_09304_ ),
    .X(\reg_module/_09576_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17346_  (.A1(\reg_module/_09572_ ),
    .A2(\reg_module/_09575_ ),
    .B1(\reg_module/_09576_ ),
    .Y(\reg_module/_00434_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17347_  (.A(\reg_module/_09571_ ),
    .B(\reg_module/gprf[435] ),
    .Y(\reg_module/_09577_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17348_  (.A(\reg_module/_08462_ ),
    .B(\reg_module/_09559_ ),
    .Y(\reg_module/_09578_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17349_  (.A(\reg_module/_09578_ ),
    .B(\reg_module/_09574_ ),
    .Y(\reg_module/_09579_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17350_  (.A1(\reg_module/_09577_ ),
    .A2(\reg_module/_09579_ ),
    .B1(\reg_module/_09576_ ),
    .Y(\reg_module/_00435_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17351_  (.A(\reg_module/_09571_ ),
    .B(net1495),
    .Y(\reg_module/_09580_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17352_  (.A(\reg_module/_09184_ ),
    .X(\reg_module/_09581_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17353_  (.A(\reg_module/_08466_ ),
    .B(\reg_module/_09581_ ),
    .Y(\reg_module/_09582_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17354_  (.A(\reg_module/_09582_ ),
    .B(\reg_module/_09574_ ),
    .Y(\reg_module/_09583_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17355_  (.A1(\reg_module/_09580_ ),
    .A2(\reg_module/_09583_ ),
    .B1(\reg_module/_09576_ ),
    .Y(\reg_module/_00436_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17356_  (.A(\reg_module/_09571_ ),
    .B(net1411),
    .Y(\reg_module/_09584_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17357_  (.A(\reg_module/_08470_ ),
    .B(\reg_module/_09581_ ),
    .Y(\reg_module/_09585_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17358_  (.A(\reg_module/_09585_ ),
    .B(\reg_module/_09574_ ),
    .Y(\reg_module/_09586_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17359_  (.A1(\reg_module/_09584_ ),
    .A2(\reg_module/_09586_ ),
    .B1(\reg_module/_09576_ ),
    .Y(\reg_module/_00437_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17360_  (.A(\reg_module/_09571_ ),
    .B(net1408),
    .Y(\reg_module/_09587_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17361_  (.A(\reg_module/_08475_ ),
    .B(\reg_module/_09581_ ),
    .Y(\reg_module/_09588_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17362_  (.A(\reg_module/_09588_ ),
    .B(\reg_module/_09574_ ),
    .Y(\reg_module/_09589_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17363_  (.A1(\reg_module/_09587_ ),
    .A2(\reg_module/_09589_ ),
    .B1(\reg_module/_09576_ ),
    .Y(\reg_module/_00438_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17364_  (.A(\reg_module/_09571_ ),
    .B(net1564),
    .Y(\reg_module/_09590_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17365_  (.A(\reg_module/_08479_ ),
    .B(\reg_module/_09581_ ),
    .Y(\reg_module/_09591_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17366_  (.A(\reg_module/_09591_ ),
    .B(\reg_module/_09574_ ),
    .Y(\reg_module/_09592_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17367_  (.A1(\reg_module/_09590_ ),
    .A2(\reg_module/_09592_ ),
    .B1(\reg_module/_09576_ ),
    .Y(\reg_module/_00439_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17368_  (.A(\reg_module/_09503_ ),
    .X(\reg_module/_09593_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17369_  (.A(\reg_module/_09593_ ),
    .B(net1753),
    .Y(\reg_module/_09594_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17370_  (.A(\reg_module/_08486_ ),
    .B(\reg_module/_09581_ ),
    .Y(\reg_module/_09595_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17371_  (.A(\reg_module/_07640_ ),
    .X(\reg_module/_09596_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17372_  (.A(\reg_module/_09595_ ),
    .B(\reg_module/_09596_ ),
    .Y(\reg_module/_09597_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17373_  (.A(\reg_module/_09304_ ),
    .X(\reg_module/_09598_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17374_  (.A1(\reg_module/_09594_ ),
    .A2(\reg_module/_09597_ ),
    .B1(\reg_module/_09598_ ),
    .Y(\reg_module/_00440_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17375_  (.A(\reg_module/_09593_ ),
    .B(net1566),
    .Y(\reg_module/_09599_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17376_  (.A(\reg_module/_08491_ ),
    .B(\reg_module/_09581_ ),
    .Y(\reg_module/_09600_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17377_  (.A(\reg_module/_09600_ ),
    .B(\reg_module/_09596_ ),
    .Y(\reg_module/_09601_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17378_  (.A1(\reg_module/_09599_ ),
    .A2(\reg_module/_09601_ ),
    .B1(\reg_module/_09598_ ),
    .Y(\reg_module/_00441_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17379_  (.A(\reg_module/_09593_ ),
    .B(net1231),
    .Y(\reg_module/_09602_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_17380_  (.A(\reg_module/_09184_ ),
    .X(\reg_module/_09603_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17381_  (.A(\reg_module/_08495_ ),
    .B(\reg_module/_09603_ ),
    .Y(\reg_module/_09604_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17382_  (.A(\reg_module/_09604_ ),
    .B(\reg_module/_09596_ ),
    .Y(\reg_module/_09605_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17383_  (.A1(\reg_module/_09602_ ),
    .A2(\reg_module/_09605_ ),
    .B1(\reg_module/_09598_ ),
    .Y(\reg_module/_00442_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17384_  (.A(\reg_module/_09593_ ),
    .B(net1236),
    .Y(\reg_module/_09606_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17385_  (.A(\reg_module/_08499_ ),
    .B(\reg_module/_09603_ ),
    .Y(\reg_module/_09607_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17386_  (.A(\reg_module/_09607_ ),
    .B(\reg_module/_09596_ ),
    .Y(\reg_module/_09608_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17387_  (.A1(\reg_module/_09606_ ),
    .A2(\reg_module/_09608_ ),
    .B1(\reg_module/_09598_ ),
    .Y(\reg_module/_00443_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17388_  (.A(\reg_module/_09593_ ),
    .B(net1249),
    .Y(\reg_module/_09609_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17389_  (.A(\reg_module/_08504_ ),
    .B(\reg_module/_09603_ ),
    .Y(\reg_module/_09610_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17390_  (.A(\reg_module/_09610_ ),
    .B(\reg_module/_09596_ ),
    .Y(\reg_module/_09611_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17391_  (.A1(\reg_module/_09609_ ),
    .A2(\reg_module/_09611_ ),
    .B1(\reg_module/_09598_ ),
    .Y(\reg_module/_00444_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17392_  (.A(\reg_module/_09593_ ),
    .B(net1588),
    .Y(\reg_module/_09612_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17393_  (.A(\reg_module/_08508_ ),
    .B(\reg_module/_09603_ ),
    .Y(\reg_module/_09613_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17394_  (.A(\reg_module/_09613_ ),
    .B(\reg_module/_09596_ ),
    .Y(\reg_module/_09614_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17395_  (.A1(\reg_module/_09612_ ),
    .A2(\reg_module/_09614_ ),
    .B1(\reg_module/_09598_ ),
    .Y(\reg_module/_00445_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17396_  (.A(\reg_module/_09504_ ),
    .B(net1468),
    .Y(\reg_module/_09615_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17397_  (.A(\reg_module/_08513_ ),
    .B(\reg_module/_09603_ ),
    .Y(\reg_module/_09616_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17398_  (.A(\reg_module/_09616_ ),
    .B(\reg_module/_07641_ ),
    .Y(\reg_module/_09617_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_17399_  (.A(\reg_module/_09303_ ),
    .X(\reg_module/_09618_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17400_  (.A(\reg_module/_09618_ ),
    .X(\reg_module/_09619_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17401_  (.A1(\reg_module/_09615_ ),
    .A2(\reg_module/_09617_ ),
    .B1(\reg_module/_09619_ ),
    .Y(\reg_module/_00446_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17402_  (.A(\reg_module/_09504_ ),
    .B(net1250),
    .Y(\reg_module/_09620_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17403_  (.A(\reg_module/_08518_ ),
    .B(\reg_module/_09603_ ),
    .Y(\reg_module/_09621_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17404_  (.A(\reg_module/_09621_ ),
    .B(\reg_module/_07641_ ),
    .Y(\reg_module/_09622_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17405_  (.A1(\reg_module/_09620_ ),
    .A2(\reg_module/_09622_ ),
    .B1(\reg_module/_09619_ ),
    .Y(\reg_module/_00447_ ));
 sky130_fd_sc_hd__and3_1 \reg_module/_17406_  (.A(\reg_module/_07808_ ),
    .B(\reg_module/_07625_ ),
    .C(\reg_module/_07817_ ),
    .X(\reg_module/_09623_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17407_  (.A(\reg_module/_07619_ ),
    .B(\reg_module/_08825_ ),
    .C(\reg_module/_09623_ ),
    .Y(\reg_module/_09624_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_17408_  (.A(\reg_module/_09624_ ),
    .X(\reg_module/_09625_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17409_  (.A(\reg_module/_09625_ ),
    .X(\reg_module/_09626_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17410_  (.A(\reg_module/_09626_ ),
    .B(net1409),
    .Y(\reg_module/_09627_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17411_  (.A(net967),
    .B(net977),
    .C(\reg_module/_07821_ ),
    .Y(\reg_module/_09628_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17412_  (.A(\reg_module/_09316_ ),
    .B(\reg_module/_09628_ ),
    .Y(\reg_module/_09629_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17413_  (.A1(\reg_module/_09627_ ),
    .A2(\reg_module/_09629_ ),
    .B1(\reg_module/_09619_ ),
    .Y(\reg_module/_00448_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17414_  (.A(\reg_module/_09626_ ),
    .B(net1252),
    .Y(\reg_module/_09630_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17415_  (.A(net968),
    .B(net980),
    .C(\reg_module/_07826_ ),
    .Y(\reg_module/_09631_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17416_  (.A(\reg_module/_09316_ ),
    .B(\reg_module/_09631_ ),
    .Y(\reg_module/_09632_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17417_  (.A1(\reg_module/_09630_ ),
    .A2(\reg_module/_09632_ ),
    .B1(\reg_module/_09619_ ),
    .Y(\reg_module/_00449_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17418_  (.A(\reg_module/_09626_ ),
    .B(net1729),
    .Y(\reg_module/_09633_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17419_  (.A(net968),
    .B(net981),
    .C(\reg_module/_07831_ ),
    .Y(\reg_module/_09634_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17420_  (.A(\reg_module/_09316_ ),
    .B(\reg_module/_09634_ ),
    .Y(\reg_module/_09635_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17421_  (.A1(\reg_module/_09633_ ),
    .A2(\reg_module/_09635_ ),
    .B1(\reg_module/_09619_ ),
    .Y(\reg_module/_00450_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17422_  (.A(\reg_module/_09626_ ),
    .B(net1776),
    .Y(\reg_module/_09636_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17423_  (.A(net968),
    .B(net981),
    .C(\reg_module/_07836_ ),
    .Y(\reg_module/_09637_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17424_  (.A(\reg_module/_09316_ ),
    .B(\reg_module/_09637_ ),
    .Y(\reg_module/_09638_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17425_  (.A1(\reg_module/_09636_ ),
    .A2(\reg_module/_09638_ ),
    .B1(\reg_module/_09619_ ),
    .Y(\reg_module/_00451_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17426_  (.A(\reg_module/_09626_ ),
    .B(net1649),
    .Y(\reg_module/_09639_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17427_  (.A(\reg_module/_09270_ ),
    .X(\reg_module/_09640_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17428_  (.A(net968),
    .B(net981),
    .C(\reg_module/_07844_ ),
    .Y(\reg_module/_09641_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17429_  (.A(\reg_module/_09640_ ),
    .B(\reg_module/_09641_ ),
    .Y(\reg_module/_09642_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17430_  (.A(\reg_module/_09618_ ),
    .X(\reg_module/_09643_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17431_  (.A1(\reg_module/_09639_ ),
    .A2(\reg_module/_09642_ ),
    .B1(\reg_module/_09643_ ),
    .Y(\reg_module/_00452_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17432_  (.A(\reg_module/_09626_ ),
    .B(net1548),
    .Y(\reg_module/_09644_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17433_  (.A(net968),
    .B(net981),
    .C(\reg_module/_07850_ ),
    .Y(\reg_module/_09645_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17434_  (.A(\reg_module/_09640_ ),
    .B(\reg_module/_09645_ ),
    .Y(\reg_module/_09646_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17435_  (.A1(\reg_module/_09644_ ),
    .A2(\reg_module/_09646_ ),
    .B1(\reg_module/_09643_ ),
    .Y(\reg_module/_00453_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17436_  (.A(\reg_module/_09625_ ),
    .X(\reg_module/_09647_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17437_  (.A(\reg_module/_09647_ ),
    .B(net1451),
    .Y(\reg_module/_09648_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17438_  (.A(net968),
    .B(net982),
    .C(\reg_module/_07858_ ),
    .Y(\reg_module/_09649_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17439_  (.A(\reg_module/_09640_ ),
    .B(\reg_module/_09649_ ),
    .Y(\reg_module/_09650_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17440_  (.A1(\reg_module/_09648_ ),
    .A2(\reg_module/_09650_ ),
    .B1(\reg_module/_09643_ ),
    .Y(\reg_module/_00454_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17441_  (.A(\reg_module/_09647_ ),
    .B(net1480),
    .Y(\reg_module/_09651_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17442_  (.A(net969),
    .B(net982),
    .C(\reg_module/_07863_ ),
    .Y(\reg_module/_09652_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17443_  (.A(\reg_module/_09640_ ),
    .B(\reg_module/_09652_ ),
    .Y(\reg_module/_09653_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17444_  (.A1(\reg_module/_09651_ ),
    .A2(\reg_module/_09653_ ),
    .B1(\reg_module/_09643_ ),
    .Y(\reg_module/_00455_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17445_  (.A(\reg_module/_09647_ ),
    .B(net1398),
    .Y(\reg_module/_09654_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17446_  (.A(net969),
    .B(net982),
    .C(\reg_module/_07868_ ),
    .Y(\reg_module/_09655_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17447_  (.A(\reg_module/_09640_ ),
    .B(\reg_module/_09655_ ),
    .Y(\reg_module/_09656_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17448_  (.A1(\reg_module/_09654_ ),
    .A2(\reg_module/_09656_ ),
    .B1(\reg_module/_09643_ ),
    .Y(\reg_module/_00456_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17449_  (.A(\reg_module/_09647_ ),
    .B(net1615),
    .Y(\reg_module/_09657_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17450_  (.A(net969),
    .B(net983),
    .C(\reg_module/_07873_ ),
    .Y(\reg_module/_09658_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17451_  (.A(\reg_module/_09640_ ),
    .B(\reg_module/_09658_ ),
    .Y(\reg_module/_09659_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17452_  (.A1(\reg_module/_09657_ ),
    .A2(\reg_module/_09659_ ),
    .B1(\reg_module/_09643_ ),
    .Y(\reg_module/_00457_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17453_  (.A(\reg_module/_09647_ ),
    .B(net1540),
    .Y(\reg_module/_09660_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17454_  (.A(\reg_module/_09270_ ),
    .X(\reg_module/_09661_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17455_  (.A(net973),
    .B(net989),
    .C(\reg_module/_07880_ ),
    .Y(\reg_module/_09662_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17456_  (.A(\reg_module/_09661_ ),
    .B(\reg_module/_09662_ ),
    .Y(\reg_module/_09663_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17457_  (.A(\reg_module/_09618_ ),
    .X(\reg_module/_09664_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17458_  (.A1(\reg_module/_09660_ ),
    .A2(\reg_module/_09663_ ),
    .B1(\reg_module/_09664_ ),
    .Y(\reg_module/_00458_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17459_  (.A(\reg_module/_09647_ ),
    .B(net1479),
    .Y(\reg_module/_09665_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17460_  (.A(net973),
    .B(net989),
    .C(\reg_module/_07886_ ),
    .Y(\reg_module/_09666_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17461_  (.A(\reg_module/_09661_ ),
    .B(\reg_module/_09666_ ),
    .Y(\reg_module/_09667_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17462_  (.A1(\reg_module/_09665_ ),
    .A2(\reg_module/_09667_ ),
    .B1(\reg_module/_09664_ ),
    .Y(\reg_module/_00459_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17463_  (.A(\reg_module/_09625_ ),
    .X(\reg_module/_09668_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17464_  (.A(\reg_module/_09668_ ),
    .B(net1488),
    .Y(\reg_module/_09669_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17465_  (.A(net973),
    .B(net988),
    .C(\reg_module/_07894_ ),
    .Y(\reg_module/_09670_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17466_  (.A(\reg_module/_09661_ ),
    .B(\reg_module/_09670_ ),
    .Y(\reg_module/_09671_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17467_  (.A1(\reg_module/_09669_ ),
    .A2(\reg_module/_09671_ ),
    .B1(\reg_module/_09664_ ),
    .Y(\reg_module/_00460_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17468_  (.A(\reg_module/_09668_ ),
    .B(net1417),
    .Y(\reg_module/_09672_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17469_  (.A(net973),
    .B(net992),
    .C(\reg_module/_07899_ ),
    .Y(\reg_module/_09673_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17470_  (.A(\reg_module/_09661_ ),
    .B(\reg_module/_09673_ ),
    .Y(\reg_module/_09674_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17471_  (.A1(\reg_module/_09672_ ),
    .A2(\reg_module/_09674_ ),
    .B1(\reg_module/_09664_ ),
    .Y(\reg_module/_00461_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17472_  (.A(\reg_module/_09668_ ),
    .B(net1725),
    .Y(\reg_module/_09675_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17473_  (.A(net973),
    .B(net991),
    .C(\reg_module/_07904_ ),
    .Y(\reg_module/_09676_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17474_  (.A(\reg_module/_09661_ ),
    .B(\reg_module/_09676_ ),
    .Y(\reg_module/_09677_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17475_  (.A1(\reg_module/_09675_ ),
    .A2(\reg_module/_09677_ ),
    .B1(\reg_module/_09664_ ),
    .Y(\reg_module/_00462_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17476_  (.A(\reg_module/_09668_ ),
    .B(net1664),
    .Y(\reg_module/_09678_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17477_  (.A(net974),
    .B(net991),
    .C(\reg_module/_07909_ ),
    .Y(\reg_module/_09679_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17478_  (.A(\reg_module/_09661_ ),
    .B(\reg_module/_09679_ ),
    .Y(\reg_module/_09680_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17479_  (.A1(\reg_module/_09678_ ),
    .A2(\reg_module/_09680_ ),
    .B1(\reg_module/_09664_ ),
    .Y(\reg_module/_00463_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17480_  (.A(\reg_module/_09668_ ),
    .B(net1586),
    .Y(\reg_module/_09681_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17481_  (.A(\reg_module/_09270_ ),
    .X(\reg_module/_09682_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17482_  (.A(net973),
    .B(net991),
    .C(\reg_module/_07916_ ),
    .Y(\reg_module/_09683_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17483_  (.A(\reg_module/_09682_ ),
    .B(\reg_module/_09683_ ),
    .Y(\reg_module/_09684_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17484_  (.A(\reg_module/_09618_ ),
    .X(\reg_module/_09685_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17485_  (.A1(\reg_module/_09681_ ),
    .A2(\reg_module/_09684_ ),
    .B1(\reg_module/_09685_ ),
    .Y(\reg_module/_00464_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17486_  (.A(\reg_module/_09668_ ),
    .B(net1593),
    .Y(\reg_module/_09686_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17487_  (.A(net975),
    .B(net991),
    .C(\reg_module/_07922_ ),
    .Y(\reg_module/_09687_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17488_  (.A(\reg_module/_09682_ ),
    .B(net280),
    .Y(\reg_module/_09688_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17489_  (.A1(\reg_module/_09686_ ),
    .A2(\reg_module/_09688_ ),
    .B1(\reg_module/_09685_ ),
    .Y(\reg_module/_00465_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17490_  (.A(\reg_module/_09625_ ),
    .X(\reg_module/_09689_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17491_  (.A(\reg_module/_09689_ ),
    .B(net1545),
    .Y(\reg_module/_09690_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17492_  (.A(net974),
    .B(net991),
    .C(\reg_module/_07930_ ),
    .Y(\reg_module/_09691_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17493_  (.A(\reg_module/_09682_ ),
    .B(\reg_module/_09691_ ),
    .Y(\reg_module/_09692_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17494_  (.A1(\reg_module/_09690_ ),
    .A2(\reg_module/_09692_ ),
    .B1(\reg_module/_09685_ ),
    .Y(\reg_module/_00466_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17495_  (.A(\reg_module/_09689_ ),
    .B(net1686),
    .Y(\reg_module/_09693_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17496_  (.A(net974),
    .B(net991),
    .C(\reg_module/_07935_ ),
    .Y(\reg_module/_09694_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17497_  (.A(\reg_module/_09682_ ),
    .B(\reg_module/_09694_ ),
    .Y(\reg_module/_09695_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17498_  (.A1(\reg_module/_09693_ ),
    .A2(\reg_module/_09695_ ),
    .B1(\reg_module/_09685_ ),
    .Y(\reg_module/_00467_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17499_  (.A(\reg_module/_09689_ ),
    .B(net1339),
    .Y(\reg_module/_09696_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17500_  (.A(net971),
    .B(net987),
    .C(\reg_module/_07940_ ),
    .Y(\reg_module/_09697_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17501_  (.A(\reg_module/_09682_ ),
    .B(\reg_module/_09697_ ),
    .Y(\reg_module/_09698_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17502_  (.A1(\reg_module/_09696_ ),
    .A2(\reg_module/_09698_ ),
    .B1(\reg_module/_09685_ ),
    .Y(\reg_module/_00468_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17503_  (.A(\reg_module/_09689_ ),
    .B(net1643),
    .Y(\reg_module/_09699_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17504_  (.A(net971),
    .B(net987),
    .C(\reg_module/_07945_ ),
    .Y(\reg_module/_09700_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17505_  (.A(\reg_module/_09682_ ),
    .B(\reg_module/_09700_ ),
    .Y(\reg_module/_09701_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17506_  (.A1(\reg_module/_09699_ ),
    .A2(\reg_module/_09701_ ),
    .B1(\reg_module/_09685_ ),
    .Y(\reg_module/_00469_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17507_  (.A(\reg_module/_09689_ ),
    .B(net1372),
    .Y(\reg_module/_09702_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_17508_  (.A(\reg_module/_08183_ ),
    .X(\reg_module/_09703_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17509_  (.A(\reg_module/_09703_ ),
    .X(\reg_module/_09704_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17510_  (.A(net971),
    .B(net985),
    .C(\reg_module/_07952_ ),
    .Y(\reg_module/_09705_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17511_  (.A(\reg_module/_09704_ ),
    .B(\reg_module/_09705_ ),
    .Y(\reg_module/_09706_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17512_  (.A(\reg_module/_09618_ ),
    .X(\reg_module/_09707_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17513_  (.A1(\reg_module/_09702_ ),
    .A2(\reg_module/_09706_ ),
    .B1(\reg_module/_09707_ ),
    .Y(\reg_module/_00470_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17514_  (.A(\reg_module/_09689_ ),
    .B(net1374),
    .Y(\reg_module/_09708_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17515_  (.A(net971),
    .B(net985),
    .C(\reg_module/_07958_ ),
    .Y(\reg_module/_09709_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17516_  (.A(\reg_module/_09704_ ),
    .B(\reg_module/_09709_ ),
    .Y(\reg_module/_09710_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17517_  (.A1(\reg_module/_09708_ ),
    .A2(\reg_module/_09710_ ),
    .B1(\reg_module/_09707_ ),
    .Y(\reg_module/_00471_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17518_  (.A(\reg_module/_09624_ ),
    .X(\reg_module/_09711_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17519_  (.A(\reg_module/_09711_ ),
    .B(net1254),
    .Y(\reg_module/_09712_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17520_  (.A(net971),
    .B(net985),
    .C(\reg_module/_07966_ ),
    .Y(\reg_module/_09713_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17521_  (.A(\reg_module/_09704_ ),
    .B(\reg_module/_09713_ ),
    .Y(\reg_module/_09714_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17522_  (.A1(\reg_module/_09712_ ),
    .A2(\reg_module/_09714_ ),
    .B1(\reg_module/_09707_ ),
    .Y(\reg_module/_00472_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17523_  (.A(\reg_module/_09711_ ),
    .B(net1394),
    .Y(\reg_module/_09715_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17524_  (.A(net971),
    .B(net985),
    .C(\reg_module/_07971_ ),
    .Y(\reg_module/_09716_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17525_  (.A(\reg_module/_09704_ ),
    .B(\reg_module/_09716_ ),
    .Y(\reg_module/_09717_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17526_  (.A1(\reg_module/_09715_ ),
    .A2(\reg_module/_09717_ ),
    .B1(\reg_module/_09707_ ),
    .Y(\reg_module/_00473_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17527_  (.A(\reg_module/_09711_ ),
    .B(net1348),
    .Y(\reg_module/_09718_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17528_  (.A(net966),
    .B(net979),
    .C(\reg_module/_07976_ ),
    .Y(\reg_module/_09719_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17529_  (.A(\reg_module/_09704_ ),
    .B(\reg_module/_09719_ ),
    .Y(\reg_module/_09720_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17530_  (.A1(\reg_module/_09718_ ),
    .A2(\reg_module/_09720_ ),
    .B1(\reg_module/_09707_ ),
    .Y(\reg_module/_00474_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17531_  (.A(\reg_module/_09711_ ),
    .B(net1599),
    .Y(\reg_module/_09721_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17532_  (.A(net966),
    .B(net979),
    .C(\reg_module/_07981_ ),
    .Y(\reg_module/_09722_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17533_  (.A(\reg_module/_09704_ ),
    .B(\reg_module/_09722_ ),
    .Y(\reg_module/_09723_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17534_  (.A1(\reg_module/_09721_ ),
    .A2(\reg_module/_09723_ ),
    .B1(\reg_module/_09707_ ),
    .Y(\reg_module/_00475_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17535_  (.A(\reg_module/_09711_ ),
    .B(net1791),
    .Y(\reg_module/_09724_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17536_  (.A(\reg_module/_09703_ ),
    .X(\reg_module/_09725_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17537_  (.A(net967),
    .B(net977),
    .C(\reg_module/_07989_ ),
    .Y(\reg_module/_09726_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17538_  (.A(\reg_module/_09725_ ),
    .B(\reg_module/_09726_ ),
    .Y(\reg_module/_09727_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17539_  (.A(\reg_module/_09618_ ),
    .X(\reg_module/_09728_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17540_  (.A1(\reg_module/_09724_ ),
    .A2(\reg_module/_09727_ ),
    .B1(\reg_module/_09728_ ),
    .Y(\reg_module/_00476_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17541_  (.A(\reg_module/_09711_ ),
    .B(net1789),
    .Y(\reg_module/_09729_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17542_  (.A(net967),
    .B(net976),
    .C(\reg_module/_07997_ ),
    .Y(\reg_module/_09730_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17543_  (.A(\reg_module/_09725_ ),
    .B(\reg_module/_09730_ ),
    .Y(\reg_module/_09731_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17544_  (.A1(\reg_module/_09729_ ),
    .A2(\reg_module/_09731_ ),
    .B1(\reg_module/_09728_ ),
    .Y(\reg_module/_00477_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17545_  (.A(\reg_module/_09625_ ),
    .B(net1544),
    .Y(\reg_module/_09732_ ));
 sky130_fd_sc_hd__nor3_1 \reg_module/_17546_  (.A(net967),
    .B(net976),
    .C(\reg_module/_08003_ ),
    .Y(\reg_module/_09733_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17547_  (.A(\reg_module/_09725_ ),
    .B(\reg_module/_09733_ ),
    .Y(\reg_module/_09734_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17548_  (.A1(\reg_module/_09732_ ),
    .A2(\reg_module/_09734_ ),
    .B1(\reg_module/_09728_ ),
    .Y(\reg_module/_00478_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17549_  (.A(\reg_module/_09625_ ),
    .B(net1402),
    .Y(\reg_module/_09735_ ));
 sky130_fd_sc_hd__nor3_2 \reg_module/_17550_  (.A(net967),
    .B(net976),
    .C(\reg_module/_08008_ ),
    .Y(\reg_module/_09736_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17551_  (.A(\reg_module/_09725_ ),
    .B(\reg_module/_09736_ ),
    .Y(\reg_module/_09737_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17552_  (.A1(\reg_module/_09735_ ),
    .A2(\reg_module/_09737_ ),
    .B1(\reg_module/_09728_ ),
    .Y(\reg_module/_00479_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17553_  (.A(\reg_module/_07504_ ),
    .B(\reg_module/_07506_ ),
    .C(\reg_module/_07816_ ),
    .Y(\reg_module/_09738_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17554_  (.A(\reg_module/_09738_ ),
    .Y(\reg_module/_09739_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17555_  (.A(\reg_module/_07619_ ),
    .B(\reg_module/_09739_ ),
    .C(\reg_module/_08825_ ),
    .Y(\reg_module/_09740_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_17556_  (.A(\reg_module/_09740_ ),
    .X(\reg_module/_09741_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17557_  (.A(\reg_module/_09741_ ),
    .X(\reg_module/_09742_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17558_  (.A(\reg_module/_09742_ ),
    .B(net1404),
    .Y(\reg_module/_09743_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_17559_  (.A(\reg_module/_07504_ ),
    .X(\reg_module/_09744_ ));
 sky130_fd_sc_hd__buf_1 \reg_module/_17560_  (.A(\reg_module/_09744_ ),
    .X(\reg_module/_09745_ ));
 sky130_fd_sc_hd__buf_1 \reg_module/_17561_  (.A(\reg_module/_07988_ ),
    .X(\reg_module/_09746_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17562_  (.A(\reg_module/_09745_ ),
    .B(\reg_module/_08639_ ),
    .C(\reg_module/_09746_ ),
    .D(net318),
    .X(\reg_module/_09747_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17563_  (.A(\reg_module/_09725_ ),
    .B(\reg_module/_09747_ ),
    .Y(\reg_module/_09748_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17564_  (.A1(\reg_module/_09743_ ),
    .A2(\reg_module/_09748_ ),
    .B1(\reg_module/_09728_ ),
    .Y(\reg_module/_00480_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17565_  (.A(\reg_module/_09742_ ),
    .B(net1431),
    .Y(\reg_module/_09749_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17566_  (.A(\reg_module/_09745_ ),
    .B(\reg_module/_08639_ ),
    .C(\reg_module/_09746_ ),
    .D(net317),
    .X(\reg_module/_09750_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17567_  (.A(\reg_module/_09725_ ),
    .B(\reg_module/_09750_ ),
    .Y(\reg_module/_09751_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17568_  (.A1(\reg_module/_09749_ ),
    .A2(\reg_module/_09751_ ),
    .B1(\reg_module/_09728_ ),
    .Y(\reg_module/_00481_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17569_  (.A(\reg_module/_09742_ ),
    .B(net1261),
    .Y(\reg_module/_09752_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17570_  (.A(\reg_module/_09703_ ),
    .X(\reg_module/_09753_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17571_  (.A(\reg_module/_09745_ ),
    .B(\reg_module/_08639_ ),
    .C(\reg_module/_09746_ ),
    .D(net316),
    .X(\reg_module/_09754_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17572_  (.A(\reg_module/_09753_ ),
    .B(\reg_module/_09754_ ),
    .Y(\reg_module/_09755_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_17573_  (.A(\reg_module/_09303_ ),
    .X(\reg_module/_09756_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17574_  (.A(\reg_module/_09756_ ),
    .X(\reg_module/_09757_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17575_  (.A1(\reg_module/_09752_ ),
    .A2(\reg_module/_09755_ ),
    .B1(\reg_module/_09757_ ),
    .Y(\reg_module/_00482_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17576_  (.A(\reg_module/_09742_ ),
    .B(net1640),
    .Y(\reg_module/_09758_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17577_  (.A(\reg_module/_09745_ ),
    .B(\reg_module/_08639_ ),
    .C(\reg_module/_09746_ ),
    .D(\wRegWrData[3] ),
    .X(\reg_module/_09759_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17578_  (.A(\reg_module/_09753_ ),
    .B(\reg_module/_09759_ ),
    .Y(\reg_module/_01034_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17579_  (.A1(\reg_module/_09758_ ),
    .A2(\reg_module/_01034_ ),
    .B1(\reg_module/_09757_ ),
    .Y(\reg_module/_00483_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17580_  (.A(\reg_module/_09742_ ),
    .B(net1428),
    .Y(\reg_module/_01035_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_17581_  (.A(\reg_module/_08573_ ),
    .X(\reg_module/_01036_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17582_  (.A(\reg_module/_09745_ ),
    .B(\reg_module/_01036_ ),
    .C(\reg_module/_09746_ ),
    .D(\wRegWrData[4] ),
    .X(\reg_module/_01037_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17583_  (.A(\reg_module/_09753_ ),
    .B(\reg_module/_01037_ ),
    .Y(\reg_module/_01038_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17584_  (.A1(\reg_module/_01035_ ),
    .A2(\reg_module/_01038_ ),
    .B1(\reg_module/_09757_ ),
    .Y(\reg_module/_00484_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17585_  (.A(\reg_module/_09742_ ),
    .B(net1416),
    .Y(\reg_module/_01039_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17586_  (.A(\reg_module/_09745_ ),
    .B(\reg_module/_01036_ ),
    .C(\reg_module/_09746_ ),
    .D(net314),
    .X(\reg_module/_01040_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17587_  (.A(\reg_module/_09753_ ),
    .B(\reg_module/_01040_ ),
    .Y(\reg_module/_01041_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17588_  (.A1(\reg_module/_01039_ ),
    .A2(\reg_module/_01041_ ),
    .B1(\reg_module/_09757_ ),
    .Y(\reg_module/_00485_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17589_  (.A(\reg_module/_09741_ ),
    .X(\reg_module/_01042_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17590_  (.A(\reg_module/_01042_ ),
    .B(net1597),
    .Y(\reg_module/_01043_ ));
 sky130_fd_sc_hd__buf_1 \reg_module/_17591_  (.A(\reg_module/_09744_ ),
    .X(\reg_module/_01044_ ));
 sky130_fd_sc_hd__buf_1 \reg_module/_17592_  (.A(\reg_module/_07988_ ),
    .X(\reg_module/_01045_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17593_  (.A(\reg_module/_01044_ ),
    .B(\reg_module/_01036_ ),
    .C(\reg_module/_01045_ ),
    .D(\wRegWrData[6] ),
    .X(\reg_module/_01046_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17594_  (.A(\reg_module/_09753_ ),
    .B(\reg_module/_01046_ ),
    .Y(\reg_module/_01047_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17595_  (.A1(\reg_module/_01043_ ),
    .A2(\reg_module/_01047_ ),
    .B1(\reg_module/_09757_ ),
    .Y(\reg_module/_00486_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17596_  (.A(\reg_module/_01042_ ),
    .B(net1654),
    .Y(\reg_module/_01048_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17597_  (.A(\reg_module/_01044_ ),
    .B(\reg_module/_01036_ ),
    .C(\reg_module/_01045_ ),
    .D(net313),
    .X(\reg_module/_01049_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17598_  (.A(\reg_module/_09753_ ),
    .B(\reg_module/_01049_ ),
    .Y(\reg_module/_01050_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17599_  (.A1(\reg_module/_01048_ ),
    .A2(\reg_module/_01050_ ),
    .B1(\reg_module/_09757_ ),
    .Y(\reg_module/_00487_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17600_  (.A(\reg_module/_01042_ ),
    .B(net1635),
    .Y(\reg_module/_01051_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_17601_  (.A(\reg_module/_09703_ ),
    .X(\reg_module/_01052_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17602_  (.A(\reg_module/_01044_ ),
    .B(\reg_module/_01036_ ),
    .C(\reg_module/_01045_ ),
    .D(\wRegWrData[8] ),
    .X(\reg_module/_01053_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17603_  (.A(\reg_module/_01052_ ),
    .B(\reg_module/_01053_ ),
    .Y(\reg_module/_01054_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17604_  (.A(\reg_module/_09756_ ),
    .X(\reg_module/_01055_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17605_  (.A1(\reg_module/_01051_ ),
    .A2(\reg_module/_01054_ ),
    .B1(\reg_module/_01055_ ),
    .Y(\reg_module/_00488_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17606_  (.A(\reg_module/_01042_ ),
    .B(net1522),
    .Y(\reg_module/_01056_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17607_  (.A(\reg_module/_01044_ ),
    .B(\reg_module/_01036_ ),
    .C(\reg_module/_01045_ ),
    .D(net312),
    .X(\reg_module/_01057_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17608_  (.A(\reg_module/_01052_ ),
    .B(\reg_module/_01057_ ),
    .Y(\reg_module/_01058_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17609_  (.A1(\reg_module/_01056_ ),
    .A2(\reg_module/_01058_ ),
    .B1(\reg_module/_01055_ ),
    .Y(\reg_module/_00489_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17610_  (.A(\reg_module/_01042_ ),
    .B(net1792),
    .Y(\reg_module/_01059_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_17611_  (.A(\reg_module/_08573_ ),
    .X(\reg_module/_01060_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17612_  (.A(\reg_module/_01044_ ),
    .B(\reg_module/_01060_ ),
    .C(\reg_module/_01045_ ),
    .D(net311),
    .X(\reg_module/_01061_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17613_  (.A(\reg_module/_01052_ ),
    .B(\reg_module/_01061_ ),
    .Y(\reg_module/_01062_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17614_  (.A1(\reg_module/_01059_ ),
    .A2(\reg_module/_01062_ ),
    .B1(\reg_module/_01055_ ),
    .Y(\reg_module/_00490_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17615_  (.A(\reg_module/_01042_ ),
    .B(net1663),
    .Y(\reg_module/_01063_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17616_  (.A(\reg_module/_01044_ ),
    .B(\reg_module/_01060_ ),
    .C(\reg_module/_01045_ ),
    .D(net310),
    .X(\reg_module/_01064_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17617_  (.A(\reg_module/_01052_ ),
    .B(\reg_module/_01064_ ),
    .Y(\reg_module/_01065_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17618_  (.A1(\reg_module/_01063_ ),
    .A2(\reg_module/_01065_ ),
    .B1(\reg_module/_01055_ ),
    .Y(\reg_module/_00491_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17619_  (.A(\reg_module/_09741_ ),
    .X(\reg_module/_01066_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17620_  (.A(\reg_module/_01066_ ),
    .B(net1568),
    .Y(\reg_module/_01067_ ));
 sky130_fd_sc_hd__buf_1 \reg_module/_17621_  (.A(\reg_module/_09744_ ),
    .X(\reg_module/_01068_ ));
 sky130_fd_sc_hd__buf_1 \reg_module/_17622_  (.A(\reg_module/_07842_ ),
    .X(\reg_module/_01069_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17623_  (.A(\reg_module/_01068_ ),
    .B(\reg_module/_01060_ ),
    .C(\reg_module/_01069_ ),
    .D(\wRegWrData[12] ),
    .X(\reg_module/_01070_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17624_  (.A(\reg_module/_01052_ ),
    .B(\reg_module/_01070_ ),
    .Y(\reg_module/_01071_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17625_  (.A1(\reg_module/_01067_ ),
    .A2(\reg_module/_01071_ ),
    .B1(\reg_module/_01055_ ),
    .Y(\reg_module/_00492_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17626_  (.A(\reg_module/_01066_ ),
    .B(net1326),
    .Y(\reg_module/_01072_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17627_  (.A(\reg_module/_01068_ ),
    .B(\reg_module/_01060_ ),
    .C(\reg_module/_01069_ ),
    .D(net309),
    .X(\reg_module/_01073_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17628_  (.A(\reg_module/_01052_ ),
    .B(\reg_module/_01073_ ),
    .Y(\reg_module/_01074_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17629_  (.A1(\reg_module/_01072_ ),
    .A2(\reg_module/_01074_ ),
    .B1(\reg_module/_01055_ ),
    .Y(\reg_module/_00493_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17630_  (.A(\reg_module/_01066_ ),
    .B(net1816),
    .Y(\reg_module/_01075_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17631_  (.A(\reg_module/_09703_ ),
    .X(\reg_module/_01076_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17632_  (.A(\reg_module/_01068_ ),
    .B(\reg_module/_01060_ ),
    .C(\reg_module/_01069_ ),
    .D(net308),
    .X(\reg_module/_01077_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17633_  (.A(\reg_module/_01076_ ),
    .B(\reg_module/_01077_ ),
    .Y(\reg_module/_01078_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17634_  (.A(\reg_module/_09756_ ),
    .X(\reg_module/_01079_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17635_  (.A1(\reg_module/_01075_ ),
    .A2(\reg_module/_01078_ ),
    .B1(\reg_module/_01079_ ),
    .Y(\reg_module/_00494_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17636_  (.A(\reg_module/_01066_ ),
    .B(net1786),
    .Y(\reg_module/_01080_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17637_  (.A(\reg_module/_01068_ ),
    .B(\reg_module/_01060_ ),
    .C(\reg_module/_01069_ ),
    .D(net306),
    .X(\reg_module/_01081_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17638_  (.A(\reg_module/_01076_ ),
    .B(\reg_module/_01081_ ),
    .Y(\reg_module/_01082_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17639_  (.A1(\reg_module/_01080_ ),
    .A2(\reg_module/_01082_ ),
    .B1(\reg_module/_01079_ ),
    .Y(\reg_module/_00495_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17640_  (.A(\reg_module/_01066_ ),
    .B(net1455),
    .Y(\reg_module/_01083_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17641_  (.A(\reg_module/_08573_ ),
    .X(\reg_module/_01084_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17642_  (.A(\reg_module/_01068_ ),
    .B(\reg_module/_01084_ ),
    .C(\reg_module/_01069_ ),
    .D(\wRegWrData[16] ),
    .X(\reg_module/_01085_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17643_  (.A(\reg_module/_01076_ ),
    .B(\reg_module/_01085_ ),
    .Y(\reg_module/_01086_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17644_  (.A1(\reg_module/_01083_ ),
    .A2(\reg_module/_01086_ ),
    .B1(\reg_module/_01079_ ),
    .Y(\reg_module/_00496_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17645_  (.A(\reg_module/_01066_ ),
    .B(net1693),
    .Y(\reg_module/_01087_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17646_  (.A(\reg_module/_01068_ ),
    .B(\reg_module/_01084_ ),
    .C(\reg_module/_01069_ ),
    .D(net305),
    .X(\reg_module/_01088_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17647_  (.A(\reg_module/_01076_ ),
    .B(\reg_module/_01088_ ),
    .Y(\reg_module/_01089_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17648_  (.A1(\reg_module/_01087_ ),
    .A2(\reg_module/_01089_ ),
    .B1(\reg_module/_01079_ ),
    .Y(\reg_module/_00497_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17649_  (.A(\reg_module/_09741_ ),
    .X(\reg_module/_01090_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17650_  (.A(\reg_module/_01090_ ),
    .B(net1858),
    .Y(\reg_module/_01091_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17651_  (.A(\reg_module/_09744_ ),
    .X(\reg_module/_01092_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17652_  (.A(\reg_module/_07842_ ),
    .X(\reg_module/_01093_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17653_  (.A(\reg_module/_01092_ ),
    .B(\reg_module/_01084_ ),
    .C(\reg_module/_01093_ ),
    .D(net304),
    .X(\reg_module/_01094_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17654_  (.A(\reg_module/_01076_ ),
    .B(\reg_module/_01094_ ),
    .Y(\reg_module/_01095_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17655_  (.A1(\reg_module/_01091_ ),
    .A2(\reg_module/_01095_ ),
    .B1(\reg_module/_01079_ ),
    .Y(\reg_module/_00498_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17656_  (.A(\reg_module/_01090_ ),
    .B(net1702),
    .Y(\reg_module/_01096_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17657_  (.A(\reg_module/_01092_ ),
    .B(\reg_module/_01084_ ),
    .C(\reg_module/_01093_ ),
    .D(net303),
    .X(\reg_module/_01097_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17658_  (.A(\reg_module/_01076_ ),
    .B(\reg_module/_01097_ ),
    .Y(\reg_module/_01098_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17659_  (.A1(\reg_module/_01096_ ),
    .A2(\reg_module/_01098_ ),
    .B1(\reg_module/_01079_ ),
    .Y(\reg_module/_00499_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17660_  (.A(\reg_module/_01090_ ),
    .B(net1493),
    .Y(\reg_module/_01099_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17661_  (.A(\reg_module/_09703_ ),
    .X(\reg_module/_01100_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17662_  (.A(\reg_module/_01092_ ),
    .B(\reg_module/_01084_ ),
    .C(\reg_module/_01093_ ),
    .D(net302),
    .X(\reg_module/_01101_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17663_  (.A(\reg_module/_01100_ ),
    .B(\reg_module/_01101_ ),
    .Y(\reg_module/_01102_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17664_  (.A(\reg_module/_09756_ ),
    .X(\reg_module/_01103_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17665_  (.A1(\reg_module/_01099_ ),
    .A2(\reg_module/_01102_ ),
    .B1(\reg_module/_01103_ ),
    .Y(\reg_module/_00500_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17666_  (.A(\reg_module/_01090_ ),
    .B(net1520),
    .Y(\reg_module/_01104_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17667_  (.A(\reg_module/_01092_ ),
    .B(\reg_module/_01084_ ),
    .C(\reg_module/_01093_ ),
    .D(net301),
    .X(\reg_module/_01105_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17668_  (.A(\reg_module/_01100_ ),
    .B(\reg_module/_01105_ ),
    .Y(\reg_module/_01106_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17669_  (.A1(\reg_module/_01104_ ),
    .A2(\reg_module/_01106_ ),
    .B1(\reg_module/_01103_ ),
    .Y(\reg_module/_00501_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17670_  (.A(\reg_module/_01090_ ),
    .B(net1325),
    .Y(\reg_module/_01107_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17671_  (.A(\reg_module/_07626_ ),
    .X(\reg_module/_01108_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17672_  (.A(\reg_module/_01092_ ),
    .B(\reg_module/_01108_ ),
    .C(\reg_module/_01093_ ),
    .D(net300),
    .X(\reg_module/_01109_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17673_  (.A(\reg_module/_01100_ ),
    .B(\reg_module/_01109_ ),
    .Y(\reg_module/_01110_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17674_  (.A1(\reg_module/_01107_ ),
    .A2(\reg_module/_01110_ ),
    .B1(\reg_module/_01103_ ),
    .Y(\reg_module/_00502_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17675_  (.A(\reg_module/_01090_ ),
    .B(net1241),
    .Y(\reg_module/_01111_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17676_  (.A(\reg_module/_01092_ ),
    .B(\reg_module/_01108_ ),
    .C(\reg_module/_01093_ ),
    .D(net299),
    .X(\reg_module/_01112_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17677_  (.A(\reg_module/_01100_ ),
    .B(\reg_module/_01112_ ),
    .Y(\reg_module/_01113_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17678_  (.A1(\reg_module/_01111_ ),
    .A2(\reg_module/_01113_ ),
    .B1(\reg_module/_01103_ ),
    .Y(\reg_module/_00503_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17679_  (.A(\reg_module/_09740_ ),
    .X(\reg_module/_01114_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17680_  (.A(\reg_module/_01114_ ),
    .B(net1243),
    .Y(\reg_module/_01115_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17681_  (.A(\reg_module/_07504_ ),
    .X(\reg_module/_01116_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17682_  (.A(\reg_module/_07842_ ),
    .X(\reg_module/_01117_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17683_  (.A(\reg_module/_01116_ ),
    .B(\reg_module/_01108_ ),
    .C(\reg_module/_01117_ ),
    .D(net298),
    .X(\reg_module/_01118_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17684_  (.A(\reg_module/_01100_ ),
    .B(\reg_module/_01118_ ),
    .Y(\reg_module/_01119_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17685_  (.A1(\reg_module/_01115_ ),
    .A2(\reg_module/_01119_ ),
    .B1(\reg_module/_01103_ ),
    .Y(\reg_module/_00504_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17686_  (.A(\reg_module/_01114_ ),
    .B(net1272),
    .Y(\reg_module/_01120_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17687_  (.A(\reg_module/_01116_ ),
    .B(\reg_module/_01108_ ),
    .C(\reg_module/_01117_ ),
    .D(net296),
    .X(\reg_module/_01121_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17688_  (.A(\reg_module/_01100_ ),
    .B(\reg_module/_01121_ ),
    .Y(\reg_module/_01122_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17689_  (.A1(\reg_module/_01120_ ),
    .A2(\reg_module/_01122_ ),
    .B1(\reg_module/_01103_ ),
    .Y(\reg_module/_00505_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17690_  (.A(\reg_module/_01114_ ),
    .B(net1437),
    .Y(\reg_module/_01123_ ));
 sky130_fd_sc_hd__buf_8 \reg_module/_17691_  (.A(\reg_module/_08183_ ),
    .X(\reg_module/_01124_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17692_  (.A(\reg_module/_01124_ ),
    .X(\reg_module/_01125_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17693_  (.A(\reg_module/_01116_ ),
    .B(\reg_module/_01108_ ),
    .C(\reg_module/_01117_ ),
    .D(net294),
    .X(\reg_module/_01126_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17694_  (.A(\reg_module/_01125_ ),
    .B(\reg_module/_01126_ ),
    .Y(\reg_module/_01127_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17695_  (.A(\reg_module/_09756_ ),
    .X(\reg_module/_01128_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17696_  (.A1(\reg_module/_01123_ ),
    .A2(\reg_module/_01127_ ),
    .B1(\reg_module/_01128_ ),
    .Y(\reg_module/_00506_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17697_  (.A(\reg_module/_01114_ ),
    .B(net1322),
    .Y(\reg_module/_01129_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17698_  (.A(\reg_module/_01116_ ),
    .B(\reg_module/_01108_ ),
    .C(\reg_module/_01117_ ),
    .D(net293),
    .X(\reg_module/_01130_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17699_  (.A(\reg_module/_01125_ ),
    .B(\reg_module/_01130_ ),
    .Y(\reg_module/_01131_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17700_  (.A1(\reg_module/_01129_ ),
    .A2(\reg_module/_01131_ ),
    .B1(\reg_module/_01128_ ),
    .Y(\reg_module/_00507_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17701_  (.A(\reg_module/_01114_ ),
    .B(net1407),
    .Y(\reg_module/_01132_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17702_  (.A(\reg_module/_01116_ ),
    .B(\reg_module/_08526_ ),
    .C(\reg_module/_01117_ ),
    .D(net292),
    .X(\reg_module/_01133_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17703_  (.A(\reg_module/_01125_ ),
    .B(\reg_module/_01133_ ),
    .Y(\reg_module/_01134_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17704_  (.A1(\reg_module/_01132_ ),
    .A2(\reg_module/_01134_ ),
    .B1(\reg_module/_01128_ ),
    .Y(\reg_module/_00508_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17705_  (.A(\reg_module/_01114_ ),
    .B(net1513),
    .Y(\reg_module/_01135_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17706_  (.A(\reg_module/_01116_ ),
    .B(\reg_module/_08526_ ),
    .C(\reg_module/_01117_ ),
    .D(net290),
    .X(\reg_module/_01136_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17707_  (.A(\reg_module/_01125_ ),
    .B(\reg_module/_01136_ ),
    .Y(\reg_module/_01137_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17708_  (.A1(\reg_module/_01135_ ),
    .A2(\reg_module/_01137_ ),
    .B1(\reg_module/_01128_ ),
    .Y(\reg_module/_00509_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17709_  (.A(\reg_module/_09741_ ),
    .B(net1273),
    .Y(\reg_module/_01138_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17710_  (.A(\reg_module/_09744_ ),
    .B(\reg_module/_08526_ ),
    .C(\reg_module/_07818_ ),
    .D(net289),
    .X(\reg_module/_01139_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17711_  (.A(\reg_module/_01125_ ),
    .B(\reg_module/_01139_ ),
    .Y(\reg_module/_01140_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17712_  (.A1(\reg_module/_01138_ ),
    .A2(\reg_module/_01140_ ),
    .B1(\reg_module/_01128_ ),
    .Y(\reg_module/_00510_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17713_  (.A(\reg_module/_09741_ ),
    .B(net1274),
    .Y(\reg_module/_01141_ ));
 sky130_fd_sc_hd__and4_1 \reg_module/_17714_  (.A(\reg_module/_09744_ ),
    .B(\reg_module/_08526_ ),
    .C(\reg_module/_07818_ ),
    .D(net287),
    .X(\reg_module/_01142_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17715_  (.A(\reg_module/_01125_ ),
    .B(\reg_module/_01142_ ),
    .Y(\reg_module/_01143_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17716_  (.A1(\reg_module/_01141_ ),
    .A2(\reg_module/_01143_ ),
    .B1(\reg_module/_01128_ ),
    .Y(\reg_module/_00511_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17717_  (.A(\reg_module/_01124_ ),
    .X(\reg_module/_01144_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_17718_  (.A(\reg_module/_08503_ ),
    .X(\reg_module/_01145_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17719_  (.A(\reg_module/_07500_ ),
    .B(\reg_module/_07501_ ),
    .Y(\reg_module/_01146_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17720_  (.A(\reg_module/_01146_ ),
    .X(\reg_module/_01147_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17721_  (.A(\reg_module/_01147_ ),
    .X(\reg_module/_01148_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17722_  (.A(\reg_module/_07513_ ),
    .B(\reg_module/_01148_ ),
    .Y(\reg_module/_01149_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17723_  (.A(\reg_module/_01144_ ),
    .B(\reg_module/_01145_ ),
    .C(\reg_module/_01149_ ),
    .Y(\reg_module/_01150_ ));
 sky130_fd_sc_hd__buf_8 \reg_module/_17724_  (.A(\reg_module/_07621_ ),
    .X(\reg_module/_01151_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17725_  (.A(\reg_module/_01151_ ),
    .X(\reg_module/_01152_ ));
 sky130_fd_sc_hd__nand3_2 \reg_module/_17726_  (.A(\reg_module/_09738_ ),
    .B(\reg_module/_07622_ ),
    .C(rRegWrEn2),
    .Y(\reg_module/_01153_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_17727_  (.A(\reg_module/_01153_ ),
    .X(\reg_module/_01154_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_17728_  (.A(\reg_module/_01154_ ),
    .X(\reg_module/_01155_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17729_  (.A(\reg_module/_01155_ ),
    .X(\reg_module/_01156_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17730_  (.A(\reg_module/_01156_ ),
    .X(\reg_module/_01157_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17731_  (.A1(\reg_module/_01152_ ),
    .A2(\reg_module/_01157_ ),
    .B1(\reg_module/gprf[512] ),
    .Y(\reg_module/_01158_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17732_  (.A(\reg_module/_09756_ ),
    .X(\reg_module/_01159_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17733_  (.A1(\reg_module/_01150_ ),
    .A2(\reg_module/_01158_ ),
    .B1(\reg_module/_01159_ ),
    .Y(\reg_module/_00512_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17734_  (.A(\reg_module/_07516_ ),
    .B(\reg_module/_01148_ ),
    .Y(\reg_module/_01160_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17735_  (.A(\reg_module/_01144_ ),
    .B(\reg_module/_01145_ ),
    .C(\reg_module/_01160_ ),
    .Y(\reg_module/_01161_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17736_  (.A1(\reg_module/_01152_ ),
    .A2(\reg_module/_01157_ ),
    .B1(\reg_module/gprf[513] ),
    .Y(\reg_module/_01162_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17737_  (.A1(\reg_module/_01161_ ),
    .A2(\reg_module/_01162_ ),
    .B1(\reg_module/_01159_ ),
    .Y(\reg_module/_00513_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17738_  (.A(\reg_module/_07519_ ),
    .B(\reg_module/_01148_ ),
    .Y(\reg_module/_01163_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17739_  (.A(\reg_module/_01144_ ),
    .B(\reg_module/_01145_ ),
    .C(\reg_module/_01163_ ),
    .Y(\reg_module/_01164_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17740_  (.A1(\reg_module/_01152_ ),
    .A2(\reg_module/_01157_ ),
    .B1(net2127),
    .Y(\reg_module/_01165_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17741_  (.A1(\reg_module/_01164_ ),
    .A2(\reg_module/_01165_ ),
    .B1(\reg_module/_01159_ ),
    .Y(\reg_module/_00514_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17742_  (.A(\reg_module/_07522_ ),
    .B(\reg_module/_01148_ ),
    .Y(\reg_module/_01166_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17743_  (.A(\reg_module/_01144_ ),
    .B(\reg_module/_01145_ ),
    .C(\reg_module/_01166_ ),
    .Y(\reg_module/_01167_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17744_  (.A1(\reg_module/_01152_ ),
    .A2(\reg_module/_01157_ ),
    .B1(net1990),
    .Y(\reg_module/_01168_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17745_  (.A1(\reg_module/_01167_ ),
    .A2(\reg_module/_01168_ ),
    .B1(\reg_module/_01159_ ),
    .Y(\reg_module/_00515_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17746_  (.A(\reg_module/_07527_ ),
    .B(\reg_module/_01148_ ),
    .Y(\reg_module/_01169_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17747_  (.A(\reg_module/_01144_ ),
    .B(\reg_module/_01145_ ),
    .C(\reg_module/_01169_ ),
    .Y(\reg_module/_01170_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17748_  (.A1(\reg_module/_01152_ ),
    .A2(\reg_module/_01157_ ),
    .B1(net2003),
    .Y(\reg_module/_01171_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17749_  (.A1(\reg_module/_01170_ ),
    .A2(\reg_module/_01171_ ),
    .B1(\reg_module/_01159_ ),
    .Y(\reg_module/_00516_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17750_  (.A(\reg_module/_07530_ ),
    .B(\reg_module/_01148_ ),
    .Y(\reg_module/_01172_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17751_  (.A(\reg_module/_01144_ ),
    .B(\reg_module/_01145_ ),
    .C(\reg_module/_01172_ ),
    .Y(\reg_module/_01173_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17752_  (.A1(\reg_module/_01152_ ),
    .A2(\reg_module/_01157_ ),
    .B1(net1996),
    .Y(\reg_module/_01174_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17753_  (.A1(\reg_module/_01173_ ),
    .A2(\reg_module/_01174_ ),
    .B1(\reg_module/_01159_ ),
    .Y(\reg_module/_00517_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17754_  (.A(\reg_module/_01124_ ),
    .X(\reg_module/_01175_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_17755_  (.A(\reg_module/_08503_ ),
    .X(\reg_module/_01176_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_17756_  (.A(\reg_module/_01147_ ),
    .X(\reg_module/_01177_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17757_  (.A(\reg_module/_07534_ ),
    .B(\reg_module/_01177_ ),
    .Y(\reg_module/_01178_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17758_  (.A(\reg_module/_01175_ ),
    .B(\reg_module/_01176_ ),
    .C(\reg_module/_01178_ ),
    .Y(\reg_module/_01179_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17759_  (.A(\reg_module/_01151_ ),
    .X(\reg_module/_01180_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17760_  (.A(\reg_module/_01156_ ),
    .X(\reg_module/_01181_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17761_  (.A1(\reg_module/_01180_ ),
    .A2(\reg_module/_01181_ ),
    .B1(net1907),
    .Y(\reg_module/_01182_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17762_  (.A(\reg_module/_09303_ ),
    .X(\reg_module/_01183_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17763_  (.A(\reg_module/_01183_ ),
    .X(\reg_module/_01184_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17764_  (.A1(\reg_module/_01179_ ),
    .A2(\reg_module/_01182_ ),
    .B1(\reg_module/_01184_ ),
    .Y(\reg_module/_00518_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17765_  (.A(\reg_module/_07537_ ),
    .B(\reg_module/_01177_ ),
    .Y(\reg_module/_01185_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17766_  (.A(\reg_module/_01175_ ),
    .B(\reg_module/_01176_ ),
    .C(\reg_module/_01185_ ),
    .Y(\reg_module/_01186_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17767_  (.A1(\reg_module/_01180_ ),
    .A2(\reg_module/_01181_ ),
    .B1(net1963),
    .Y(\reg_module/_01187_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17768_  (.A1(\reg_module/_01186_ ),
    .A2(\reg_module/_01187_ ),
    .B1(\reg_module/_01184_ ),
    .Y(\reg_module/_00519_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17769_  (.A(\reg_module/_07540_ ),
    .B(\reg_module/_01177_ ),
    .Y(\reg_module/_01188_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17770_  (.A(\reg_module/_01175_ ),
    .B(\reg_module/_01176_ ),
    .C(\reg_module/_01188_ ),
    .Y(\reg_module/_01189_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17771_  (.A1(\reg_module/_01180_ ),
    .A2(\reg_module/_01181_ ),
    .B1(net2078),
    .Y(\reg_module/_01190_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17772_  (.A1(\reg_module/_01189_ ),
    .A2(\reg_module/_01190_ ),
    .B1(\reg_module/_01184_ ),
    .Y(\reg_module/_00520_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17773_  (.A(\reg_module/_07543_ ),
    .B(\reg_module/_01177_ ),
    .Y(\reg_module/_01191_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17774_  (.A(\reg_module/_01175_ ),
    .B(\reg_module/_01176_ ),
    .C(\reg_module/_01191_ ),
    .Y(\reg_module/_01192_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17775_  (.A1(\reg_module/_01180_ ),
    .A2(\reg_module/_01181_ ),
    .B1(net1812),
    .Y(\reg_module/_01193_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17776_  (.A1(\reg_module/_01192_ ),
    .A2(\reg_module/_01193_ ),
    .B1(\reg_module/_01184_ ),
    .Y(\reg_module/_00521_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17777_  (.A(\reg_module/_07547_ ),
    .B(\reg_module/_01177_ ),
    .Y(\reg_module/_01194_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17778_  (.A(\reg_module/_01175_ ),
    .B(\reg_module/_01176_ ),
    .C(\reg_module/_01194_ ),
    .Y(\reg_module/_01195_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17779_  (.A1(\reg_module/_01180_ ),
    .A2(\reg_module/_01181_ ),
    .B1(net1952),
    .Y(\reg_module/_01196_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17780_  (.A1(\reg_module/_01195_ ),
    .A2(\reg_module/_01196_ ),
    .B1(\reg_module/_01184_ ),
    .Y(\reg_module/_00522_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17781_  (.A(\reg_module/_07550_ ),
    .B(\reg_module/_01177_ ),
    .Y(\reg_module/_01197_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17782_  (.A(\reg_module/_01175_ ),
    .B(\reg_module/_01176_ ),
    .C(\reg_module/_01197_ ),
    .Y(\reg_module/_01198_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17783_  (.A1(\reg_module/_01180_ ),
    .A2(\reg_module/_01181_ ),
    .B1(net2133),
    .Y(\reg_module/_01199_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17784_  (.A1(\reg_module/_01198_ ),
    .A2(\reg_module/_01199_ ),
    .B1(\reg_module/_01184_ ),
    .Y(\reg_module/_00523_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17785_  (.A(\reg_module/_01124_ ),
    .X(\reg_module/_01200_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_17786_  (.A(\reg_module/_08028_ ),
    .X(\reg_module/_01201_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_17787_  (.A(\reg_module/_01147_ ),
    .X(\reg_module/_01202_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17788_  (.A(\reg_module/_07554_ ),
    .B(\reg_module/_01202_ ),
    .Y(\reg_module/_01203_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17789_  (.A(\reg_module/_01200_ ),
    .B(\reg_module/_01201_ ),
    .C(\reg_module/_01203_ ),
    .Y(\reg_module/_01204_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17790_  (.A(\reg_module/_01151_ ),
    .X(\reg_module/_01205_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17791_  (.A(\reg_module/_01156_ ),
    .X(\reg_module/_01206_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17792_  (.A1(\reg_module/_01205_ ),
    .A2(\reg_module/_01206_ ),
    .B1(net2006),
    .Y(\reg_module/_01207_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17793_  (.A(\reg_module/_01183_ ),
    .X(\reg_module/_01208_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17794_  (.A1(\reg_module/_01204_ ),
    .A2(\reg_module/_01207_ ),
    .B1(\reg_module/_01208_ ),
    .Y(\reg_module/_00524_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17795_  (.A(\reg_module/_07557_ ),
    .B(\reg_module/_01202_ ),
    .Y(\reg_module/_01209_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17796_  (.A(\reg_module/_01200_ ),
    .B(\reg_module/_01201_ ),
    .C(\reg_module/_01209_ ),
    .Y(\reg_module/_01210_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17797_  (.A1(\reg_module/_01205_ ),
    .A2(\reg_module/_01206_ ),
    .B1(net2061),
    .Y(\reg_module/_01211_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17798_  (.A1(\reg_module/_01210_ ),
    .A2(\reg_module/_01211_ ),
    .B1(\reg_module/_01208_ ),
    .Y(\reg_module/_00525_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17799_  (.A(\reg_module/_07560_ ),
    .B(\reg_module/_01202_ ),
    .Y(\reg_module/_01212_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17800_  (.A(\reg_module/_01200_ ),
    .B(\reg_module/_01201_ ),
    .C(\reg_module/_01212_ ),
    .Y(\reg_module/_01213_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17801_  (.A1(\reg_module/_01205_ ),
    .A2(\reg_module/_01206_ ),
    .B1(net2110),
    .Y(\reg_module/_01214_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17802_  (.A1(\reg_module/_01213_ ),
    .A2(\reg_module/_01214_ ),
    .B1(\reg_module/_01208_ ),
    .Y(\reg_module/_00526_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17803_  (.A(\reg_module/_07563_ ),
    .B(\reg_module/_01202_ ),
    .Y(\reg_module/_01215_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17804_  (.A(\reg_module/_01200_ ),
    .B(\reg_module/_01201_ ),
    .C(\reg_module/_01215_ ),
    .Y(\reg_module/_01216_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17805_  (.A1(\reg_module/_01205_ ),
    .A2(\reg_module/_01206_ ),
    .B1(net1969),
    .Y(\reg_module/_01217_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17806_  (.A1(\reg_module/_01216_ ),
    .A2(\reg_module/_01217_ ),
    .B1(\reg_module/_01208_ ),
    .Y(\reg_module/_00527_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17807_  (.A(\reg_module/_07567_ ),
    .B(\reg_module/_01202_ ),
    .Y(\reg_module/_01218_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17808_  (.A(\reg_module/_01200_ ),
    .B(\reg_module/_01201_ ),
    .C(\reg_module/_01218_ ),
    .Y(\reg_module/_01219_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17809_  (.A1(\reg_module/_01205_ ),
    .A2(\reg_module/_01206_ ),
    .B1(net1868),
    .Y(\reg_module/_01220_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17810_  (.A1(\reg_module/_01219_ ),
    .A2(\reg_module/_01220_ ),
    .B1(\reg_module/_01208_ ),
    .Y(\reg_module/_00528_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17811_  (.A(\reg_module/_07570_ ),
    .B(\reg_module/_01202_ ),
    .Y(\reg_module/_01221_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17812_  (.A(\reg_module/_01200_ ),
    .B(\reg_module/_01201_ ),
    .C(\reg_module/_01221_ ),
    .Y(\reg_module/_01222_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17813_  (.A1(\reg_module/_01205_ ),
    .A2(\reg_module/_01206_ ),
    .B1(net2119),
    .Y(\reg_module/_01223_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17814_  (.A1(\reg_module/_01222_ ),
    .A2(\reg_module/_01223_ ),
    .B1(\reg_module/_01208_ ),
    .Y(\reg_module/_00529_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17815_  (.A(\reg_module/_01124_ ),
    .X(\reg_module/_01224_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_17816_  (.A(\reg_module/_08028_ ),
    .X(\reg_module/_01225_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_17817_  (.A(\reg_module/_01147_ ),
    .X(\reg_module/_01226_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17818_  (.A(\reg_module/_07574_ ),
    .B(\reg_module/_01226_ ),
    .Y(\reg_module/_01227_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17819_  (.A(\reg_module/_01224_ ),
    .B(\reg_module/_01225_ ),
    .C(\reg_module/_01227_ ),
    .Y(\reg_module/_01228_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17820_  (.A(\reg_module/_01151_ ),
    .X(\reg_module/_01229_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17821_  (.A(\reg_module/_01156_ ),
    .X(\reg_module/_01230_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17822_  (.A1(\reg_module/_01229_ ),
    .A2(\reg_module/_01230_ ),
    .B1(net2194),
    .Y(\reg_module/_01231_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17823_  (.A(\reg_module/_01183_ ),
    .X(\reg_module/_01232_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17824_  (.A1(\reg_module/_01228_ ),
    .A2(\reg_module/_01231_ ),
    .B1(\reg_module/_01232_ ),
    .Y(\reg_module/_00530_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17825_  (.A(\reg_module/_07577_ ),
    .B(\reg_module/_01226_ ),
    .Y(\reg_module/_01233_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17826_  (.A(\reg_module/_01224_ ),
    .B(\reg_module/_01225_ ),
    .C(\reg_module/_01233_ ),
    .Y(\reg_module/_01234_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17827_  (.A1(\reg_module/_01229_ ),
    .A2(\reg_module/_01230_ ),
    .B1(net2124),
    .Y(\reg_module/_01235_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17828_  (.A1(\reg_module/_01234_ ),
    .A2(\reg_module/_01235_ ),
    .B1(\reg_module/_01232_ ),
    .Y(\reg_module/_00531_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17829_  (.A(\reg_module/_07580_ ),
    .B(\reg_module/_01226_ ),
    .Y(\reg_module/_01236_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17830_  (.A(\reg_module/_01224_ ),
    .B(\reg_module/_01225_ ),
    .C(\reg_module/_01236_ ),
    .Y(\reg_module/_01237_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17831_  (.A1(\reg_module/_01229_ ),
    .A2(\reg_module/_01230_ ),
    .B1(net2143),
    .Y(\reg_module/_01238_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17832_  (.A1(\reg_module/_01237_ ),
    .A2(\reg_module/_01238_ ),
    .B1(\reg_module/_01232_ ),
    .Y(\reg_module/_00532_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17833_  (.A(\reg_module/_07583_ ),
    .B(\reg_module/_01226_ ),
    .Y(\reg_module/_01239_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17834_  (.A(\reg_module/_01224_ ),
    .B(\reg_module/_01225_ ),
    .C(\reg_module/_01239_ ),
    .Y(\reg_module/_01240_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17835_  (.A1(\reg_module/_01229_ ),
    .A2(\reg_module/_01230_ ),
    .B1(net1750),
    .Y(\reg_module/_01241_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17836_  (.A1(\reg_module/_01240_ ),
    .A2(\reg_module/_01241_ ),
    .B1(\reg_module/_01232_ ),
    .Y(\reg_module/_00533_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17837_  (.A(\reg_module/_07587_ ),
    .B(\reg_module/_01226_ ),
    .Y(\reg_module/_01242_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17838_  (.A(\reg_module/_01224_ ),
    .B(\reg_module/_01225_ ),
    .C(\reg_module/_01242_ ),
    .Y(\reg_module/_01243_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17839_  (.A1(\reg_module/_01229_ ),
    .A2(\reg_module/_01230_ ),
    .B1(net1793),
    .Y(\reg_module/_01244_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17840_  (.A1(\reg_module/_01243_ ),
    .A2(\reg_module/_01244_ ),
    .B1(\reg_module/_01232_ ),
    .Y(\reg_module/_00534_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17841_  (.A(\reg_module/_07590_ ),
    .B(\reg_module/_01226_ ),
    .Y(\reg_module/_01245_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17842_  (.A(\reg_module/_01224_ ),
    .B(\reg_module/_01225_ ),
    .C(\reg_module/_01245_ ),
    .Y(\reg_module/_01246_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17843_  (.A1(\reg_module/_01229_ ),
    .A2(\reg_module/_01230_ ),
    .B1(net1986),
    .Y(\reg_module/_01247_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17844_  (.A1(\reg_module/_01246_ ),
    .A2(\reg_module/_01247_ ),
    .B1(\reg_module/_01232_ ),
    .Y(\reg_module/_00535_ ));
 sky130_fd_sc_hd__buf_6 \reg_module/_17845_  (.A(\reg_module/_01124_ ),
    .X(\reg_module/_01248_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_17846_  (.A(\reg_module/_08028_ ),
    .X(\reg_module/_01249_ ));
 sky130_fd_sc_hd__dlymetal6s2s_1 \reg_module/_17847_  (.A(\reg_module/_01146_ ),
    .X(\reg_module/_01250_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17848_  (.A(\reg_module/_07594_ ),
    .B(\reg_module/_01250_ ),
    .Y(\reg_module/_01251_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17849_  (.A(\reg_module/_01248_ ),
    .B(\reg_module/_01249_ ),
    .C(\reg_module/_01251_ ),
    .Y(\reg_module/_01252_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17850_  (.A(\reg_module/_07621_ ),
    .X(\reg_module/_01253_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_17851_  (.A(\reg_module/_01154_ ),
    .X(\reg_module/_01254_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17852_  (.A(\reg_module/_01254_ ),
    .X(\reg_module/_01255_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17853_  (.A1(\reg_module/_01253_ ),
    .A2(\reg_module/_01255_ ),
    .B1(net2001),
    .Y(\reg_module/_01256_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17854_  (.A(\reg_module/_01183_ ),
    .X(\reg_module/_01257_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17855_  (.A1(\reg_module/_01252_ ),
    .A2(\reg_module/_01256_ ),
    .B1(\reg_module/_01257_ ),
    .Y(\reg_module/_00536_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17856_  (.A(\reg_module/_07597_ ),
    .B(\reg_module/_01250_ ),
    .Y(\reg_module/_01258_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17857_  (.A(\reg_module/_01248_ ),
    .B(\reg_module/_01249_ ),
    .C(\reg_module/_01258_ ),
    .Y(\reg_module/_01259_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17858_  (.A1(\reg_module/_01253_ ),
    .A2(\reg_module/_01255_ ),
    .B1(net2039),
    .Y(\reg_module/_01260_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17859_  (.A1(\reg_module/_01259_ ),
    .A2(\reg_module/_01260_ ),
    .B1(\reg_module/_01257_ ),
    .Y(\reg_module/_00537_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17860_  (.A(\reg_module/_07600_ ),
    .B(\reg_module/_01250_ ),
    .Y(\reg_module/_01261_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17861_  (.A(\reg_module/_01248_ ),
    .B(\reg_module/_01249_ ),
    .C(\reg_module/_01261_ ),
    .Y(\reg_module/_01262_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17862_  (.A1(\reg_module/_01253_ ),
    .A2(\reg_module/_01255_ ),
    .B1(net1894),
    .Y(\reg_module/_01263_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17863_  (.A1(\reg_module/_01262_ ),
    .A2(\reg_module/_01263_ ),
    .B1(\reg_module/_01257_ ),
    .Y(\reg_module/_00538_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17864_  (.A(\reg_module/_07603_ ),
    .B(\reg_module/_01250_ ),
    .Y(\reg_module/_01264_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17865_  (.A(\reg_module/_01248_ ),
    .B(\reg_module/_01249_ ),
    .C(\reg_module/_01264_ ),
    .Y(\reg_module/_01265_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17866_  (.A1(\reg_module/_01253_ ),
    .A2(\reg_module/_01255_ ),
    .B1(net1857),
    .Y(\reg_module/_01266_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17867_  (.A1(\reg_module/_01265_ ),
    .A2(\reg_module/_01266_ ),
    .B1(\reg_module/_01257_ ),
    .Y(\reg_module/_00539_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17868_  (.A(\reg_module/_07606_ ),
    .B(\reg_module/_01250_ ),
    .Y(\reg_module/_01267_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17869_  (.A(\reg_module/_01248_ ),
    .B(\reg_module/_01249_ ),
    .C(\reg_module/_01267_ ),
    .Y(\reg_module/_01268_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17870_  (.A1(\reg_module/_01253_ ),
    .A2(\reg_module/_01255_ ),
    .B1(net1982),
    .Y(\reg_module/_01269_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17871_  (.A1(\reg_module/_01268_ ),
    .A2(\reg_module/_01269_ ),
    .B1(\reg_module/_01257_ ),
    .Y(\reg_module/_00540_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17872_  (.A(\reg_module/_07609_ ),
    .B(\reg_module/_01250_ ),
    .Y(\reg_module/_01270_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17873_  (.A(\reg_module/_01248_ ),
    .B(\reg_module/_01249_ ),
    .C(\reg_module/_01270_ ),
    .Y(\reg_module/_01271_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17874_  (.A1(\reg_module/_01253_ ),
    .A2(\reg_module/_01255_ ),
    .B1(net2004),
    .Y(\reg_module/_01272_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17875_  (.A1(\reg_module/_01271_ ),
    .A2(\reg_module/_01272_ ),
    .B1(\reg_module/_01257_ ),
    .Y(\reg_module/_00541_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17876_  (.A(\reg_module/_07612_ ),
    .B(\reg_module/_01147_ ),
    .Y(\reg_module/_01273_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17877_  (.A(\reg_module/_08185_ ),
    .B(\reg_module/_08023_ ),
    .C(\reg_module/_01273_ ),
    .Y(\reg_module/_01274_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17878_  (.A(\reg_module/_01254_ ),
    .X(\reg_module/_01275_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17879_  (.A1(\reg_module/_01151_ ),
    .A2(\reg_module/_01275_ ),
    .B1(net1743),
    .Y(\reg_module/_01276_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17880_  (.A(\reg_module/_01183_ ),
    .X(\reg_module/_01277_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17881_  (.A1(\reg_module/_01274_ ),
    .A2(\reg_module/_01276_ ),
    .B1(\reg_module/_01277_ ),
    .Y(\reg_module/_00542_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_17882_  (.A(\reg_module/_07615_ ),
    .B(\reg_module/_01147_ ),
    .Y(\reg_module/_01278_ ));
 sky130_fd_sc_hd__nand3_1 \reg_module/_17883_  (.A(\reg_module/_08185_ ),
    .B(\reg_module/_08023_ ),
    .C(\reg_module/_01278_ ),
    .Y(\reg_module/_01279_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_17884_  (.A1(\reg_module/_01151_ ),
    .A2(\reg_module/_01275_ ),
    .B1(net1770),
    .Y(\reg_module/_01280_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17885_  (.A1(\reg_module/_01279_ ),
    .A2(\reg_module/_01280_ ),
    .B1(\reg_module/_01277_ ),
    .Y(\reg_module/_00543_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_17886_  (.A(\reg_module/_07635_ ),
    .B(\reg_module/_01153_ ),
    .Y(\reg_module/_01281_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17887_  (.A(\reg_module/_01281_ ),
    .B(\reg_module/_07630_ ),
    .Y(\reg_module/_01282_ ));
 sky130_fd_sc_hd__buf_8 \reg_module/_17888_  (.A(\reg_module/_01282_ ),
    .X(\reg_module/_01283_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17889_  (.A(\reg_module/_01283_ ),
    .X(\reg_module/_01284_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17890_  (.A(\reg_module/_01284_ ),
    .B(net1684),
    .Y(\reg_module/_01285_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_17891_  (.A(\reg_module/_01153_ ),
    .Y(\reg_module/_01286_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_17892_  (.A(\reg_module/_01286_ ),
    .X(\reg_module/_01287_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17893_  (.A(\reg_module/_01287_ ),
    .X(\reg_module/_01288_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17894_  (.A(\reg_module/_07651_ ),
    .B(\reg_module/_01288_ ),
    .Y(\reg_module/_01289_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17895_  (.A1(\reg_module/_01285_ ),
    .A2(\reg_module/_01289_ ),
    .B1(\reg_module/_01277_ ),
    .Y(\reg_module/_00544_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17896_  (.A(\reg_module/_01284_ ),
    .B(net1320),
    .Y(\reg_module/_01290_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17897_  (.A(\reg_module/_07659_ ),
    .B(\reg_module/_01288_ ),
    .Y(\reg_module/_01291_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17898_  (.A1(\reg_module/_01290_ ),
    .A2(\reg_module/_01291_ ),
    .B1(\reg_module/_01277_ ),
    .Y(\reg_module/_00545_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17899_  (.A(\reg_module/_01284_ ),
    .B(net1642),
    .Y(\reg_module/_01292_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17900_  (.A(\reg_module/_07665_ ),
    .B(\reg_module/_01288_ ),
    .Y(\reg_module/_01293_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17901_  (.A1(\reg_module/_01292_ ),
    .A2(\reg_module/_01293_ ),
    .B1(\reg_module/_01277_ ),
    .Y(\reg_module/_00546_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17902_  (.A(\reg_module/_01284_ ),
    .B(net2041),
    .Y(\reg_module/_01294_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17903_  (.A(\reg_module/_07669_ ),
    .B(\reg_module/_01288_ ),
    .Y(\reg_module/_01295_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17904_  (.A1(\reg_module/_01294_ ),
    .A2(\reg_module/_01295_ ),
    .B1(\reg_module/_01277_ ),
    .Y(\reg_module/_00547_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17905_  (.A(\reg_module/_01284_ ),
    .B(net1570),
    .Y(\reg_module/_01296_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17906_  (.A(\reg_module/_07673_ ),
    .B(\reg_module/_01288_ ),
    .Y(\reg_module/_01297_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17907_  (.A(\reg_module/_01183_ ),
    .X(\reg_module/_01298_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17908_  (.A1(\reg_module/_01296_ ),
    .A2(\reg_module/_01297_ ),
    .B1(\reg_module/_01298_ ),
    .Y(\reg_module/_00548_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17909_  (.A(\reg_module/_01284_ ),
    .B(net1589),
    .Y(\reg_module/_01299_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17910_  (.A(\reg_module/_01286_ ),
    .X(\reg_module/_01300_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_17911_  (.A(\reg_module/_01300_ ),
    .X(\reg_module/_01301_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17912_  (.A(\reg_module/_01301_ ),
    .X(\reg_module/_01302_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17913_  (.A(\reg_module/_07677_ ),
    .B(\reg_module/_01302_ ),
    .Y(\reg_module/_01303_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17914_  (.A1(\reg_module/_01299_ ),
    .A2(\reg_module/_01303_ ),
    .B1(\reg_module/_01298_ ),
    .Y(\reg_module/_00549_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17915_  (.A(\reg_module/_01283_ ),
    .X(\reg_module/_01304_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17916_  (.A(\reg_module/_01304_ ),
    .B(net1358),
    .Y(\reg_module/_01305_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17917_  (.A(\reg_module/_07684_ ),
    .B(\reg_module/_01302_ ),
    .Y(\reg_module/_01306_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17918_  (.A1(\reg_module/_01305_ ),
    .A2(\reg_module/_01306_ ),
    .B1(\reg_module/_01298_ ),
    .Y(\reg_module/_00550_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17919_  (.A(\reg_module/_01304_ ),
    .B(net1440),
    .Y(\reg_module/_01307_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17920_  (.A(\reg_module/_07689_ ),
    .B(\reg_module/_01302_ ),
    .Y(\reg_module/_01308_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17921_  (.A1(\reg_module/_01307_ ),
    .A2(\reg_module/_01308_ ),
    .B1(\reg_module/_01298_ ),
    .Y(\reg_module/_00551_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17922_  (.A(\reg_module/_01304_ ),
    .B(net1944),
    .Y(\reg_module/_01309_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17923_  (.A(\reg_module/_07694_ ),
    .B(\reg_module/_01302_ ),
    .Y(\reg_module/_01310_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17924_  (.A1(\reg_module/_01309_ ),
    .A2(\reg_module/_01310_ ),
    .B1(\reg_module/_01298_ ),
    .Y(\reg_module/_00552_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17925_  (.A(\reg_module/_01304_ ),
    .B(net1712),
    .Y(\reg_module/_01311_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17926_  (.A(\reg_module/_07698_ ),
    .B(\reg_module/_01302_ ),
    .Y(\reg_module/_01312_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17927_  (.A1(\reg_module/_01311_ ),
    .A2(\reg_module/_01312_ ),
    .B1(\reg_module/_01298_ ),
    .Y(\reg_module/_00553_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17928_  (.A(\reg_module/_01304_ ),
    .B(net1574),
    .Y(\reg_module/_01313_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17929_  (.A(\reg_module/_07702_ ),
    .B(\reg_module/_01302_ ),
    .Y(\reg_module/_01314_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_17930_  (.A(\reg_module/_09303_ ),
    .X(\reg_module/_01315_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17931_  (.A(\reg_module/_01315_ ),
    .X(\reg_module/_01316_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17932_  (.A1(\reg_module/_01313_ ),
    .A2(\reg_module/_01314_ ),
    .B1(\reg_module/_01316_ ),
    .Y(\reg_module/_00554_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17933_  (.A(\reg_module/_01304_ ),
    .B(net1842),
    .Y(\reg_module/_01317_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17934_  (.A(\reg_module/_01301_ ),
    .X(\reg_module/_01318_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17935_  (.A(\reg_module/_07706_ ),
    .B(\reg_module/_01318_ ),
    .Y(\reg_module/_01319_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17936_  (.A1(\reg_module/_01317_ ),
    .A2(\reg_module/_01319_ ),
    .B1(\reg_module/_01316_ ),
    .Y(\reg_module/_00555_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17937_  (.A(\reg_module/_01283_ ),
    .X(\reg_module/_01320_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17938_  (.A(\reg_module/_01320_ ),
    .B(net2023),
    .Y(\reg_module/_01321_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17939_  (.A(\reg_module/_07713_ ),
    .B(\reg_module/_01318_ ),
    .Y(\reg_module/_01322_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17940_  (.A1(\reg_module/_01321_ ),
    .A2(\reg_module/_01322_ ),
    .B1(\reg_module/_01316_ ),
    .Y(\reg_module/_00556_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17941_  (.A(\reg_module/_01320_ ),
    .B(net1998),
    .Y(\reg_module/_01323_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17942_  (.A(\reg_module/_07718_ ),
    .B(\reg_module/_01318_ ),
    .Y(\reg_module/_01324_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17943_  (.A1(\reg_module/_01323_ ),
    .A2(\reg_module/_01324_ ),
    .B1(\reg_module/_01316_ ),
    .Y(\reg_module/_00557_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17944_  (.A(\reg_module/_01320_ ),
    .B(net2134),
    .Y(\reg_module/_01325_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17945_  (.A(\reg_module/_07723_ ),
    .B(\reg_module/_01318_ ),
    .Y(\reg_module/_01326_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17946_  (.A1(\reg_module/_01325_ ),
    .A2(\reg_module/_01326_ ),
    .B1(\reg_module/_01316_ ),
    .Y(\reg_module/_00558_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17947_  (.A(\reg_module/_01320_ ),
    .B(net1956),
    .Y(\reg_module/_01327_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17948_  (.A(\reg_module/_07727_ ),
    .B(\reg_module/_01318_ ),
    .Y(\reg_module/_01328_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17949_  (.A1(\reg_module/_01327_ ),
    .A2(\reg_module/_01328_ ),
    .B1(\reg_module/_01316_ ),
    .Y(\reg_module/_00559_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17950_  (.A(\reg_module/_01320_ ),
    .B(net2021),
    .Y(\reg_module/_01329_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17951_  (.A(\reg_module/_07731_ ),
    .B(\reg_module/_01318_ ),
    .Y(\reg_module/_01330_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_17952_  (.A(\reg_module/_01315_ ),
    .X(\reg_module/_01331_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17953_  (.A1(\reg_module/_01329_ ),
    .A2(\reg_module/_01330_ ),
    .B1(\reg_module/_01331_ ),
    .Y(\reg_module/_00560_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17954_  (.A(\reg_module/_01320_ ),
    .B(net2097),
    .Y(\reg_module/_01332_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_17955_  (.A(\reg_module/_01301_ ),
    .X(\reg_module/_01333_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17956_  (.A(\reg_module/_07735_ ),
    .B(\reg_module/_01333_ ),
    .Y(\reg_module/_01334_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17957_  (.A1(\reg_module/_01332_ ),
    .A2(\reg_module/_01334_ ),
    .B1(\reg_module/_01331_ ),
    .Y(\reg_module/_00561_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17958_  (.A(\reg_module/_01283_ ),
    .X(\reg_module/_01335_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17959_  (.A(\reg_module/_01335_ ),
    .B(net2014),
    .Y(\reg_module/_01336_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17960_  (.A(\reg_module/_07742_ ),
    .B(\reg_module/_01333_ ),
    .Y(\reg_module/_01337_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17961_  (.A1(\reg_module/_01336_ ),
    .A2(\reg_module/_01337_ ),
    .B1(\reg_module/_01331_ ),
    .Y(\reg_module/_00562_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17962_  (.A(\reg_module/_01335_ ),
    .B(net2007),
    .Y(\reg_module/_01338_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17963_  (.A(\reg_module/_07747_ ),
    .B(\reg_module/_01333_ ),
    .Y(\reg_module/_01339_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17964_  (.A1(\reg_module/_01338_ ),
    .A2(\reg_module/_01339_ ),
    .B1(\reg_module/_01331_ ),
    .Y(\reg_module/_00563_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17965_  (.A(\reg_module/_01335_ ),
    .B(net1980),
    .Y(\reg_module/_01340_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17966_  (.A(\reg_module/_07752_ ),
    .B(\reg_module/_01333_ ),
    .Y(\reg_module/_01341_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17967_  (.A1(\reg_module/_01340_ ),
    .A2(\reg_module/_01341_ ),
    .B1(\reg_module/_01331_ ),
    .Y(\reg_module/_00564_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17968_  (.A(\reg_module/_01335_ ),
    .B(net1999),
    .Y(\reg_module/_01342_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17969_  (.A(\reg_module/_07756_ ),
    .B(\reg_module/_01333_ ),
    .Y(\reg_module/_01343_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17970_  (.A1(\reg_module/_01342_ ),
    .A2(\reg_module/_01343_ ),
    .B1(\reg_module/_01331_ ),
    .Y(\reg_module/_00565_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17971_  (.A(\reg_module/_01335_ ),
    .B(net1972),
    .Y(\reg_module/_01344_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17972_  (.A(\reg_module/_07760_ ),
    .B(\reg_module/_01333_ ),
    .Y(\reg_module/_01345_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17973_  (.A(\reg_module/_01315_ ),
    .X(\reg_module/_01346_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17974_  (.A1(\reg_module/_01344_ ),
    .A2(\reg_module/_01345_ ),
    .B1(\reg_module/_01346_ ),
    .Y(\reg_module/_00566_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17975_  (.A(\reg_module/_01335_ ),
    .B(net1860),
    .Y(\reg_module/_01347_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_17976_  (.A(\reg_module/_01300_ ),
    .X(\reg_module/_01348_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17977_  (.A(\reg_module/_01348_ ),
    .X(\reg_module/_01349_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17978_  (.A(\reg_module/_07764_ ),
    .B(\reg_module/_01349_ ),
    .Y(\reg_module/_01350_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17979_  (.A1(\reg_module/_01347_ ),
    .A2(\reg_module/_01350_ ),
    .B1(\reg_module/_01346_ ),
    .Y(\reg_module/_00567_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_17980_  (.A(\reg_module/_01282_ ),
    .X(\reg_module/_01351_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17981_  (.A(\reg_module/_01351_ ),
    .B(net1443),
    .Y(\reg_module/_01352_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17982_  (.A(\reg_module/_07772_ ),
    .B(\reg_module/_01349_ ),
    .Y(\reg_module/_01353_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17983_  (.A1(\reg_module/_01352_ ),
    .A2(\reg_module/_01353_ ),
    .B1(\reg_module/_01346_ ),
    .Y(\reg_module/_00568_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17984_  (.A(\reg_module/_01351_ ),
    .B(net1309),
    .Y(\reg_module/_01354_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17985_  (.A(\reg_module/_07778_ ),
    .B(\reg_module/_01349_ ),
    .Y(\reg_module/_01355_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17986_  (.A1(\reg_module/_01354_ ),
    .A2(\reg_module/_01355_ ),
    .B1(\reg_module/_01346_ ),
    .Y(\reg_module/_00569_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17987_  (.A(\reg_module/_01351_ ),
    .B(net1824),
    .Y(\reg_module/_01356_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17988_  (.A(\reg_module/_07784_ ),
    .B(\reg_module/_01349_ ),
    .Y(\reg_module/_01357_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17989_  (.A1(\reg_module/_01356_ ),
    .A2(\reg_module/_01357_ ),
    .B1(\reg_module/_01346_ ),
    .Y(\reg_module/_00570_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17990_  (.A(\reg_module/_01351_ ),
    .B(net1896),
    .Y(\reg_module/_01358_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17991_  (.A(\reg_module/_07788_ ),
    .B(\reg_module/_01349_ ),
    .Y(\reg_module/_01359_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17992_  (.A1(\reg_module/_01358_ ),
    .A2(\reg_module/_01359_ ),
    .B1(\reg_module/_01346_ ),
    .Y(\reg_module/_00571_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17993_  (.A(\reg_module/_01351_ ),
    .B(net1516),
    .Y(\reg_module/_01360_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17994_  (.A(\reg_module/_07792_ ),
    .B(\reg_module/_01349_ ),
    .Y(\reg_module/_01361_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_17995_  (.A(\reg_module/_01315_ ),
    .X(\reg_module/_01362_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_17996_  (.A1(\reg_module/_01360_ ),
    .A2(\reg_module/_01361_ ),
    .B1(\reg_module/_01362_ ),
    .Y(\reg_module/_00572_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17997_  (.A(\reg_module/_01351_ ),
    .B(net1636),
    .Y(\reg_module/_01363_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_17998_  (.A(\reg_module/_01348_ ),
    .X(\reg_module/_01364_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_17999_  (.A(\reg_module/_07796_ ),
    .B(\reg_module/_01364_ ),
    .Y(\reg_module/_01365_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18000_  (.A1(\reg_module/_01363_ ),
    .A2(\reg_module/_01365_ ),
    .B1(\reg_module/_01362_ ),
    .Y(\reg_module/_00573_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18001_  (.A(\reg_module/_01283_ ),
    .B(net1284),
    .Y(\reg_module/_01366_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18002_  (.A(\reg_module/_07801_ ),
    .B(\reg_module/_01364_ ),
    .Y(\reg_module/_01367_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18003_  (.A1(\reg_module/_01366_ ),
    .A2(\reg_module/_01367_ ),
    .B1(\reg_module/_01362_ ),
    .Y(\reg_module/_00574_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18004_  (.A(\reg_module/_01283_ ),
    .B(net1271),
    .Y(\reg_module/_01368_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18005_  (.A(\reg_module/_07806_ ),
    .B(\reg_module/_01364_ ),
    .Y(\reg_module/_01369_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18006_  (.A1(\reg_module/_01368_ ),
    .A2(\reg_module/_01369_ ),
    .B1(\reg_module/_01362_ ),
    .Y(\reg_module/_00575_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18007_  (.A(\reg_module/_01281_ ),
    .B(\reg_module/_07810_ ),
    .Y(\reg_module/_01370_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_18008_  (.A(\reg_module/_01370_ ),
    .X(\reg_module/_01371_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18009_  (.A(\reg_module/_01371_ ),
    .X(\reg_module/_01372_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18010_  (.A(\reg_module/_01372_ ),
    .B(net1652),
    .Y(\reg_module/_01373_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18011_  (.A(\reg_module/_07823_ ),
    .B(\reg_module/_01364_ ),
    .Y(\reg_module/_01374_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18012_  (.A1(\reg_module/_01373_ ),
    .A2(\reg_module/_01374_ ),
    .B1(\reg_module/_01362_ ),
    .Y(\reg_module/_00576_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18013_  (.A(\reg_module/_01372_ ),
    .B(net1960),
    .Y(\reg_module/_01375_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18014_  (.A(\reg_module/_07828_ ),
    .B(\reg_module/_01364_ ),
    .Y(\reg_module/_01376_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18015_  (.A1(\reg_module/_01375_ ),
    .A2(\reg_module/_01376_ ),
    .B1(\reg_module/_01362_ ),
    .Y(\reg_module/_00577_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18016_  (.A(\reg_module/_01372_ ),
    .B(net1655),
    .Y(\reg_module/_01377_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18017_  (.A(\reg_module/_07833_ ),
    .B(\reg_module/_01364_ ),
    .Y(\reg_module/_01378_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18018_  (.A(\reg_module/_01315_ ),
    .X(\reg_module/_01379_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18019_  (.A1(\reg_module/_01377_ ),
    .A2(\reg_module/_01378_ ),
    .B1(\reg_module/_01379_ ),
    .Y(\reg_module/_00578_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18020_  (.A(\reg_module/_01372_ ),
    .B(net1614),
    .Y(\reg_module/_01380_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18021_  (.A(\reg_module/_01281_ ),
    .X(\reg_module/_01381_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_18022_  (.A(\reg_module/_01381_ ),
    .X(\reg_module/_01382_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18023_  (.A(\reg_module/_07838_ ),
    .B(\reg_module/_01382_ ),
    .Y(\reg_module/_01383_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18024_  (.A1(\reg_module/_01380_ ),
    .A2(\reg_module/_01383_ ),
    .B1(\reg_module/_01379_ ),
    .Y(\reg_module/_00579_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18025_  (.A(\reg_module/_01372_ ),
    .B(net1724),
    .Y(\reg_module/_01384_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18026_  (.A(\reg_module/_01348_ ),
    .X(\reg_module/_01385_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18027_  (.A(\reg_module/_07846_ ),
    .B(\reg_module/_01385_ ),
    .Y(\reg_module/_01386_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18028_  (.A1(\reg_module/_01384_ ),
    .A2(\reg_module/_01386_ ),
    .B1(\reg_module/_01379_ ),
    .Y(\reg_module/_00580_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18029_  (.A(\reg_module/_01372_ ),
    .B(net1814),
    .Y(\reg_module/_01387_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18030_  (.A(\reg_module/_07852_ ),
    .B(\reg_module/_01385_ ),
    .Y(\reg_module/_01388_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18031_  (.A1(\reg_module/_01387_ ),
    .A2(\reg_module/_01388_ ),
    .B1(\reg_module/_01379_ ),
    .Y(\reg_module/_00581_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18032_  (.A(\reg_module/_01371_ ),
    .X(\reg_module/_01389_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18033_  (.A(\reg_module/_01389_ ),
    .B(net1830),
    .Y(\reg_module/_01390_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18034_  (.A(\reg_module/_07860_ ),
    .B(\reg_module/_01385_ ),
    .Y(\reg_module/_01391_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18035_  (.A1(\reg_module/_01390_ ),
    .A2(\reg_module/_01391_ ),
    .B1(\reg_module/_01379_ ),
    .Y(\reg_module/_00582_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18036_  (.A(\reg_module/_01389_ ),
    .B(net1616),
    .Y(\reg_module/_01392_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18037_  (.A(\reg_module/_07865_ ),
    .B(\reg_module/_01385_ ),
    .Y(\reg_module/_01393_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18038_  (.A1(\reg_module/_01392_ ),
    .A2(\reg_module/_01393_ ),
    .B1(\reg_module/_01379_ ),
    .Y(\reg_module/_00583_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18039_  (.A(\reg_module/_01389_ ),
    .B(net2182),
    .Y(\reg_module/_01394_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18040_  (.A(\reg_module/_07870_ ),
    .B(\reg_module/_01385_ ),
    .Y(\reg_module/_01395_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18041_  (.A(\reg_module/_01315_ ),
    .X(\reg_module/_01396_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18042_  (.A1(\reg_module/_01394_ ),
    .A2(\reg_module/_01395_ ),
    .B1(\reg_module/_01396_ ),
    .Y(\reg_module/_00584_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18043_  (.A(\reg_module/_01389_ ),
    .B(net1749),
    .Y(\reg_module/_01397_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18044_  (.A(\reg_module/_07875_ ),
    .B(\reg_module/_01385_ ),
    .Y(\reg_module/_01398_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18045_  (.A1(\reg_module/_01397_ ),
    .A2(\reg_module/_01398_ ),
    .B1(\reg_module/_01396_ ),
    .Y(\reg_module/_00585_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18046_  (.A(\reg_module/_01389_ ),
    .B(net1687),
    .Y(\reg_module/_01399_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18047_  (.A(\reg_module/_07882_ ),
    .B(\reg_module/_01382_ ),
    .Y(\reg_module/_01400_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18048_  (.A1(\reg_module/_01399_ ),
    .A2(\reg_module/_01400_ ),
    .B1(\reg_module/_01396_ ),
    .Y(\reg_module/_00586_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18049_  (.A(\reg_module/_01389_ ),
    .B(net2107),
    .Y(\reg_module/_01401_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18050_  (.A(\reg_module/_01348_ ),
    .X(\reg_module/_01402_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18051_  (.A(\reg_module/_07888_ ),
    .B(\reg_module/_01402_ ),
    .Y(\reg_module/_01403_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18052_  (.A1(\reg_module/_01401_ ),
    .A2(\reg_module/_01403_ ),
    .B1(\reg_module/_01396_ ),
    .Y(\reg_module/_00587_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18053_  (.A(\reg_module/_01371_ ),
    .X(\reg_module/_01404_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18054_  (.A(\reg_module/_01404_ ),
    .B(net1669),
    .Y(\reg_module/_01405_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18055_  (.A(\reg_module/_07896_ ),
    .B(\reg_module/_01402_ ),
    .Y(\reg_module/_01406_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18056_  (.A1(\reg_module/_01405_ ),
    .A2(\reg_module/_01406_ ),
    .B1(\reg_module/_01396_ ),
    .Y(\reg_module/_00588_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18057_  (.A(\reg_module/_01404_ ),
    .B(net1466),
    .Y(\reg_module/_01407_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_18058_  (.A(\reg_module/_01381_ ),
    .X(\reg_module/_01408_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18059_  (.A(\reg_module/_07901_ ),
    .B(\reg_module/_01408_ ),
    .Y(\reg_module/_01409_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18060_  (.A1(\reg_module/_01407_ ),
    .A2(\reg_module/_01409_ ),
    .B1(\reg_module/_01396_ ),
    .Y(\reg_module/_00589_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18061_  (.A(\reg_module/_01404_ ),
    .B(net1943),
    .Y(\reg_module/_01410_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18062_  (.A(\reg_module/_07906_ ),
    .B(\reg_module/_01402_ ),
    .Y(\reg_module/_01411_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_18063_  (.A(\reg_module/_09303_ ),
    .X(\reg_module/_01412_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18064_  (.A(\reg_module/_01412_ ),
    .X(\reg_module/_01413_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18065_  (.A1(\reg_module/_01410_ ),
    .A2(\reg_module/_01411_ ),
    .B1(\reg_module/_01413_ ),
    .Y(\reg_module/_00590_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18066_  (.A(\reg_module/_01404_ ),
    .B(net1445),
    .Y(\reg_module/_01414_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18067_  (.A(\reg_module/_07911_ ),
    .B(\reg_module/_01402_ ),
    .Y(\reg_module/_01415_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18068_  (.A1(\reg_module/_01414_ ),
    .A2(\reg_module/_01415_ ),
    .B1(\reg_module/_01413_ ),
    .Y(\reg_module/_00591_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18069_  (.A(\reg_module/_01404_ ),
    .B(net1594),
    .Y(\reg_module/_01416_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18070_  (.A(\reg_module/_07918_ ),
    .B(\reg_module/_01402_ ),
    .Y(\reg_module/_01417_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18071_  (.A1(\reg_module/_01416_ ),
    .A2(\reg_module/_01417_ ),
    .B1(\reg_module/_01413_ ),
    .Y(\reg_module/_00592_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18072_  (.A(\reg_module/_01404_ ),
    .B(net2011),
    .Y(\reg_module/_01418_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18073_  (.A(\reg_module/_07924_ ),
    .B(\reg_module/_01402_ ),
    .Y(\reg_module/_01419_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18074_  (.A1(\reg_module/_01418_ ),
    .A2(\reg_module/_01419_ ),
    .B1(\reg_module/_01413_ ),
    .Y(\reg_module/_00593_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18075_  (.A(\reg_module/_01371_ ),
    .X(\reg_module/_01420_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18076_  (.A(\reg_module/_01420_ ),
    .B(net1446),
    .Y(\reg_module/_01421_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18077_  (.A(\reg_module/_07932_ ),
    .B(\reg_module/_01408_ ),
    .Y(\reg_module/_01422_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18078_  (.A1(\reg_module/_01421_ ),
    .A2(\reg_module/_01422_ ),
    .B1(\reg_module/_01413_ ),
    .Y(\reg_module/_00594_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18079_  (.A(\reg_module/_01420_ ),
    .B(net1485),
    .Y(\reg_module/_01423_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18080_  (.A(\reg_module/_01348_ ),
    .X(\reg_module/_01424_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18081_  (.A(\reg_module/_07937_ ),
    .B(\reg_module/_01424_ ),
    .Y(\reg_module/_01425_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18082_  (.A1(\reg_module/_01423_ ),
    .A2(\reg_module/_01425_ ),
    .B1(\reg_module/_01413_ ),
    .Y(\reg_module/_00595_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18083_  (.A(\reg_module/_01420_ ),
    .B(net1695),
    .Y(\reg_module/_01426_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18084_  (.A(\reg_module/_07942_ ),
    .B(\reg_module/_01424_ ),
    .Y(\reg_module/_01427_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18085_  (.A(\reg_module/_01412_ ),
    .X(\reg_module/_01428_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18086_  (.A1(\reg_module/_01426_ ),
    .A2(\reg_module/_01427_ ),
    .B1(\reg_module/_01428_ ),
    .Y(\reg_module/_00596_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18087_  (.A(\reg_module/_01420_ ),
    .B(net1618),
    .Y(\reg_module/_01429_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18088_  (.A(\reg_module/_07947_ ),
    .B(\reg_module/_01424_ ),
    .Y(\reg_module/_01430_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18089_  (.A1(\reg_module/_01429_ ),
    .A2(\reg_module/_01430_ ),
    .B1(\reg_module/_01428_ ),
    .Y(\reg_module/_00597_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18090_  (.A(\reg_module/_01420_ ),
    .B(net1700),
    .Y(\reg_module/_01431_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18091_  (.A(\reg_module/_07954_ ),
    .B(\reg_module/_01424_ ),
    .Y(\reg_module/_01432_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18092_  (.A1(\reg_module/_01431_ ),
    .A2(\reg_module/_01432_ ),
    .B1(\reg_module/_01428_ ),
    .Y(\reg_module/_00598_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18093_  (.A(\reg_module/_01420_ ),
    .B(net1690),
    .Y(\reg_module/_01433_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18094_  (.A(\reg_module/_07960_ ),
    .B(\reg_module/_01408_ ),
    .Y(\reg_module/_01434_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18095_  (.A1(\reg_module/_01433_ ),
    .A2(\reg_module/_01434_ ),
    .B1(\reg_module/_01428_ ),
    .Y(\reg_module/_00599_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18096_  (.A(\reg_module/_01370_ ),
    .X(\reg_module/_01435_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18097_  (.A(\reg_module/_01435_ ),
    .B(net1833),
    .Y(\reg_module/_01436_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18098_  (.A(\reg_module/_07968_ ),
    .B(\reg_module/_01424_ ),
    .Y(\reg_module/_01437_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18099_  (.A1(\reg_module/_01436_ ),
    .A2(\reg_module/_01437_ ),
    .B1(\reg_module/_01428_ ),
    .Y(\reg_module/_00600_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18100_  (.A(\reg_module/_01435_ ),
    .B(net1939),
    .Y(\reg_module/_01438_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18101_  (.A(\reg_module/_07973_ ),
    .B(\reg_module/_01424_ ),
    .Y(\reg_module/_01439_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18102_  (.A1(\reg_module/_01438_ ),
    .A2(\reg_module/_01439_ ),
    .B1(\reg_module/_01428_ ),
    .Y(\reg_module/_00601_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18103_  (.A(\reg_module/_01435_ ),
    .B(net1932),
    .Y(\reg_module/_01440_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18104_  (.A(\reg_module/_01348_ ),
    .X(\reg_module/_01441_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18105_  (.A(\reg_module/_07978_ ),
    .B(\reg_module/_01441_ ),
    .Y(\reg_module/_01442_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18106_  (.A(\reg_module/_01412_ ),
    .X(\reg_module/_01443_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18107_  (.A1(\reg_module/_01440_ ),
    .A2(\reg_module/_01442_ ),
    .B1(\reg_module/_01443_ ),
    .Y(\reg_module/_00602_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18108_  (.A(\reg_module/_01435_ ),
    .B(net1992),
    .Y(\reg_module/_01444_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18109_  (.A(\reg_module/_07983_ ),
    .B(\reg_module/_01441_ ),
    .Y(\reg_module/_01445_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18110_  (.A1(\reg_module/_01444_ ),
    .A2(\reg_module/_01445_ ),
    .B1(\reg_module/_01443_ ),
    .Y(\reg_module/_00603_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18111_  (.A(\reg_module/_01435_ ),
    .B(net1839),
    .Y(\reg_module/_01446_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18112_  (.A(\reg_module/_07991_ ),
    .B(\reg_module/_01441_ ),
    .Y(\reg_module/_01447_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18113_  (.A1(\reg_module/_01446_ ),
    .A2(\reg_module/_01447_ ),
    .B1(\reg_module/_01443_ ),
    .Y(\reg_module/_00604_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18114_  (.A(\reg_module/_01435_ ),
    .B(net2054),
    .Y(\reg_module/_01448_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18115_  (.A(\reg_module/_07999_ ),
    .B(\reg_module/_01441_ ),
    .Y(\reg_module/_01449_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18116_  (.A1(\reg_module/_01448_ ),
    .A2(\reg_module/_01449_ ),
    .B1(\reg_module/_01443_ ),
    .Y(\reg_module/_00605_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18117_  (.A(\reg_module/_01371_ ),
    .B(net1703),
    .Y(\reg_module/_01450_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18118_  (.A(\reg_module/_08005_ ),
    .B(\reg_module/_01441_ ),
    .Y(\reg_module/_01451_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18119_  (.A1(\reg_module/_01450_ ),
    .A2(\reg_module/_01451_ ),
    .B1(\reg_module/_01443_ ),
    .Y(\reg_module/_00606_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18120_  (.A(\reg_module/_01371_ ),
    .B(net1639),
    .Y(\reg_module/_01452_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18121_  (.A(\reg_module/_08010_ ),
    .B(\reg_module/_01441_ ),
    .Y(\reg_module/_01453_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18122_  (.A1(\reg_module/_01452_ ),
    .A2(\reg_module/_01453_ ),
    .B1(\reg_module/_01443_ ),
    .Y(\reg_module/_00607_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18123_  (.A(\reg_module/_01281_ ),
    .B(\reg_module/_08015_ ),
    .Y(\reg_module/_01454_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_18124_  (.A(\reg_module/_01454_ ),
    .X(\reg_module/_01455_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18125_  (.A(\reg_module/_01455_ ),
    .X(\reg_module/_01456_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18126_  (.A(\reg_module/_01456_ ),
    .B(net1846),
    .Y(\reg_module/_01457_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18127_  (.A(\reg_module/_01300_ ),
    .X(\reg_module/_01458_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18128_  (.A(\reg_module/_01458_ ),
    .X(\reg_module/_01459_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18129_  (.A(\reg_module/_08024_ ),
    .B(\reg_module/_01459_ ),
    .Y(\reg_module/_01460_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18130_  (.A(\reg_module/_01412_ ),
    .X(\reg_module/_01461_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18131_  (.A1(\reg_module/_01457_ ),
    .A2(\reg_module/_01460_ ),
    .B1(\reg_module/_01461_ ),
    .Y(\reg_module/_00608_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18132_  (.A(\reg_module/_01456_ ),
    .B(net1511),
    .Y(\reg_module/_01462_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18133_  (.A(\reg_module/_08030_ ),
    .B(\reg_module/_01459_ ),
    .Y(\reg_module/_01463_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18134_  (.A1(\reg_module/_01462_ ),
    .A2(\reg_module/_01463_ ),
    .B1(\reg_module/_01461_ ),
    .Y(\reg_module/_00609_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18135_  (.A(\reg_module/_01456_ ),
    .B(net1905),
    .Y(\reg_module/_01464_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18136_  (.A(\reg_module/_08035_ ),
    .B(\reg_module/_01459_ ),
    .Y(\reg_module/_01465_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18137_  (.A1(\reg_module/_01464_ ),
    .A2(\reg_module/_01465_ ),
    .B1(\reg_module/_01461_ ),
    .Y(\reg_module/_00610_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18138_  (.A(\reg_module/_01456_ ),
    .B(net1361),
    .Y(\reg_module/_01466_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18139_  (.A(\reg_module/_08040_ ),
    .B(\reg_module/_01459_ ),
    .Y(\reg_module/_01467_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18140_  (.A1(\reg_module/_01466_ ),
    .A2(\reg_module/_01467_ ),
    .B1(\reg_module/_01461_ ),
    .Y(\reg_module/_00611_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18141_  (.A(\reg_module/_01456_ ),
    .B(net1256),
    .Y(\reg_module/_01468_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18142_  (.A(\reg_module/_08044_ ),
    .B(\reg_module/_01459_ ),
    .Y(\reg_module/_01469_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18143_  (.A1(\reg_module/_01468_ ),
    .A2(\reg_module/_01469_ ),
    .B1(\reg_module/_01461_ ),
    .Y(\reg_module/_00612_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18144_  (.A(\reg_module/_01456_ ),
    .B(net1427),
    .Y(\reg_module/_01470_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18145_  (.A(\reg_module/_01408_ ),
    .X(\reg_module/_01471_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18146_  (.A(\reg_module/_01471_ ),
    .B(\reg_module/_08048_ ),
    .Y(\reg_module/_01472_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18147_  (.A1(\reg_module/_01470_ ),
    .A2(\reg_module/_01472_ ),
    .B1(\reg_module/_01461_ ),
    .Y(\reg_module/_00613_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18148_  (.A(\reg_module/_01455_ ),
    .X(\reg_module/_01473_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18149_  (.A(\reg_module/_01473_ ),
    .B(net1441),
    .Y(\reg_module/_01474_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18150_  (.A(\reg_module/_08054_ ),
    .B(\reg_module/_01459_ ),
    .Y(\reg_module/_01475_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18151_  (.A(\reg_module/_01412_ ),
    .X(\reg_module/_01476_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18152_  (.A1(\reg_module/_01474_ ),
    .A2(\reg_module/_01475_ ),
    .B1(\reg_module/_01476_ ),
    .Y(\reg_module/_00614_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18153_  (.A(\reg_module/_01473_ ),
    .B(net1240),
    .Y(\reg_module/_01477_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18154_  (.A(\reg_module/_01458_ ),
    .X(\reg_module/_01478_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18155_  (.A(\reg_module/_08058_ ),
    .B(\reg_module/_01478_ ),
    .Y(\reg_module/_01479_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18156_  (.A1(\reg_module/_01477_ ),
    .A2(\reg_module/_01479_ ),
    .B1(\reg_module/_01476_ ),
    .Y(\reg_module/_00615_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18157_  (.A(\reg_module/_01473_ ),
    .B(net2056),
    .Y(\reg_module/_01480_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18158_  (.A(\reg_module/_08064_ ),
    .B(\reg_module/_01478_ ),
    .Y(\reg_module/_01481_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18159_  (.A1(\reg_module/_01480_ ),
    .A2(\reg_module/_01481_ ),
    .B1(\reg_module/_01476_ ),
    .Y(\reg_module/_00616_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18160_  (.A(\reg_module/_01473_ ),
    .B(net1251),
    .Y(\reg_module/_01482_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18161_  (.A(\reg_module/_08069_ ),
    .B(\reg_module/_01478_ ),
    .Y(\reg_module/_01483_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18162_  (.A1(\reg_module/_01482_ ),
    .A2(\reg_module/_01483_ ),
    .B1(\reg_module/_01476_ ),
    .Y(\reg_module/_00617_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18163_  (.A(\reg_module/_01473_ ),
    .B(net1291),
    .Y(\reg_module/_01484_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18164_  (.A(\reg_module/_08073_ ),
    .B(\reg_module/_01478_ ),
    .Y(\reg_module/_01485_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18165_  (.A1(\reg_module/_01484_ ),
    .A2(\reg_module/_01485_ ),
    .B1(\reg_module/_01476_ ),
    .Y(\reg_module/_00618_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18166_  (.A(\reg_module/_01473_ ),
    .B(net1836),
    .Y(\reg_module/_01486_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18167_  (.A(\reg_module/_08077_ ),
    .B(\reg_module/_01478_ ),
    .Y(\reg_module/_01487_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18168_  (.A1(\reg_module/_01486_ ),
    .A2(\reg_module/_01487_ ),
    .B1(\reg_module/_01476_ ),
    .Y(\reg_module/_00619_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18169_  (.A(\reg_module/_01455_ ),
    .X(\reg_module/_01488_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18170_  (.A(\reg_module/_01488_ ),
    .B(net1454),
    .Y(\reg_module/_01489_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18171_  (.A(\reg_module/_01471_ ),
    .B(\reg_module/_08083_ ),
    .Y(\reg_module/_01490_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18172_  (.A(\reg_module/_01412_ ),
    .X(\reg_module/_01491_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18173_  (.A1(\reg_module/_01489_ ),
    .A2(\reg_module/_01490_ ),
    .B1(\reg_module/_01491_ ),
    .Y(\reg_module/_00620_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18174_  (.A(\reg_module/_01488_ ),
    .B(net1282),
    .Y(\reg_module/_01492_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18175_  (.A(\reg_module/_08087_ ),
    .B(\reg_module/_01478_ ),
    .Y(\reg_module/_01493_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18176_  (.A1(\reg_module/_01492_ ),
    .A2(\reg_module/_01493_ ),
    .B1(\reg_module/_01491_ ),
    .Y(\reg_module/_00621_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18177_  (.A(\reg_module/_01488_ ),
    .B(net1780),
    .Y(\reg_module/_01494_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18178_  (.A(\reg_module/_01458_ ),
    .X(\reg_module/_01495_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18179_  (.A(\reg_module/_08092_ ),
    .B(\reg_module/_01495_ ),
    .Y(\reg_module/_01496_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18180_  (.A1(\reg_module/_01494_ ),
    .A2(\reg_module/_01496_ ),
    .B1(\reg_module/_01491_ ),
    .Y(\reg_module/_00622_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18181_  (.A(\reg_module/_01488_ ),
    .B(net1330),
    .Y(\reg_module/_01497_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18182_  (.A(\reg_module/_08098_ ),
    .B(\reg_module/_01495_ ),
    .Y(\reg_module/_01498_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18183_  (.A1(\reg_module/_01497_ ),
    .A2(\reg_module/_01498_ ),
    .B1(\reg_module/_01491_ ),
    .Y(\reg_module/_00623_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18184_  (.A(\reg_module/_01488_ ),
    .B(net1263),
    .Y(\reg_module/_01499_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18185_  (.A(\reg_module/_08102_ ),
    .B(\reg_module/_01495_ ),
    .Y(\reg_module/_01500_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18186_  (.A1(\reg_module/_01499_ ),
    .A2(\reg_module/_01500_ ),
    .B1(\reg_module/_01491_ ),
    .Y(\reg_module/_00624_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18187_  (.A(\reg_module/_01488_ ),
    .B(net1890),
    .Y(\reg_module/_01501_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18188_  (.A(\reg_module/_08106_ ),
    .B(\reg_module/_01495_ ),
    .Y(\reg_module/_01502_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18189_  (.A1(\reg_module/_01501_ ),
    .A2(\reg_module/_01502_ ),
    .B1(\reg_module/_01491_ ),
    .Y(\reg_module/_00625_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18190_  (.A(\reg_module/_01455_ ),
    .X(\reg_module/_01503_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18191_  (.A(\reg_module/_01503_ ),
    .B(net1704),
    .Y(\reg_module/_01504_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18192_  (.A(\reg_module/_08112_ ),
    .B(\reg_module/_01495_ ),
    .Y(\reg_module/_01505_ ));
 sky130_fd_sc_hd__buf_1 \reg_module/_18193_  (.A(\reg_module/_07653_ ),
    .X(\reg_module/_01506_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18194_  (.A(\reg_module/_01506_ ),
    .X(\reg_module/_01507_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18195_  (.A(\reg_module/_01507_ ),
    .X(\reg_module/_01508_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18196_  (.A1(\reg_module/_01504_ ),
    .A2(\reg_module/_01505_ ),
    .B1(\reg_module/_01508_ ),
    .Y(\reg_module/_00626_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18197_  (.A(\reg_module/_01503_ ),
    .B(net1731),
    .Y(\reg_module/_01509_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18198_  (.A(\reg_module/_08116_ ),
    .B(\reg_module/_01495_ ),
    .Y(\reg_module/_01510_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18199_  (.A1(\reg_module/_01509_ ),
    .A2(\reg_module/_01510_ ),
    .B1(\reg_module/_01508_ ),
    .Y(\reg_module/_00627_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18200_  (.A(\reg_module/_01503_ ),
    .B(net1629),
    .Y(\reg_module/_01511_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18201_  (.A(\reg_module/_01458_ ),
    .X(\reg_module/_01512_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18202_  (.A(\reg_module/_08121_ ),
    .B(\reg_module/_01512_ ),
    .Y(\reg_module/_01513_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18203_  (.A1(\reg_module/_01511_ ),
    .A2(\reg_module/_01513_ ),
    .B1(\reg_module/_01508_ ),
    .Y(\reg_module/_00628_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18204_  (.A(\reg_module/_01503_ ),
    .B(net1682),
    .Y(\reg_module/_01514_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18205_  (.A(\reg_module/_08127_ ),
    .B(\reg_module/_01512_ ),
    .Y(\reg_module/_01515_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18206_  (.A1(\reg_module/_01514_ ),
    .A2(\reg_module/_01515_ ),
    .B1(\reg_module/_01508_ ),
    .Y(\reg_module/_00629_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18207_  (.A(\reg_module/_01503_ ),
    .B(net1696),
    .Y(\reg_module/_01516_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18208_  (.A(\reg_module/_08131_ ),
    .B(\reg_module/_01512_ ),
    .Y(\reg_module/_01517_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18209_  (.A1(\reg_module/_01516_ ),
    .A2(\reg_module/_01517_ ),
    .B1(\reg_module/_01508_ ),
    .Y(\reg_module/_00630_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18210_  (.A(\reg_module/_01503_ ),
    .B(net1595),
    .Y(\reg_module/_01518_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18211_  (.A(\reg_module/_08135_ ),
    .B(\reg_module/_01512_ ),
    .Y(\reg_module/_01519_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18212_  (.A1(\reg_module/_01518_ ),
    .A2(\reg_module/_01519_ ),
    .B1(\reg_module/_01508_ ),
    .Y(\reg_module/_00631_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18213_  (.A(\reg_module/_01454_ ),
    .X(\reg_module/_01520_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18214_  (.A(\reg_module/_01520_ ),
    .B(net1299),
    .Y(\reg_module/_01521_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18215_  (.A(\reg_module/_08141_ ),
    .B(\reg_module/_01512_ ),
    .Y(\reg_module/_01522_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18216_  (.A(\reg_module/_01507_ ),
    .X(\reg_module/_01523_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18217_  (.A1(\reg_module/_01521_ ),
    .A2(\reg_module/_01522_ ),
    .B1(\reg_module/_01523_ ),
    .Y(\reg_module/_00632_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18218_  (.A(\reg_module/_01520_ ),
    .B(net1232),
    .Y(\reg_module/_01524_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18219_  (.A(\reg_module/_08145_ ),
    .B(\reg_module/_01512_ ),
    .Y(\reg_module/_01525_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18220_  (.A1(\reg_module/_01524_ ),
    .A2(\reg_module/_01525_ ),
    .B1(\reg_module/_01523_ ),
    .Y(\reg_module/_00633_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18221_  (.A(\reg_module/_01520_ ),
    .B(net1638),
    .Y(\reg_module/_01526_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18222_  (.A(\reg_module/_01458_ ),
    .X(\reg_module/_01527_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18223_  (.A(\reg_module/_08150_ ),
    .B(\reg_module/_01527_ ),
    .Y(\reg_module/_01528_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18224_  (.A1(\reg_module/_01526_ ),
    .A2(\reg_module/_01528_ ),
    .B1(\reg_module/_01523_ ),
    .Y(\reg_module/_00634_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18225_  (.A(\reg_module/_01520_ ),
    .B(net1376),
    .Y(\reg_module/_01529_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18226_  (.A(\reg_module/_08155_ ),
    .B(\reg_module/_01527_ ),
    .Y(\reg_module/_01530_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18227_  (.A1(\reg_module/_01529_ ),
    .A2(\reg_module/_01530_ ),
    .B1(\reg_module/_01523_ ),
    .Y(\reg_module/_00635_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18228_  (.A(\reg_module/_01520_ ),
    .B(net1304),
    .Y(\reg_module/_01531_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18229_  (.A(\reg_module/_01471_ ),
    .B(\reg_module/_08159_ ),
    .Y(\reg_module/_01532_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18230_  (.A1(\reg_module/_01531_ ),
    .A2(\reg_module/_01532_ ),
    .B1(\reg_module/_01523_ ),
    .Y(\reg_module/_00636_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18231_  (.A(\reg_module/_01520_ ),
    .B(net1554),
    .Y(\reg_module/_01533_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18232_  (.A(\reg_module/_08163_ ),
    .B(\reg_module/_01527_ ),
    .Y(\reg_module/_01534_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18233_  (.A1(\reg_module/_01533_ ),
    .A2(\reg_module/_01534_ ),
    .B1(\reg_module/_01523_ ),
    .Y(\reg_module/_00637_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18234_  (.A(\reg_module/_01455_ ),
    .B(net1293),
    .Y(\reg_module/_01535_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18235_  (.A(\reg_module/_08167_ ),
    .B(\reg_module/_01527_ ),
    .Y(\reg_module/_01536_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18236_  (.A(\reg_module/_01507_ ),
    .X(\reg_module/_01537_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18237_  (.A1(\reg_module/_01535_ ),
    .A2(\reg_module/_01536_ ),
    .B1(\reg_module/_01537_ ),
    .Y(\reg_module/_00638_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18238_  (.A(\reg_module/_01455_ ),
    .B(net1388),
    .Y(\reg_module/_01538_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18239_  (.A(\reg_module/_08171_ ),
    .B(\reg_module/_01527_ ),
    .Y(\reg_module/_01539_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18240_  (.A1(\reg_module/_01538_ ),
    .A2(\reg_module/_01539_ ),
    .B1(\reg_module/_01537_ ),
    .Y(\reg_module/_00639_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18241_  (.A(\reg_module/_08175_ ),
    .B(\reg_module/_01153_ ),
    .Y(\reg_module/_01540_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18242_  (.A(\reg_module/_01540_ ),
    .X(\reg_module/_01541_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18243_  (.A(\reg_module/_01541_ ),
    .X(\reg_module/_01542_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18244_  (.A(net1774),
    .B(\reg_module/_01542_ ),
    .Y(\reg_module/_01543_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18245_  (.A(\reg_module/_01540_ ),
    .X(\reg_module/_01544_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18246_  (.A(\reg_module/_07653_ ),
    .X(\reg_module/_01545_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18247_  (.A(\reg_module/_01545_ ),
    .X(\reg_module/_01546_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18248_  (.A1(\reg_module/_01544_ ),
    .A2(\reg_module/_07513_ ),
    .B1(\reg_module/_01546_ ),
    .X(\reg_module/_01547_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18249_  (.A(\reg_module/_01543_ ),
    .B(\reg_module/_01547_ ),
    .Y(\reg_module/_00640_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18250_  (.A(\reg_module/_01540_ ),
    .X(\reg_module/_01548_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18251_  (.A(\reg_module/_01548_ ),
    .X(\reg_module/_01549_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18252_  (.A(net2193),
    .B(\reg_module/_01549_ ),
    .Y(\reg_module/_01550_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18253_  (.A(\reg_module/_01545_ ),
    .X(\reg_module/_01551_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18254_  (.A1(\reg_module/_01544_ ),
    .A2(\reg_module/_07517_ ),
    .B1(\reg_module/_01551_ ),
    .X(\reg_module/_01552_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18255_  (.A(\reg_module/_01550_ ),
    .B(\reg_module/_01552_ ),
    .Y(\reg_module/_00641_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18256_  (.A(net2002),
    .B(\reg_module/_01549_ ),
    .Y(\reg_module/_01553_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18257_  (.A1(\reg_module/_01544_ ),
    .A2(\reg_module/_07520_ ),
    .B1(\reg_module/_01551_ ),
    .X(\reg_module/_01554_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18258_  (.A(\reg_module/_01553_ ),
    .B(\reg_module/_01554_ ),
    .Y(\reg_module/_00642_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_18259_  (.A(\reg_module/_01541_ ),
    .X(\reg_module/_01555_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18260_  (.A1(net1820),
    .A2(\reg_module/_01555_ ),
    .B1(net1047),
    .Y(\reg_module/_01556_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18261_  (.A1(\reg_module/_07523_ ),
    .A2(\reg_module/_01542_ ),
    .B1(\reg_module/_01556_ ),
    .Y(\reg_module/_00643_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18262_  (.A(net1721),
    .B(\reg_module/_01549_ ),
    .Y(\reg_module/_01557_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18263_  (.A1(\reg_module/_01544_ ),
    .A2(\reg_module/_07528_ ),
    .B1(\reg_module/_01551_ ),
    .X(\reg_module/_01558_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18264_  (.A(\reg_module/_01557_ ),
    .B(\reg_module/_01558_ ),
    .Y(\reg_module/_00644_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18265_  (.A(net1953),
    .B(\reg_module/_01549_ ),
    .Y(\reg_module/_01559_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18266_  (.A1(\reg_module/_01544_ ),
    .A2(\reg_module/_07531_ ),
    .B1(\reg_module/_01551_ ),
    .X(\reg_module/_01560_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18267_  (.A(\reg_module/_01559_ ),
    .B(\reg_module/_01560_ ),
    .Y(\reg_module/_00645_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18268_  (.A(net1827),
    .B(\reg_module/_01549_ ),
    .Y(\reg_module/_01561_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18269_  (.A(\reg_module/_01541_ ),
    .X(\reg_module/_01562_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18270_  (.A1(\reg_module/_01562_ ),
    .A2(\reg_module/_07535_ ),
    .B1(\reg_module/_01551_ ),
    .X(\reg_module/_01563_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18271_  (.A(\reg_module/_01561_ ),
    .B(\reg_module/_01563_ ),
    .Y(\reg_module/_00646_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18272_  (.A(net1838),
    .B(\reg_module/_01549_ ),
    .Y(\reg_module/_01564_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18273_  (.A1(\reg_module/_01562_ ),
    .A2(\reg_module/_07538_ ),
    .B1(\reg_module/_01551_ ),
    .X(\reg_module/_01565_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18274_  (.A(\reg_module/_01564_ ),
    .B(\reg_module/_01565_ ),
    .Y(\reg_module/_00647_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18275_  (.A(\reg_module/_01548_ ),
    .X(\reg_module/_01566_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18276_  (.A(net1840),
    .B(\reg_module/_01566_ ),
    .Y(\reg_module/_01567_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18277_  (.A(\reg_module/_01545_ ),
    .X(\reg_module/_01568_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18278_  (.A1(\reg_module/_01562_ ),
    .A2(\reg_module/_07541_ ),
    .B1(\reg_module/_01568_ ),
    .X(\reg_module/_01569_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18279_  (.A(\reg_module/_01567_ ),
    .B(\reg_module/_01569_ ),
    .Y(\reg_module/_00648_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18280_  (.A(net1632),
    .B(\reg_module/_01566_ ),
    .Y(\reg_module/_01570_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18281_  (.A1(\reg_module/_01562_ ),
    .A2(\reg_module/_07544_ ),
    .B1(\reg_module/_01568_ ),
    .X(\reg_module/_01571_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18282_  (.A(\reg_module/_01570_ ),
    .B(\reg_module/_01571_ ),
    .Y(\reg_module/_00649_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18283_  (.A1(net1665),
    .A2(\reg_module/_01555_ ),
    .B1(net1053),
    .Y(\reg_module/_01572_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18284_  (.A1(\reg_module/_07548_ ),
    .A2(\reg_module/_01542_ ),
    .B1(\reg_module/_01572_ ),
    .Y(\reg_module/_00650_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18285_  (.A(net1707),
    .B(\reg_module/_01566_ ),
    .Y(\reg_module/_01573_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18286_  (.A1(\reg_module/_01562_ ),
    .A2(\reg_module/_07551_ ),
    .B1(\reg_module/_01568_ ),
    .X(\reg_module/_01574_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18287_  (.A(\reg_module/_01573_ ),
    .B(\reg_module/_01574_ ),
    .Y(\reg_module/_00651_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18288_  (.A(net1892),
    .B(\reg_module/_01566_ ),
    .Y(\reg_module/_01575_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18289_  (.A1(\reg_module/_01562_ ),
    .A2(\reg_module/_07555_ ),
    .B1(\reg_module/_01568_ ),
    .X(\reg_module/_01576_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18290_  (.A(\reg_module/_01575_ ),
    .B(\reg_module/_01576_ ),
    .Y(\reg_module/_00652_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18291_  (.A1(net1856),
    .A2(\reg_module/_01555_ ),
    .B1(net1053),
    .Y(\reg_module/_01577_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18292_  (.A1(\reg_module/_07558_ ),
    .A2(\reg_module/_01542_ ),
    .B1(\reg_module/_01577_ ),
    .Y(\reg_module/_00653_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18293_  (.A(net1689),
    .B(\reg_module/_01566_ ),
    .Y(\reg_module/_01578_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18294_  (.A(\reg_module/_01541_ ),
    .X(\reg_module/_01579_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18295_  (.A1(\reg_module/_01579_ ),
    .A2(\reg_module/_07561_ ),
    .B1(\reg_module/_01568_ ),
    .X(\reg_module/_01580_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18296_  (.A(\reg_module/_01578_ ),
    .B(\reg_module/_01580_ ),
    .Y(\reg_module/_00654_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18297_  (.A(net1880),
    .B(\reg_module/_01566_ ),
    .Y(\reg_module/_01581_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18298_  (.A1(\reg_module/_01579_ ),
    .A2(\reg_module/_07564_ ),
    .B1(\reg_module/_01568_ ),
    .X(\reg_module/_01582_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18299_  (.A(\reg_module/_01581_ ),
    .B(\reg_module/_01582_ ),
    .Y(\reg_module/_00655_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18300_  (.A(\reg_module/_01541_ ),
    .X(\reg_module/_01583_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18301_  (.A(net1967),
    .B(\reg_module/_01583_ ),
    .Y(\reg_module/_01584_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18302_  (.A(\reg_module/_01545_ ),
    .X(\reg_module/_01585_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18303_  (.A1(\reg_module/_01579_ ),
    .A2(\reg_module/_07568_ ),
    .B1(\reg_module/_01585_ ),
    .X(\reg_module/_01586_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18304_  (.A(\reg_module/_01584_ ),
    .B(\reg_module/_01586_ ),
    .Y(\reg_module/_00656_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18305_  (.A(net1845),
    .B(\reg_module/_01583_ ),
    .Y(\reg_module/_01587_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18306_  (.A1(\reg_module/_01579_ ),
    .A2(\reg_module/_07571_ ),
    .B1(\reg_module/_01585_ ),
    .X(\reg_module/_01588_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18307_  (.A(\reg_module/_01587_ ),
    .B(\reg_module/_01588_ ),
    .Y(\reg_module/_00657_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18308_  (.A1(net1879),
    .A2(\reg_module/_01555_ ),
    .B1(net1044),
    .Y(\reg_module/_01589_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18309_  (.A1(\reg_module/_07575_ ),
    .A2(\reg_module/_01542_ ),
    .B1(\reg_module/_01589_ ),
    .Y(\reg_module/_00658_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18310_  (.A(net1777),
    .B(\reg_module/_01583_ ),
    .Y(\reg_module/_01590_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18311_  (.A1(\reg_module/_01579_ ),
    .A2(\reg_module/_07578_ ),
    .B1(\reg_module/_01585_ ),
    .X(\reg_module/_01591_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18312_  (.A(\reg_module/_01590_ ),
    .B(\reg_module/_01591_ ),
    .Y(\reg_module/_00659_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18313_  (.A(net1718),
    .B(\reg_module/_01583_ ),
    .Y(\reg_module/_01592_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18314_  (.A1(\reg_module/_01579_ ),
    .A2(\reg_module/_07581_ ),
    .B1(\reg_module/_01585_ ),
    .X(\reg_module/_01593_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18315_  (.A(\reg_module/_01592_ ),
    .B(\reg_module/_01593_ ),
    .Y(\reg_module/_00660_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18316_  (.A(net1794),
    .B(\reg_module/_01583_ ),
    .Y(\reg_module/_01594_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18317_  (.A(\reg_module/_01540_ ),
    .X(\reg_module/_01595_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18318_  (.A1(\reg_module/_01595_ ),
    .A2(\reg_module/_07584_ ),
    .B1(\reg_module/_01585_ ),
    .X(\reg_module/_01596_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18319_  (.A(\reg_module/_01594_ ),
    .B(\reg_module/_01596_ ),
    .Y(\reg_module/_00661_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18320_  (.A(net1788),
    .B(\reg_module/_01583_ ),
    .Y(\reg_module/_01597_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18321_  (.A1(\reg_module/_01595_ ),
    .A2(\reg_module/_07588_ ),
    .B1(\reg_module/_01585_ ),
    .X(\reg_module/_01598_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18322_  (.A(\reg_module/_01597_ ),
    .B(\reg_module/_01598_ ),
    .Y(\reg_module/_00662_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18323_  (.A1(\reg_module/gprf[663] ),
    .A2(\reg_module/_01544_ ),
    .B1(net1038),
    .Y(\reg_module/_01599_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18324_  (.A1(\reg_module/_07591_ ),
    .A2(\reg_module/_01542_ ),
    .B1(\reg_module/_01599_ ),
    .Y(\reg_module/_00663_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18325_  (.A(\reg_module/_01541_ ),
    .X(\reg_module/_01600_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18326_  (.A(net1767),
    .B(\reg_module/_01600_ ),
    .Y(\reg_module/_01601_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18327_  (.A(\reg_module/_01545_ ),
    .X(\reg_module/_01602_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18328_  (.A1(\reg_module/_01595_ ),
    .A2(\reg_module/_07595_ ),
    .B1(\reg_module/_01602_ ),
    .X(\reg_module/_01603_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18329_  (.A(\reg_module/_01601_ ),
    .B(\reg_module/_01603_ ),
    .Y(\reg_module/_00664_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18330_  (.A(net1869),
    .B(\reg_module/_01600_ ),
    .Y(\reg_module/_01604_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18331_  (.A1(\reg_module/_01595_ ),
    .A2(\reg_module/_07598_ ),
    .B1(\reg_module/_01602_ ),
    .X(\reg_module/_01605_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18332_  (.A(\reg_module/_01604_ ),
    .B(\reg_module/_01605_ ),
    .Y(\reg_module/_00665_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18333_  (.A(net1678),
    .B(\reg_module/_01600_ ),
    .Y(\reg_module/_01606_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18334_  (.A1(\reg_module/_01595_ ),
    .A2(\reg_module/_07601_ ),
    .B1(\reg_module/_01602_ ),
    .X(\reg_module/_01607_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18335_  (.A(\reg_module/_01606_ ),
    .B(\reg_module/_01607_ ),
    .Y(\reg_module/_00666_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18336_  (.A(net1717),
    .B(\reg_module/_01600_ ),
    .Y(\reg_module/_01608_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18337_  (.A1(\reg_module/_01595_ ),
    .A2(\reg_module/_07604_ ),
    .B1(\reg_module/_01602_ ),
    .X(\reg_module/_01609_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18338_  (.A(\reg_module/_01608_ ),
    .B(\reg_module/_01609_ ),
    .Y(\reg_module/_00667_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18339_  (.A(net1728),
    .B(\reg_module/_01600_ ),
    .Y(\reg_module/_01610_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18340_  (.A1(\reg_module/_01548_ ),
    .A2(\reg_module/_07607_ ),
    .B1(\reg_module/_01602_ ),
    .X(\reg_module/_01611_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18341_  (.A(\reg_module/_01610_ ),
    .B(\reg_module/_01611_ ),
    .Y(\reg_module/_00668_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18342_  (.A(net1804),
    .B(\reg_module/_01600_ ),
    .Y(\reg_module/_01612_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18343_  (.A1(\reg_module/_01548_ ),
    .A2(\reg_module/_07610_ ),
    .B1(\reg_module/_01602_ ),
    .X(\reg_module/_01613_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18344_  (.A(\reg_module/_01612_ ),
    .B(\reg_module/_01613_ ),
    .Y(\reg_module/_00669_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18345_  (.A(net1647),
    .B(\reg_module/_01555_ ),
    .Y(\reg_module/_01614_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18346_  (.A1(\reg_module/_01548_ ),
    .A2(\reg_module/_07613_ ),
    .B1(\reg_module/_07655_ ),
    .X(\reg_module/_01615_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18347_  (.A(\reg_module/_01614_ ),
    .B(\reg_module/_01615_ ),
    .Y(\reg_module/_00670_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18348_  (.A(net1883),
    .B(\reg_module/_01555_ ),
    .Y(\reg_module/_01616_ ));
 sky130_fd_sc_hd__a21o_1 \reg_module/_18349_  (.A1(\reg_module/_01548_ ),
    .A2(\reg_module/_07616_ ),
    .B1(\reg_module/_07655_ ),
    .X(\reg_module/_01617_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18350_  (.A(\reg_module/_01616_ ),
    .B(\reg_module/_01617_ ),
    .Y(\reg_module/_00671_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18351_  (.A(\reg_module/_01281_ ),
    .B(\reg_module/_08359_ ),
    .Y(\reg_module/_01618_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18352_  (.A(\reg_module/_01618_ ),
    .X(\reg_module/_01619_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18353_  (.A(\reg_module/_01619_ ),
    .X(\reg_module/_01620_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18354_  (.A(\reg_module/_01620_ ),
    .B(net1235),
    .Y(\reg_module/_01621_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18355_  (.A(\reg_module/_08370_ ),
    .B(\reg_module/_01527_ ),
    .Y(\reg_module/_01622_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18356_  (.A1(\reg_module/_01621_ ),
    .A2(\reg_module/_01622_ ),
    .B1(\reg_module/_01537_ ),
    .Y(\reg_module/_00672_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18357_  (.A(\reg_module/_01620_ ),
    .B(net1248),
    .Y(\reg_module/_01623_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18358_  (.A(\reg_module/_01458_ ),
    .X(\reg_module/_01624_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18359_  (.A(\reg_module/_08376_ ),
    .B(\reg_module/_01624_ ),
    .Y(\reg_module/_01625_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18360_  (.A1(\reg_module/_01623_ ),
    .A2(\reg_module/_01625_ ),
    .B1(\reg_module/_01537_ ),
    .Y(\reg_module/_00673_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18361_  (.A(\reg_module/_01620_ ),
    .B(net1484),
    .Y(\reg_module/_01626_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18362_  (.A(\reg_module/_08380_ ),
    .B(\reg_module/_01624_ ),
    .Y(\reg_module/_01627_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18363_  (.A1(\reg_module/_01626_ ),
    .A2(\reg_module/_01627_ ),
    .B1(\reg_module/_01537_ ),
    .Y(\reg_module/_00674_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18364_  (.A(\reg_module/_01620_ ),
    .B(net1734),
    .Y(\reg_module/_01628_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18365_  (.A(\reg_module/_08384_ ),
    .B(\reg_module/_01624_ ),
    .Y(\reg_module/_01629_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18366_  (.A1(\reg_module/_01628_ ),
    .A2(\reg_module/_01629_ ),
    .B1(\reg_module/_01537_ ),
    .Y(\reg_module/_00675_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18367_  (.A(\reg_module/_01620_ ),
    .B(net1298),
    .Y(\reg_module/_01630_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18368_  (.A(\reg_module/_08389_ ),
    .B(\reg_module/_01624_ ),
    .Y(\reg_module/_01631_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18369_  (.A(\reg_module/_01507_ ),
    .X(\reg_module/_01632_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18370_  (.A1(\reg_module/_01630_ ),
    .A2(\reg_module/_01631_ ),
    .B1(\reg_module/_01632_ ),
    .Y(\reg_module/_00676_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18371_  (.A(\reg_module/_01620_ ),
    .B(net1338),
    .Y(\reg_module/_01633_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18372_  (.A(\reg_module/_08393_ ),
    .B(\reg_module/_01624_ ),
    .Y(\reg_module/_01634_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18373_  (.A1(\reg_module/_01633_ ),
    .A2(\reg_module/_01634_ ),
    .B1(\reg_module/_01632_ ),
    .Y(\reg_module/_00677_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18374_  (.A(\reg_module/_01619_ ),
    .X(\reg_module/_01635_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18375_  (.A(\reg_module/_01635_ ),
    .B(net1579),
    .Y(\reg_module/_01636_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18376_  (.A(\reg_module/_08400_ ),
    .B(\reg_module/_01624_ ),
    .Y(\reg_module/_01637_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18377_  (.A1(\reg_module/_01636_ ),
    .A2(\reg_module/_01637_ ),
    .B1(\reg_module/_01632_ ),
    .Y(\reg_module/_00678_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18378_  (.A(\reg_module/_01635_ ),
    .B(net1582),
    .Y(\reg_module/_01638_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18379_  (.A(\reg_module/_01287_ ),
    .X(\reg_module/_01639_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18380_  (.A(\reg_module/_08405_ ),
    .B(\reg_module/_01639_ ),
    .Y(\reg_module/_01640_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18381_  (.A1(\reg_module/_01638_ ),
    .A2(\reg_module/_01640_ ),
    .B1(\reg_module/_01632_ ),
    .Y(\reg_module/_00679_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18382_  (.A(\reg_module/_01635_ ),
    .B(net1922),
    .Y(\reg_module/_01641_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18383_  (.A(\reg_module/_08409_ ),
    .B(\reg_module/_01639_ ),
    .Y(\reg_module/_01642_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18384_  (.A1(\reg_module/_01641_ ),
    .A2(\reg_module/_01642_ ),
    .B1(\reg_module/_01632_ ),
    .Y(\reg_module/_00680_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18385_  (.A(\reg_module/_01635_ ),
    .B(net2034),
    .Y(\reg_module/_01643_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18386_  (.A(\reg_module/_08413_ ),
    .B(\reg_module/_01639_ ),
    .Y(\reg_module/_01644_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18387_  (.A1(\reg_module/_01643_ ),
    .A2(\reg_module/_01644_ ),
    .B1(\reg_module/_01632_ ),
    .Y(\reg_module/_00681_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18388_  (.A(\reg_module/_01635_ ),
    .B(net1934),
    .Y(\reg_module/_01645_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18389_  (.A(\reg_module/_08418_ ),
    .B(\reg_module/_01639_ ),
    .Y(\reg_module/_01646_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18390_  (.A(\reg_module/_01507_ ),
    .X(\reg_module/_01647_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18391_  (.A1(\reg_module/_01645_ ),
    .A2(\reg_module/_01646_ ),
    .B1(\reg_module/_01647_ ),
    .Y(\reg_module/_00682_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18392_  (.A(\reg_module/_01635_ ),
    .B(net1714),
    .Y(\reg_module/_01648_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18393_  (.A(\reg_module/_08422_ ),
    .B(\reg_module/_01639_ ),
    .Y(\reg_module/_01649_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18394_  (.A1(\reg_module/_01648_ ),
    .A2(\reg_module/_01649_ ),
    .B1(\reg_module/_01647_ ),
    .Y(\reg_module/_00683_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18395_  (.A(\reg_module/_01619_ ),
    .X(\reg_module/_01650_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18396_  (.A(\reg_module/_01650_ ),
    .B(net1854),
    .Y(\reg_module/_01651_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18397_  (.A(\reg_module/_08429_ ),
    .B(\reg_module/_01639_ ),
    .Y(\reg_module/_01652_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18398_  (.A1(\reg_module/_01651_ ),
    .A2(\reg_module/_01652_ ),
    .B1(\reg_module/_01647_ ),
    .Y(\reg_module/_00684_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18399_  (.A(\reg_module/_01650_ ),
    .B(net1924),
    .Y(\reg_module/_01653_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18400_  (.A(\reg_module/_01287_ ),
    .X(\reg_module/_01654_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18401_  (.A(\reg_module/_08434_ ),
    .B(\reg_module/_01654_ ),
    .Y(\reg_module/_01655_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18402_  (.A1(\reg_module/_01653_ ),
    .A2(\reg_module/_01655_ ),
    .B1(\reg_module/_01647_ ),
    .Y(\reg_module/_00685_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18403_  (.A(\reg_module/_01650_ ),
    .B(net1268),
    .Y(\reg_module/_01656_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18404_  (.A(\reg_module/_08438_ ),
    .B(\reg_module/_01654_ ),
    .Y(\reg_module/_01657_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18405_  (.A1(\reg_module/_01656_ ),
    .A2(\reg_module/_01657_ ),
    .B1(\reg_module/_01647_ ),
    .Y(\reg_module/_00686_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18406_  (.A(\reg_module/_01650_ ),
    .B(net1832),
    .Y(\reg_module/_01658_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18407_  (.A(\reg_module/_08442_ ),
    .B(\reg_module/_01654_ ),
    .Y(\reg_module/_01659_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18408_  (.A1(\reg_module/_01658_ ),
    .A2(\reg_module/_01659_ ),
    .B1(\reg_module/_01647_ ),
    .Y(\reg_module/_00687_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18409_  (.A(\reg_module/_01650_ ),
    .B(net1519),
    .Y(\reg_module/_01660_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18410_  (.A(\reg_module/_08447_ ),
    .B(\reg_module/_01654_ ),
    .Y(\reg_module/_01661_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18411_  (.A(\reg_module/_01507_ ),
    .X(\reg_module/_01662_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18412_  (.A1(\reg_module/_01660_ ),
    .A2(\reg_module/_01661_ ),
    .B1(\reg_module/_01662_ ),
    .Y(\reg_module/_00688_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18413_  (.A(\reg_module/_01650_ ),
    .B(net1258),
    .Y(\reg_module/_01663_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18414_  (.A(\reg_module/_08451_ ),
    .B(\reg_module/_01654_ ),
    .Y(\reg_module/_01664_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18415_  (.A1(\reg_module/_01663_ ),
    .A2(\reg_module/_01664_ ),
    .B1(\reg_module/_01662_ ),
    .Y(\reg_module/_00689_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18416_  (.A(\reg_module/_01619_ ),
    .X(\reg_module/_01665_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18417_  (.A(\reg_module/_01665_ ),
    .B(net1474),
    .Y(\reg_module/_01666_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18418_  (.A(\reg_module/_08458_ ),
    .B(\reg_module/_01654_ ),
    .Y(\reg_module/_01667_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18419_  (.A1(\reg_module/_01666_ ),
    .A2(\reg_module/_01667_ ),
    .B1(\reg_module/_01662_ ),
    .Y(\reg_module/_00690_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18420_  (.A(\reg_module/_01665_ ),
    .B(net1280),
    .Y(\reg_module/_01668_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18421_  (.A(\reg_module/_01287_ ),
    .X(\reg_module/_01669_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18422_  (.A(\reg_module/_08463_ ),
    .B(\reg_module/_01669_ ),
    .Y(\reg_module/_01670_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18423_  (.A1(\reg_module/_01668_ ),
    .A2(\reg_module/_01670_ ),
    .B1(\reg_module/_01662_ ),
    .Y(\reg_module/_00691_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18424_  (.A(\reg_module/_01665_ ),
    .B(net1294),
    .Y(\reg_module/_01671_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18425_  (.A(\reg_module/_08467_ ),
    .B(\reg_module/_01669_ ),
    .Y(\reg_module/_01672_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18426_  (.A1(\reg_module/_01671_ ),
    .A2(\reg_module/_01672_ ),
    .B1(\reg_module/_01662_ ),
    .Y(\reg_module/_00692_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18427_  (.A(\reg_module/_01665_ ),
    .B(net1253),
    .Y(\reg_module/_01673_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18428_  (.A(\reg_module/_08471_ ),
    .B(\reg_module/_01669_ ),
    .Y(\reg_module/_01674_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18429_  (.A1(\reg_module/_01673_ ),
    .A2(\reg_module/_01674_ ),
    .B1(\reg_module/_01662_ ),
    .Y(\reg_module/_00693_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18430_  (.A(\reg_module/_01665_ ),
    .B(net1233),
    .Y(\reg_module/_01675_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18431_  (.A(\reg_module/_08476_ ),
    .B(\reg_module/_01669_ ),
    .Y(\reg_module/_01676_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18432_  (.A(\reg_module/_01506_ ),
    .X(\reg_module/_01677_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18433_  (.A(\reg_module/_01677_ ),
    .X(\reg_module/_01678_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18434_  (.A1(\reg_module/_01675_ ),
    .A2(\reg_module/_01676_ ),
    .B1(\reg_module/_01678_ ),
    .Y(\reg_module/_00694_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18435_  (.A(\reg_module/_01665_ ),
    .B(net1242),
    .Y(\reg_module/_01679_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18436_  (.A(\reg_module/_08480_ ),
    .B(\reg_module/_01669_ ),
    .Y(\reg_module/_01680_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18437_  (.A1(\reg_module/_01679_ ),
    .A2(\reg_module/_01680_ ),
    .B1(\reg_module/_01678_ ),
    .Y(\reg_module/_00695_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18438_  (.A(\reg_module/_01618_ ),
    .X(\reg_module/_01681_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18439_  (.A(\reg_module/_01681_ ),
    .B(net1478),
    .Y(\reg_module/_01682_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18440_  (.A(\reg_module/_08487_ ),
    .B(\reg_module/_01669_ ),
    .Y(\reg_module/_01683_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18441_  (.A1(\reg_module/_01682_ ),
    .A2(\reg_module/_01683_ ),
    .B1(\reg_module/_01678_ ),
    .Y(\reg_module/_00696_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18442_  (.A(\reg_module/_01681_ ),
    .B(net1289),
    .Y(\reg_module/_01684_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18443_  (.A(\reg_module/_01287_ ),
    .X(\reg_module/_01685_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18444_  (.A(\reg_module/_08492_ ),
    .B(\reg_module/_01685_ ),
    .Y(\reg_module/_01686_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18445_  (.A1(\reg_module/_01684_ ),
    .A2(\reg_module/_01686_ ),
    .B1(\reg_module/_01678_ ),
    .Y(\reg_module/_00697_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18446_  (.A(\reg_module/_01681_ ),
    .B(net1287),
    .Y(\reg_module/_01687_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18447_  (.A(\reg_module/_08496_ ),
    .B(\reg_module/_01685_ ),
    .Y(\reg_module/_01688_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18448_  (.A1(\reg_module/_01687_ ),
    .A2(\reg_module/_01688_ ),
    .B1(\reg_module/_01678_ ),
    .Y(\reg_module/_00698_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18449_  (.A(\reg_module/_01681_ ),
    .B(net1764),
    .Y(\reg_module/_01689_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18450_  (.A(\reg_module/_08500_ ),
    .B(\reg_module/_01685_ ),
    .Y(\reg_module/_01690_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18451_  (.A1(\reg_module/_01689_ ),
    .A2(\reg_module/_01690_ ),
    .B1(\reg_module/_01678_ ),
    .Y(\reg_module/_00699_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18452_  (.A(\reg_module/_01681_ ),
    .B(net1897),
    .Y(\reg_module/_01691_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18453_  (.A(\reg_module/_08505_ ),
    .B(\reg_module/_01685_ ),
    .Y(\reg_module/_01692_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18454_  (.A(\reg_module/_01677_ ),
    .X(\reg_module/_01693_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18455_  (.A1(\reg_module/_01691_ ),
    .A2(\reg_module/_01692_ ),
    .B1(\reg_module/_01693_ ),
    .Y(\reg_module/_00700_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18456_  (.A(\reg_module/_01681_ ),
    .B(net1561),
    .Y(\reg_module/_01694_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18457_  (.A(\reg_module/_08509_ ),
    .B(\reg_module/_01685_ ),
    .Y(\reg_module/_01695_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18458_  (.A1(\reg_module/_01694_ ),
    .A2(\reg_module/_01695_ ),
    .B1(\reg_module/_01693_ ),
    .Y(\reg_module/_00701_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18459_  (.A(\reg_module/_01619_ ),
    .B(net1585),
    .Y(\reg_module/_01696_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18460_  (.A(\reg_module/_08514_ ),
    .B(\reg_module/_01685_ ),
    .Y(\reg_module/_01697_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18461_  (.A1(\reg_module/_01696_ ),
    .A2(\reg_module/_01697_ ),
    .B1(\reg_module/_01693_ ),
    .Y(\reg_module/_00702_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18462_  (.A(\reg_module/_01619_ ),
    .B(net1469),
    .Y(\reg_module/_01698_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_18463_  (.A(\reg_module/_01287_ ),
    .X(\reg_module/_01699_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18464_  (.A(\reg_module/_08519_ ),
    .B(\reg_module/_01699_ ),
    .Y(\reg_module/_01700_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18465_  (.A1(\reg_module/_01698_ ),
    .A2(\reg_module/_01700_ ),
    .B1(\reg_module/_01693_ ),
    .Y(\reg_module/_00703_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18466_  (.A(\reg_module/_01281_ ),
    .B(\reg_module/_08521_ ),
    .Y(\reg_module/_01701_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_18467_  (.A(\reg_module/_01701_ ),
    .X(\reg_module/_01702_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18468_  (.A(\reg_module/_01702_ ),
    .X(\reg_module/_01703_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18469_  (.A(\reg_module/_01703_ ),
    .B(net1395),
    .Y(\reg_module/_01704_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18470_  (.A(\reg_module/_01699_ ),
    .X(\reg_module/_01705_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18471_  (.A(\reg_module/_01705_ ),
    .B(\reg_module/_08528_ ),
    .Y(\reg_module/_01706_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18472_  (.A1(\reg_module/_01704_ ),
    .A2(\reg_module/_01706_ ),
    .B1(\reg_module/_01693_ ),
    .Y(\reg_module/_00704_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18473_  (.A(\reg_module/_01703_ ),
    .B(net1413),
    .Y(\reg_module/_01707_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18474_  (.A(\reg_module/_01705_ ),
    .B(\reg_module/_08531_ ),
    .Y(\reg_module/_01708_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18475_  (.A1(\reg_module/_01707_ ),
    .A2(\reg_module/_01708_ ),
    .B1(\reg_module/_01693_ ),
    .Y(\reg_module/_00705_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18476_  (.A(\reg_module/_01703_ ),
    .B(net1369),
    .Y(\reg_module/_01709_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18477_  (.A(\reg_module/_01705_ ),
    .B(net285),
    .Y(\reg_module/_01710_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18478_  (.A(\reg_module/_01677_ ),
    .X(\reg_module/_01711_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18479_  (.A1(\reg_module/_01709_ ),
    .A2(\reg_module/_01710_ ),
    .B1(\reg_module/_01711_ ),
    .Y(\reg_module/_00706_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18480_  (.A(\reg_module/_01703_ ),
    .B(net1381),
    .Y(\reg_module/_01712_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18481_  (.A(\reg_module/_01471_ ),
    .B(\reg_module/_08537_ ),
    .Y(\reg_module/_01713_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18482_  (.A1(\reg_module/_01712_ ),
    .A2(\reg_module/_01713_ ),
    .B1(\reg_module/_01711_ ),
    .Y(\reg_module/_00707_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18483_  (.A(\reg_module/_01703_ ),
    .B(net1246),
    .Y(\reg_module/_01714_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18484_  (.A(\reg_module/_01705_ ),
    .B(net284),
    .Y(\reg_module/_01715_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18485_  (.A1(\reg_module/_01714_ ),
    .A2(\reg_module/_01715_ ),
    .B1(\reg_module/_01711_ ),
    .Y(\reg_module/_00708_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18486_  (.A(\reg_module/_01703_ ),
    .B(net1917),
    .Y(\reg_module/_01716_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18487_  (.A(\reg_module/_01705_ ),
    .B(net283),
    .Y(\reg_module/_01717_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18488_  (.A1(\reg_module/_01716_ ),
    .A2(\reg_module/_01717_ ),
    .B1(\reg_module/_01711_ ),
    .Y(\reg_module/_00709_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18489_  (.A(\reg_module/_01702_ ),
    .X(\reg_module/_01718_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18490_  (.A(\reg_module/_01718_ ),
    .B(net1538),
    .Y(\reg_module/_01719_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18491_  (.A(\reg_module/_01705_ ),
    .B(\reg_module/_08552_ ),
    .Y(\reg_module/_01720_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18492_  (.A1(\reg_module/_01719_ ),
    .A2(\reg_module/_01720_ ),
    .B1(\reg_module/_01711_ ),
    .Y(\reg_module/_00710_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18493_  (.A(\reg_module/_01718_ ),
    .B(net1460),
    .Y(\reg_module/_01721_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18494_  (.A(\reg_module/_01699_ ),
    .X(\reg_module/_01722_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18495_  (.A(\reg_module/_01722_ ),
    .B(\reg_module/_08555_ ),
    .Y(\reg_module/_01723_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18496_  (.A1(\reg_module/_01721_ ),
    .A2(\reg_module/_01723_ ),
    .B1(\reg_module/_01711_ ),
    .Y(\reg_module/_00711_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18497_  (.A(\reg_module/_01718_ ),
    .B(net1886),
    .Y(\reg_module/_01724_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18498_  (.A(\reg_module/_01722_ ),
    .B(\reg_module/_08558_ ),
    .Y(\reg_module/_01725_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18499_  (.A(\reg_module/_01677_ ),
    .X(\reg_module/_01726_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18500_  (.A1(\reg_module/_01724_ ),
    .A2(\reg_module/_01725_ ),
    .B1(\reg_module/_01726_ ),
    .Y(\reg_module/_00712_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18501_  (.A(\reg_module/_01718_ ),
    .B(net1802),
    .Y(\reg_module/_01727_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18502_  (.A(\reg_module/_01722_ ),
    .B(\reg_module/_08561_ ),
    .Y(\reg_module/_01728_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18503_  (.A1(\reg_module/_01727_ ),
    .A2(\reg_module/_01728_ ),
    .B1(\reg_module/_01726_ ),
    .Y(\reg_module/_00713_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18504_  (.A(\reg_module/_01718_ ),
    .B(net1382),
    .Y(\reg_module/_01729_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18505_  (.A(\reg_module/_01471_ ),
    .B(\reg_module/_08565_ ),
    .Y(\reg_module/_01730_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18506_  (.A1(\reg_module/_01729_ ),
    .A2(\reg_module/_01730_ ),
    .B1(\reg_module/_01726_ ),
    .Y(\reg_module/_00714_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18507_  (.A(\reg_module/_01718_ ),
    .B(net2022),
    .Y(\reg_module/_01731_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18508_  (.A(\reg_module/_01722_ ),
    .B(\reg_module/_08569_ ),
    .Y(\reg_module/_01732_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18509_  (.A1(\reg_module/_01731_ ),
    .A2(\reg_module/_01732_ ),
    .B1(\reg_module/_01726_ ),
    .Y(\reg_module/_00715_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18510_  (.A(\reg_module/_01702_ ),
    .X(\reg_module/_01733_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18511_  (.A(\reg_module/_01733_ ),
    .B(net1587),
    .Y(\reg_module/_01734_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18512_  (.A(\reg_module/_01722_ ),
    .B(\reg_module/_08575_ ),
    .Y(\reg_module/_01735_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18513_  (.A1(\reg_module/_01734_ ),
    .A2(\reg_module/_01735_ ),
    .B1(\reg_module/_01726_ ),
    .Y(\reg_module/_00716_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18514_  (.A(\reg_module/_01733_ ),
    .B(net1771),
    .Y(\reg_module/_01736_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18515_  (.A(\reg_module/_01471_ ),
    .B(\reg_module/_08578_ ),
    .Y(\reg_module/_01737_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18516_  (.A1(\reg_module/_01736_ ),
    .A2(\reg_module/_01737_ ),
    .B1(\reg_module/_01726_ ),
    .Y(\reg_module/_00717_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18517_  (.A(\reg_module/_01733_ ),
    .B(net1920),
    .Y(\reg_module/_01738_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18518_  (.A(\reg_module/_01722_ ),
    .B(\reg_module/_08581_ ),
    .Y(\reg_module/_01739_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18519_  (.A(\reg_module/_01677_ ),
    .X(\reg_module/_01740_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18520_  (.A1(\reg_module/_01738_ ),
    .A2(\reg_module/_01739_ ),
    .B1(\reg_module/_01740_ ),
    .Y(\reg_module/_00718_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18521_  (.A(\reg_module/_01733_ ),
    .B(net1667),
    .Y(\reg_module/_01741_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18522_  (.A(\reg_module/_01699_ ),
    .X(\reg_module/_01742_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18523_  (.A(\reg_module/_01742_ ),
    .B(\reg_module/_08584_ ),
    .Y(\reg_module/_01743_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18524_  (.A1(\reg_module/_01741_ ),
    .A2(\reg_module/_01743_ ),
    .B1(\reg_module/_01740_ ),
    .Y(\reg_module/_00719_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18525_  (.A(\reg_module/_01733_ ),
    .B(net1558),
    .Y(\reg_module/_01744_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18526_  (.A(\reg_module/_01742_ ),
    .B(\reg_module/_08588_ ),
    .Y(\reg_module/_01745_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18527_  (.A1(\reg_module/_01744_ ),
    .A2(\reg_module/_01745_ ),
    .B1(\reg_module/_01740_ ),
    .Y(\reg_module/_00720_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18528_  (.A(\reg_module/_01733_ ),
    .B(net1979),
    .Y(\reg_module/_01746_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18529_  (.A(\reg_module/_01742_ ),
    .B(\reg_module/_08592_ ),
    .Y(\reg_module/_01747_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18530_  (.A1(\reg_module/_01746_ ),
    .A2(\reg_module/_01747_ ),
    .B1(\reg_module/_01740_ ),
    .Y(\reg_module/_00721_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18531_  (.A(\reg_module/_01702_ ),
    .X(\reg_module/_01748_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18532_  (.A(\reg_module/_01748_ ),
    .B(net1461),
    .Y(\reg_module/_01749_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18533_  (.A(\reg_module/_01381_ ),
    .X(\reg_module/_01750_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18534_  (.A(\reg_module/_01750_ ),
    .B(\reg_module/_08597_ ),
    .Y(\reg_module/_01751_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18535_  (.A1(\reg_module/_01749_ ),
    .A2(\reg_module/_01751_ ),
    .B1(\reg_module/_01740_ ),
    .Y(\reg_module/_00722_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18536_  (.A(\reg_module/_01748_ ),
    .B(net1453),
    .Y(\reg_module/_01752_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18537_  (.A(\reg_module/_01742_ ),
    .B(\reg_module/_08600_ ),
    .Y(\reg_module/_01753_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18538_  (.A1(\reg_module/_01752_ ),
    .A2(\reg_module/_01753_ ),
    .B1(\reg_module/_01740_ ),
    .Y(\reg_module/_00723_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18539_  (.A(\reg_module/_01748_ ),
    .B(net1432),
    .Y(\reg_module/_01754_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18540_  (.A(\reg_module/_01742_ ),
    .B(net282),
    .Y(\reg_module/_01755_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18541_  (.A(\reg_module/_01677_ ),
    .X(\reg_module/_01756_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18542_  (.A1(\reg_module/_01754_ ),
    .A2(\reg_module/_01755_ ),
    .B1(\reg_module/_01756_ ),
    .Y(\reg_module/_00724_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18543_  (.A(\reg_module/_01748_ ),
    .B(net1301),
    .Y(\reg_module/_01757_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18544_  (.A(\reg_module/_01742_ ),
    .B(net281),
    .Y(\reg_module/_01758_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18545_  (.A1(\reg_module/_01757_ ),
    .A2(\reg_module/_01758_ ),
    .B1(\reg_module/_01756_ ),
    .Y(\reg_module/_00725_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18546_  (.A(\reg_module/_01748_ ),
    .B(net1335),
    .Y(\reg_module/_01759_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18547_  (.A(\reg_module/_01699_ ),
    .X(\reg_module/_01760_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18548_  (.A(\reg_module/_01760_ ),
    .B(\reg_module/_08610_ ),
    .Y(\reg_module/_01761_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18549_  (.A1(\reg_module/_01759_ ),
    .A2(\reg_module/_01761_ ),
    .B1(\reg_module/_01756_ ),
    .Y(\reg_module/_00726_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18550_  (.A(\reg_module/_01748_ ),
    .B(net1389),
    .Y(\reg_module/_01762_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18551_  (.A(\reg_module/_01750_ ),
    .B(\reg_module/_08614_ ),
    .Y(\reg_module/_01763_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18552_  (.A1(\reg_module/_01762_ ),
    .A2(\reg_module/_01763_ ),
    .B1(\reg_module/_01756_ ),
    .Y(\reg_module/_00727_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18553_  (.A(\reg_module/_01701_ ),
    .X(\reg_module/_01764_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18554_  (.A(\reg_module/_01764_ ),
    .B(net1834),
    .Y(\reg_module/_01765_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18555_  (.A(\reg_module/_01760_ ),
    .B(\reg_module/_08619_ ),
    .Y(\reg_module/_01766_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18556_  (.A1(\reg_module/_01765_ ),
    .A2(\reg_module/_01766_ ),
    .B1(\reg_module/_01756_ ),
    .Y(\reg_module/_00728_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18557_  (.A(\reg_module/_01764_ ),
    .B(net1837),
    .Y(\reg_module/_01767_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18558_  (.A(\reg_module/_01760_ ),
    .B(\reg_module/_08622_ ),
    .Y(\reg_module/_01768_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18559_  (.A1(\reg_module/_01767_ ),
    .A2(\reg_module/_01768_ ),
    .B1(\reg_module/_01756_ ),
    .Y(\reg_module/_00729_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18560_  (.A(\reg_module/_01764_ ),
    .B(net1308),
    .Y(\reg_module/_01769_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18561_  (.A(\reg_module/_01760_ ),
    .B(\reg_module/_08625_ ),
    .Y(\reg_module/_01770_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18562_  (.A(\reg_module/_01506_ ),
    .X(\reg_module/_01771_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18563_  (.A(\reg_module/_01771_ ),
    .X(\reg_module/_01772_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18564_  (.A1(\reg_module/_01769_ ),
    .A2(\reg_module/_01770_ ),
    .B1(\reg_module/_01772_ ),
    .Y(\reg_module/_00730_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18565_  (.A(\reg_module/_01764_ ),
    .B(net1921),
    .Y(\reg_module/_01773_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18566_  (.A(\reg_module/_01760_ ),
    .B(\reg_module/_08628_ ),
    .Y(\reg_module/_01774_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18567_  (.A1(\reg_module/_01773_ ),
    .A2(\reg_module/_01774_ ),
    .B1(\reg_module/_01772_ ),
    .Y(\reg_module/_00731_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18568_  (.A(\reg_module/_01764_ ),
    .B(net1978),
    .Y(\reg_module/_01775_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18569_  (.A(\reg_module/_01760_ ),
    .B(\reg_module/_08632_ ),
    .Y(\reg_module/_01776_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18570_  (.A1(\reg_module/_01775_ ),
    .A2(\reg_module/_01776_ ),
    .B1(\reg_module/_01772_ ),
    .Y(\reg_module/_00732_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18571_  (.A(\reg_module/_01764_ ),
    .B(net1634),
    .Y(\reg_module/_01777_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18572_  (.A(\reg_module/_01699_ ),
    .X(\reg_module/_01778_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18573_  (.A(\reg_module/_01778_ ),
    .B(\reg_module/_08636_ ),
    .Y(\reg_module/_01779_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18574_  (.A1(\reg_module/_01777_ ),
    .A2(\reg_module/_01779_ ),
    .B1(\reg_module/_01772_ ),
    .Y(\reg_module/_00733_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18575_  (.A(\reg_module/_01702_ ),
    .B(net1705),
    .Y(\reg_module/_01780_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18576_  (.A(\reg_module/_01778_ ),
    .B(\reg_module/_08640_ ),
    .Y(\reg_module/_01781_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18577_  (.A1(\reg_module/_01780_ ),
    .A2(\reg_module/_01781_ ),
    .B1(\reg_module/_01772_ ),
    .Y(\reg_module/_00734_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18578_  (.A(\reg_module/_01702_ ),
    .B(net1968),
    .Y(\reg_module/_01782_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18579_  (.A(\reg_module/_01778_ ),
    .B(\reg_module/_08643_ ),
    .Y(\reg_module/_01783_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18580_  (.A1(\reg_module/_01782_ ),
    .A2(\reg_module/_01783_ ),
    .B1(\reg_module/_01772_ ),
    .Y(\reg_module/_00735_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_18581_  (.A(\reg_module/_08646_ ),
    .B(\reg_module/_01154_ ),
    .Y(\reg_module/_01784_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_18582_  (.A(\reg_module/_01784_ ),
    .Y(\reg_module/_01785_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18583_  (.A(\reg_module/_01785_ ),
    .X(\reg_module/_01786_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18584_  (.A(\reg_module/_01786_ ),
    .B(net1757),
    .Y(\reg_module/_01787_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18585_  (.A(\reg_module/_01784_ ),
    .X(\reg_module/_01788_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18586_  (.A(\reg_module/_01788_ ),
    .X(\reg_module/_01789_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18587_  (.A(\reg_module/_01789_ ),
    .B(net318),
    .Y(\reg_module/_01790_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18588_  (.A(\reg_module/_01771_ ),
    .X(\reg_module/_01791_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18589_  (.A1(\reg_module/_01787_ ),
    .A2(\reg_module/_01790_ ),
    .B1(\reg_module/_01791_ ),
    .Y(\reg_module/_00736_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18590_  (.A(\reg_module/_01786_ ),
    .B(net1418),
    .Y(\reg_module/_01792_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18591_  (.A(\reg_module/_01789_ ),
    .B(net317),
    .Y(\reg_module/_01793_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18592_  (.A1(\reg_module/_01792_ ),
    .A2(\reg_module/_01793_ ),
    .B1(\reg_module/_01791_ ),
    .Y(\reg_module/_00737_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18593_  (.A(\reg_module/_01786_ ),
    .B(net1499),
    .Y(\reg_module/_01794_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18594_  (.A(\reg_module/_01788_ ),
    .X(\reg_module/_01795_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18595_  (.A(\reg_module/_01795_ ),
    .B(net316),
    .Y(\reg_module/_01796_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18596_  (.A1(\reg_module/_01794_ ),
    .A2(\reg_module/_01796_ ),
    .B1(\reg_module/_01791_ ),
    .Y(\reg_module/_00738_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18597_  (.A(\reg_module/_01786_ ),
    .B(net1311),
    .Y(\reg_module/_01797_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18598_  (.A(\reg_module/_01795_ ),
    .B(net315),
    .Y(\reg_module/_01798_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18599_  (.A1(\reg_module/_01797_ ),
    .A2(\reg_module/_01798_ ),
    .B1(\reg_module/_01791_ ),
    .Y(\reg_module/_00739_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18600_  (.A(\reg_module/_01788_ ),
    .X(\reg_module/_01799_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18601_  (.A(\reg_module/_01788_ ),
    .X(\reg_module/_01800_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18602_  (.A1(net1899),
    .A2(\reg_module/_01800_ ),
    .B1(net1037),
    .Y(\reg_module/_01801_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18603_  (.A1(\reg_module/_07528_ ),
    .A2(\reg_module/_01799_ ),
    .B1(\reg_module/_01801_ ),
    .Y(\reg_module/_00740_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18604_  (.A(\reg_module/_01786_ ),
    .B(net1379),
    .Y(\reg_module/_01802_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18605_  (.A(\reg_module/_01795_ ),
    .B(net314),
    .Y(\reg_module/_01803_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18606_  (.A1(\reg_module/_01802_ ),
    .A2(\reg_module/_01803_ ),
    .B1(\reg_module/_01791_ ),
    .Y(\reg_module/_00741_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18607_  (.A(\reg_module/_01788_ ),
    .X(\reg_module/_01804_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18608_  (.A1(net1567),
    .A2(\reg_module/_01804_ ),
    .B1(net1047),
    .Y(\reg_module/_01805_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18609_  (.A1(\reg_module/_07535_ ),
    .A2(\reg_module/_01799_ ),
    .B1(\reg_module/_01805_ ),
    .Y(\reg_module/_00742_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18610_  (.A(\reg_module/_01786_ ),
    .B(net1580),
    .Y(\reg_module/_01806_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18611_  (.A(\reg_module/_01795_ ),
    .B(net313),
    .Y(\reg_module/_01807_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18612_  (.A1(\reg_module/_01806_ ),
    .A2(\reg_module/_01807_ ),
    .B1(\reg_module/_01791_ ),
    .Y(\reg_module/_00743_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18613_  (.A1(net1709),
    .A2(\reg_module/_01804_ ),
    .B1(net1043),
    .Y(\reg_module/_01808_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18614_  (.A1(\reg_module/_07541_ ),
    .A2(\reg_module/_01799_ ),
    .B1(\reg_module/_01808_ ),
    .Y(\reg_module/_00744_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18615_  (.A(\reg_module/_01785_ ),
    .X(\reg_module/_01809_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18616_  (.A(\reg_module/_01809_ ),
    .B(net1237),
    .Y(\reg_module/_01810_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18617_  (.A(\reg_module/_01795_ ),
    .B(net312),
    .Y(\reg_module/_01811_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18618_  (.A(\reg_module/_01771_ ),
    .X(\reg_module/_01812_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18619_  (.A1(\reg_module/_01810_ ),
    .A2(\reg_module/_01811_ ),
    .B1(\reg_module/_01812_ ),
    .Y(\reg_module/_00745_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18620_  (.A(\reg_module/_01809_ ),
    .B(net1403),
    .Y(\reg_module/_01813_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18621_  (.A(\reg_module/_01795_ ),
    .B(net311),
    .Y(\reg_module/_01814_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18622_  (.A1(\reg_module/_01813_ ),
    .A2(\reg_module/_01814_ ),
    .B1(\reg_module/_01812_ ),
    .Y(\reg_module/_00746_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18623_  (.A(\reg_module/_01809_ ),
    .B(net1244),
    .Y(\reg_module/_01815_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18624_  (.A(\reg_module/_01784_ ),
    .X(\reg_module/_01816_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18625_  (.A(\reg_module/_01816_ ),
    .B(net310),
    .Y(\reg_module/_01817_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18626_  (.A1(\reg_module/_01815_ ),
    .A2(\reg_module/_01817_ ),
    .B1(\reg_module/_01812_ ),
    .Y(\reg_module/_00747_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18627_  (.A1(net1801),
    .A2(\reg_module/_01804_ ),
    .B1(net1053),
    .Y(\reg_module/_01818_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18628_  (.A1(\reg_module/_07555_ ),
    .A2(\reg_module/_01799_ ),
    .B1(\reg_module/_01818_ ),
    .Y(\reg_module/_00748_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18629_  (.A(\reg_module/_01809_ ),
    .B(net1622),
    .Y(\reg_module/_01819_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18630_  (.A(\reg_module/_01816_ ),
    .B(net309),
    .Y(\reg_module/_01820_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18631_  (.A1(\reg_module/_01819_ ),
    .A2(\reg_module/_01820_ ),
    .B1(\reg_module/_01812_ ),
    .Y(\reg_module/_00749_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18632_  (.A1(net1716),
    .A2(\reg_module/_01804_ ),
    .B1(net1044),
    .Y(\reg_module/_01821_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18633_  (.A1(\reg_module/_07561_ ),
    .A2(\reg_module/_01799_ ),
    .B1(\reg_module/_01821_ ),
    .Y(\reg_module/_00750_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18634_  (.A(\reg_module/_01809_ ),
    .B(net1334),
    .Y(\reg_module/_01822_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18635_  (.A(\reg_module/_01816_ ),
    .B(net306),
    .Y(\reg_module/_01823_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18636_  (.A1(\reg_module/_01822_ ),
    .A2(\reg_module/_01823_ ),
    .B1(\reg_module/_01812_ ),
    .Y(\reg_module/_00751_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18637_  (.A1(net1660),
    .A2(\reg_module/_01804_ ),
    .B1(net1053),
    .Y(\reg_module/_01824_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18638_  (.A1(\reg_module/_07568_ ),
    .A2(\reg_module/_01799_ ),
    .B1(\reg_module/_01824_ ),
    .Y(\reg_module/_00752_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18639_  (.A(\reg_module/_01809_ ),
    .B(net1270),
    .Y(\reg_module/_01825_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18640_  (.A(\reg_module/_01816_ ),
    .B(net305),
    .Y(\reg_module/_01826_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18641_  (.A1(\reg_module/_01825_ ),
    .A2(\reg_module/_01826_ ),
    .B1(\reg_module/_01812_ ),
    .Y(\reg_module/_00753_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18642_  (.A(\reg_module/_01785_ ),
    .X(\reg_module/_01827_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18643_  (.A(\reg_module/_01827_ ),
    .B(net1759),
    .Y(\reg_module/_01828_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18644_  (.A(\reg_module/_01816_ ),
    .B(net304),
    .Y(\reg_module/_01829_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18645_  (.A(\reg_module/_01771_ ),
    .X(\reg_module/_01830_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18646_  (.A1(\reg_module/_01828_ ),
    .A2(\reg_module/_01829_ ),
    .B1(\reg_module/_01830_ ),
    .Y(\reg_module/_00754_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18647_  (.A(\reg_module/_01827_ ),
    .B(net1316),
    .Y(\reg_module/_01831_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18648_  (.A(\reg_module/_01816_ ),
    .B(net303),
    .Y(\reg_module/_01832_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18649_  (.A1(\reg_module/_01831_ ),
    .A2(\reg_module/_01832_ ),
    .B1(\reg_module/_01830_ ),
    .Y(\reg_module/_00755_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18650_  (.A1(net1988),
    .A2(\reg_module/_01804_ ),
    .B1(net1041),
    .Y(\reg_module/_01833_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18651_  (.A1(\reg_module/_07581_ ),
    .A2(\reg_module/_01800_ ),
    .B1(\reg_module/_01833_ ),
    .Y(\reg_module/_00756_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18652_  (.A(\reg_module/_01827_ ),
    .B(net1719),
    .Y(\reg_module/_01834_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18653_  (.A(\reg_module/_01784_ ),
    .X(\reg_module/_01835_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18654_  (.A(\reg_module/_01835_ ),
    .B(net301),
    .Y(\reg_module/_01836_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18655_  (.A1(\reg_module/_01834_ ),
    .A2(\reg_module/_01836_ ),
    .B1(\reg_module/_01830_ ),
    .Y(\reg_module/_00757_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18656_  (.A1(net2036),
    .A2(\reg_module/_01789_ ),
    .B1(net1040),
    .Y(\reg_module/_01837_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18657_  (.A1(\reg_module/_07588_ ),
    .A2(\reg_module/_01800_ ),
    .B1(\reg_module/_01837_ ),
    .Y(\reg_module/_00758_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18658_  (.A(\reg_module/_01827_ ),
    .B(net1286),
    .Y(\reg_module/_01838_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18659_  (.A(\reg_module/_01835_ ),
    .B(net299),
    .Y(\reg_module/_01839_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18660_  (.A1(\reg_module/_01838_ ),
    .A2(\reg_module/_01839_ ),
    .B1(\reg_module/_01830_ ),
    .Y(\reg_module/_00759_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18661_  (.A1(net1826),
    .A2(\reg_module/_01789_ ),
    .B1(net1014),
    .Y(\reg_module/_01840_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18662_  (.A1(\reg_module/_07595_ ),
    .A2(\reg_module/_01800_ ),
    .B1(\reg_module/_01840_ ),
    .Y(\reg_module/_00760_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18663_  (.A(\reg_module/_01827_ ),
    .B(net1281),
    .Y(\reg_module/_01841_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18664_  (.A(\reg_module/_01835_ ),
    .B(net297),
    .Y(\reg_module/_01842_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18665_  (.A1(\reg_module/_01841_ ),
    .A2(\reg_module/_01842_ ),
    .B1(\reg_module/_01830_ ),
    .Y(\reg_module/_00761_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18666_  (.A(\reg_module/_01827_ ),
    .B(net1964),
    .Y(\reg_module/_01843_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18667_  (.A(\reg_module/_01835_ ),
    .B(net295),
    .Y(\reg_module/_01844_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18668_  (.A1(\reg_module/_01843_ ),
    .A2(\reg_module/_01844_ ),
    .B1(\reg_module/_01830_ ),
    .Y(\reg_module/_00762_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18669_  (.A(\reg_module/_01785_ ),
    .B(net1364),
    .Y(\reg_module/_01845_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18670_  (.A(\reg_module/_01835_ ),
    .B(net293),
    .Y(\reg_module/_01846_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18671_  (.A(\reg_module/_01771_ ),
    .X(\reg_module/_01847_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18672_  (.A1(\reg_module/_01845_ ),
    .A2(\reg_module/_01846_ ),
    .B1(\reg_module/_01847_ ),
    .Y(\reg_module/_00763_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18673_  (.A1(net1685),
    .A2(\reg_module/_01789_ ),
    .B1(net1012),
    .Y(\reg_module/_01848_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18674_  (.A1(\reg_module/_07607_ ),
    .A2(\reg_module/_01800_ ),
    .B1(\reg_module/_01848_ ),
    .Y(\reg_module/_00764_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18675_  (.A(\reg_module/_01785_ ),
    .B(net1505),
    .Y(\reg_module/_01849_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18676_  (.A(\reg_module/_01835_ ),
    .B(net291),
    .Y(\reg_module/_01850_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18677_  (.A1(\reg_module/_01849_ ),
    .A2(\reg_module/_01850_ ),
    .B1(\reg_module/_01847_ ),
    .Y(\reg_module/_00765_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18678_  (.A1(net1648),
    .A2(\reg_module/_01789_ ),
    .B1(net1012),
    .Y(\reg_module/_01851_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18679_  (.A1(\reg_module/_07613_ ),
    .A2(\reg_module/_01800_ ),
    .B1(\reg_module/_01851_ ),
    .Y(\reg_module/_00766_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18680_  (.A(\reg_module/_01785_ ),
    .B(\reg_module/gprf[767] ),
    .Y(\reg_module/_01852_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18681_  (.A(\reg_module/_01788_ ),
    .B(net288),
    .Y(\reg_module/_01853_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18682_  (.A1(\reg_module/_01852_ ),
    .A2(\reg_module/_01853_ ),
    .B1(\reg_module/_01847_ ),
    .Y(\reg_module/_00767_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_18683_  (.A(\reg_module/_08836_ ),
    .B(\reg_module/_01154_ ),
    .Y(\reg_module/_01854_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18684_  (.A(\reg_module/_01854_ ),
    .X(\reg_module/_01855_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18685_  (.A(\reg_module/_01854_ ),
    .X(\reg_module/_01856_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18686_  (.A1(net1740),
    .A2(\reg_module/_01856_ ),
    .B1(net1039),
    .Y(\reg_module/_01857_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18687_  (.A1(\reg_module/_07514_ ),
    .A2(\reg_module/_01855_ ),
    .B1(\reg_module/_01857_ ),
    .Y(\reg_module/_00768_ ));
 sky130_fd_sc_hd__inv_4 \reg_module/_18688_  (.A(\reg_module/_01854_ ),
    .Y(\reg_module/_01858_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18689_  (.A(\reg_module/_01858_ ),
    .X(\reg_module/_01859_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18690_  (.A(\reg_module/_01859_ ),
    .B(net1559),
    .Y(\reg_module/_01860_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18691_  (.A(\reg_module/_01778_ ),
    .B(\reg_module/_08839_ ),
    .Y(\reg_module/_01861_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18692_  (.A1(\reg_module/_01860_ ),
    .A2(\reg_module/_01861_ ),
    .B1(\reg_module/_01847_ ),
    .Y(\reg_module/_00769_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18693_  (.A(\reg_module/_01859_ ),
    .B(net1305),
    .Y(\reg_module/_01862_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18694_  (.A(\reg_module/_01778_ ),
    .B(\reg_module/_08842_ ),
    .Y(\reg_module/_01863_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18695_  (.A1(\reg_module/_01862_ ),
    .A2(\reg_module/_01863_ ),
    .B1(\reg_module/_01847_ ),
    .Y(\reg_module/_00770_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18696_  (.A1(net1936),
    .A2(\reg_module/_01856_ ),
    .B1(net1042),
    .Y(\reg_module/_01864_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18697_  (.A1(\reg_module/_07523_ ),
    .A2(\reg_module/_01855_ ),
    .B1(\reg_module/_01864_ ),
    .Y(\reg_module/_00771_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18698_  (.A(\reg_module/_01859_ ),
    .B(net1681),
    .Y(\reg_module/_01865_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18699_  (.A(\reg_module/_01778_ ),
    .B(\reg_module/_08849_ ),
    .Y(\reg_module/_01866_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18700_  (.A1(\reg_module/_01865_ ),
    .A2(\reg_module/_01866_ ),
    .B1(\reg_module/_01847_ ),
    .Y(\reg_module/_00772_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18701_  (.A(\reg_module/_01859_ ),
    .B(net1583),
    .Y(\reg_module/_01867_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18702_  (.A(\reg_module/_01300_ ),
    .X(\reg_module/_01868_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18703_  (.A(\reg_module/_01868_ ),
    .X(\reg_module/_01869_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18704_  (.A(\reg_module/_01869_ ),
    .B(\reg_module/_08853_ ),
    .Y(\reg_module/_01870_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18705_  (.A(\reg_module/_01771_ ),
    .X(\reg_module/_01871_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18706_  (.A1(\reg_module/_01867_ ),
    .A2(\reg_module/_01870_ ),
    .B1(\reg_module/_01871_ ),
    .Y(\reg_module/_00773_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18707_  (.A(\reg_module/_01859_ ),
    .B(net1476),
    .Y(\reg_module/_01872_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18708_  (.A(\reg_module/_01869_ ),
    .B(\reg_module/_08856_ ),
    .Y(\reg_module/_01873_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18709_  (.A1(\reg_module/_01872_ ),
    .A2(\reg_module/_01873_ ),
    .B1(\reg_module/_01871_ ),
    .Y(\reg_module/_00774_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18710_  (.A(\reg_module/_01859_ ),
    .B(net1974),
    .Y(\reg_module/_01874_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18711_  (.A(\reg_module/_01869_ ),
    .B(\reg_module/_08859_ ),
    .Y(\reg_module/_01875_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18712_  (.A1(\reg_module/_01874_ ),
    .A2(\reg_module/_01875_ ),
    .B1(\reg_module/_01871_ ),
    .Y(\reg_module/_00775_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18713_  (.A(\reg_module/_01858_ ),
    .X(\reg_module/_01876_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18714_  (.A(\reg_module/_01876_ ),
    .B(net1347),
    .Y(\reg_module/_01877_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18715_  (.A(\reg_module/_01869_ ),
    .B(\reg_module/_08864_ ),
    .Y(\reg_module/_01878_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18716_  (.A1(\reg_module/_01877_ ),
    .A2(\reg_module/_01878_ ),
    .B1(\reg_module/_01871_ ),
    .Y(\reg_module/_00776_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18717_  (.A(\reg_module/_01876_ ),
    .B(net1448),
    .Y(\reg_module/_01879_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18718_  (.A(\reg_module/_01869_ ),
    .B(\reg_module/_08867_ ),
    .Y(\reg_module/_01880_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18719_  (.A1(\reg_module/_01879_ ),
    .A2(\reg_module/_01880_ ),
    .B1(\reg_module/_01871_ ),
    .Y(\reg_module/_00777_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18720_  (.A1(net1698),
    .A2(\reg_module/_01856_ ),
    .B1(net1053),
    .Y(\reg_module/_01881_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18721_  (.A1(\reg_module/_07548_ ),
    .A2(\reg_module/_01855_ ),
    .B1(\reg_module/_01881_ ),
    .Y(\reg_module/_00778_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18722_  (.A(\reg_module/_01876_ ),
    .B(net1769),
    .Y(\reg_module/_01882_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18723_  (.A(\reg_module/_01869_ ),
    .B(\reg_module/_08875_ ),
    .Y(\reg_module/_01883_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18724_  (.A1(\reg_module/_01882_ ),
    .A2(\reg_module/_01883_ ),
    .B1(\reg_module/_01871_ ),
    .Y(\reg_module/_00779_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18725_  (.A(\reg_module/_01876_ ),
    .B(net1904),
    .Y(\reg_module/_01884_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18726_  (.A(\reg_module/_01868_ ),
    .X(\reg_module/_01885_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18727_  (.A(\reg_module/_01885_ ),
    .B(\reg_module/_08880_ ),
    .Y(\reg_module/_01886_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18728_  (.A(\reg_module/_01506_ ),
    .X(\reg_module/_01887_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18729_  (.A(\reg_module/_01887_ ),
    .X(\reg_module/_01888_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18730_  (.A1(\reg_module/_01884_ ),
    .A2(\reg_module/_01886_ ),
    .B1(\reg_module/_01888_ ),
    .Y(\reg_module/_00780_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18731_  (.A1(net1706),
    .A2(\reg_module/_01856_ ),
    .B1(net1066),
    .Y(\reg_module/_01889_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18732_  (.A1(\reg_module/_07558_ ),
    .A2(\reg_module/_01855_ ),
    .B1(\reg_module/_01889_ ),
    .Y(\reg_module/_00781_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18733_  (.A(\reg_module/_01876_ ),
    .B(net1490),
    .Y(\reg_module/_01890_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18734_  (.A(\reg_module/_01885_ ),
    .B(\reg_module/_08886_ ),
    .Y(\reg_module/_01891_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18735_  (.A1(\reg_module/_01890_ ),
    .A2(\reg_module/_01891_ ),
    .B1(\reg_module/_01888_ ),
    .Y(\reg_module/_00782_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18736_  (.A(\reg_module/_01876_ ),
    .B(net1419),
    .Y(\reg_module/_01892_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18737_  (.A(\reg_module/_01885_ ),
    .B(\reg_module/_08889_ ),
    .Y(\reg_module/_01893_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18738_  (.A1(\reg_module/_01892_ ),
    .A2(\reg_module/_01893_ ),
    .B1(\reg_module/_01888_ ),
    .Y(\reg_module/_00783_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18739_  (.A(\reg_module/_01858_ ),
    .X(\reg_module/_01894_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18740_  (.A(\reg_module/_01894_ ),
    .B(net1340),
    .Y(\reg_module/_01895_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18741_  (.A(\reg_module/_01885_ ),
    .B(\reg_module/_08894_ ),
    .Y(\reg_module/_01896_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18742_  (.A1(\reg_module/_01895_ ),
    .A2(\reg_module/_01896_ ),
    .B1(\reg_module/_01888_ ),
    .Y(\reg_module/_00784_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18743_  (.A(\reg_module/_01894_ ),
    .B(net1535),
    .Y(\reg_module/_01897_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18744_  (.A(\reg_module/_01885_ ),
    .B(\reg_module/_08897_ ),
    .Y(\reg_module/_01898_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18745_  (.A1(\reg_module/_01897_ ),
    .A2(\reg_module/_01898_ ),
    .B1(\reg_module/_01888_ ),
    .Y(\reg_module/_00785_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18746_  (.A1(net2005),
    .A2(\reg_module/_01856_ ),
    .B1(net1058),
    .Y(\reg_module/_01899_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18747_  (.A1(\reg_module/_07575_ ),
    .A2(\reg_module/_01855_ ),
    .B1(\reg_module/_01899_ ),
    .Y(\reg_module/_00786_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18748_  (.A(\reg_module/_01894_ ),
    .B(net2129),
    .Y(\reg_module/_01900_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18749_  (.A(\reg_module/_01885_ ),
    .B(\reg_module/_08904_ ),
    .Y(\reg_module/_01901_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18750_  (.A1(\reg_module/_01900_ ),
    .A2(\reg_module/_01901_ ),
    .B1(\reg_module/_01888_ ),
    .Y(\reg_module/_00787_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18751_  (.A(\reg_module/_01894_ ),
    .B(net1878),
    .Y(\reg_module/_01902_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18752_  (.A(\reg_module/_01868_ ),
    .X(\reg_module/_01903_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18753_  (.A(\reg_module/_01903_ ),
    .B(\reg_module/_08908_ ),
    .Y(\reg_module/_01904_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18754_  (.A(\reg_module/_01887_ ),
    .X(\reg_module/_01905_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18755_  (.A1(\reg_module/_01902_ ),
    .A2(\reg_module/_01904_ ),
    .B1(\reg_module/_01905_ ),
    .Y(\reg_module/_00788_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18756_  (.A(\reg_module/_01894_ ),
    .B(net1349),
    .Y(\reg_module/_01906_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18757_  (.A(\reg_module/_01903_ ),
    .B(\reg_module/_08911_ ),
    .Y(\reg_module/_01907_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18758_  (.A1(\reg_module/_01906_ ),
    .A2(\reg_module/_01907_ ),
    .B1(\reg_module/_01905_ ),
    .Y(\reg_module/_00789_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18759_  (.A(\reg_module/_01894_ ),
    .B(net1497),
    .Y(\reg_module/_01908_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18760_  (.A(\reg_module/_01903_ ),
    .B(\reg_module/_08914_ ),
    .Y(\reg_module/_01909_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18761_  (.A1(\reg_module/_01908_ ),
    .A2(\reg_module/_01909_ ),
    .B1(\reg_module/_01905_ ),
    .Y(\reg_module/_00790_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18762_  (.A1(net2144),
    .A2(\reg_module/_01856_ ),
    .B1(net1058),
    .Y(\reg_module/_01910_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18763_  (.A1(\reg_module/_07591_ ),
    .A2(\reg_module/_01855_ ),
    .B1(\reg_module/_01910_ ),
    .Y(\reg_module/_00791_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18764_  (.A(\reg_module/_01858_ ),
    .X(\reg_module/_01911_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18765_  (.A(\reg_module/_01911_ ),
    .B(net1515),
    .Y(\reg_module/_01912_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18766_  (.A(\reg_module/_01903_ ),
    .B(\reg_module/_08922_ ),
    .Y(\reg_module/_01913_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18767_  (.A1(\reg_module/_01912_ ),
    .A2(\reg_module/_01913_ ),
    .B1(\reg_module/_01905_ ),
    .Y(\reg_module/_00792_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18768_  (.A(\reg_module/_01911_ ),
    .B(net1354),
    .Y(\reg_module/_01914_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18769_  (.A(\reg_module/_01903_ ),
    .B(\reg_module/_08925_ ),
    .Y(\reg_module/_01915_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18770_  (.A1(\reg_module/_01914_ ),
    .A2(\reg_module/_01915_ ),
    .B1(\reg_module/_01905_ ),
    .Y(\reg_module/_00793_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18771_  (.A(\reg_module/_01911_ ),
    .B(net1366),
    .Y(\reg_module/_01916_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18772_  (.A(\reg_module/_01903_ ),
    .B(\reg_module/_08929_ ),
    .Y(\reg_module/_01917_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18773_  (.A1(\reg_module/_01916_ ),
    .A2(\reg_module/_01917_ ),
    .B1(\reg_module/_01905_ ),
    .Y(\reg_module/_00794_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18774_  (.A(\reg_module/_01911_ ),
    .B(net1300),
    .Y(\reg_module/_01918_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18775_  (.A(\reg_module/_01868_ ),
    .X(\reg_module/_01919_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18776_  (.A(\reg_module/_01919_ ),
    .B(\reg_module/_08933_ ),
    .Y(\reg_module/_01920_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18777_  (.A(\reg_module/_01887_ ),
    .X(\reg_module/_01921_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18778_  (.A1(\reg_module/_01918_ ),
    .A2(\reg_module/_01920_ ),
    .B1(\reg_module/_01921_ ),
    .Y(\reg_module/_00795_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18779_  (.A(\reg_module/_01911_ ),
    .B(net1264),
    .Y(\reg_module/_01922_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18780_  (.A(\reg_module/_01919_ ),
    .B(\reg_module/_08936_ ),
    .Y(\reg_module/_01923_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18781_  (.A1(\reg_module/_01922_ ),
    .A2(\reg_module/_01923_ ),
    .B1(\reg_module/_01921_ ),
    .Y(\reg_module/_00796_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18782_  (.A(\reg_module/_01911_ ),
    .B(net1502),
    .Y(\reg_module/_01924_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18783_  (.A(\reg_module/_01919_ ),
    .B(\reg_module/_08939_ ),
    .Y(\reg_module/_01925_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18784_  (.A1(\reg_module/_01924_ ),
    .A2(\reg_module/_01925_ ),
    .B1(\reg_module/_01921_ ),
    .Y(\reg_module/_00797_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18785_  (.A(\reg_module/_01858_ ),
    .B(net1342),
    .Y(\reg_module/_01926_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18786_  (.A(\reg_module/_01919_ ),
    .B(\reg_module/_08942_ ),
    .Y(\reg_module/_01927_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18787_  (.A1(\reg_module/_01926_ ),
    .A2(\reg_module/_01927_ ),
    .B1(\reg_module/_01921_ ),
    .Y(\reg_module/_00798_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18788_  (.A(\reg_module/_01858_ ),
    .B(net1346),
    .Y(\reg_module/_01928_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18789_  (.A(\reg_module/_01919_ ),
    .B(\reg_module/_08945_ ),
    .Y(\reg_module/_01929_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18790_  (.A1(\reg_module/_01928_ ),
    .A2(\reg_module/_01929_ ),
    .B1(\reg_module/_01921_ ),
    .Y(\reg_module/_00799_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18791_  (.A(\reg_module/_08956_ ),
    .B(\reg_module/_01750_ ),
    .Y(\reg_module/_01930_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18792_  (.A(\reg_module/_07647_ ),
    .B(\reg_module/_07626_ ),
    .Y(\reg_module/_01931_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_18793_  (.A(\reg_module/_01931_ ),
    .X(\reg_module/_01932_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18794_  (.A(\reg_module/_01932_ ),
    .X(\reg_module/_01933_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18795_  (.A1(\reg_module/_01275_ ),
    .A2(\reg_module/_01933_ ),
    .B1(net1821),
    .Y(\reg_module/_01934_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18796_  (.A1(\reg_module/_01930_ ),
    .A2(\reg_module/_01934_ ),
    .B1(\reg_module/_01921_ ),
    .Y(\reg_module/_00800_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18797_  (.A(\reg_module/_08962_ ),
    .B(\reg_module/_01750_ ),
    .Y(\reg_module/_01935_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18798_  (.A1(\reg_module/_01275_ ),
    .A2(\reg_module/_01933_ ),
    .B1(net1958),
    .Y(\reg_module/_01936_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18799_  (.A(\reg_module/_01887_ ),
    .X(\reg_module/_01937_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18800_  (.A1(\reg_module/_01935_ ),
    .A2(\reg_module/_01936_ ),
    .B1(\reg_module/_01937_ ),
    .Y(\reg_module/_00801_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18801_  (.A(\reg_module/_08965_ ),
    .B(\reg_module/_01750_ ),
    .Y(\reg_module/_01938_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18802_  (.A1(\reg_module/_01275_ ),
    .A2(\reg_module/_01933_ ),
    .B1(net2026),
    .Y(\reg_module/_01939_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18803_  (.A1(\reg_module/_01938_ ),
    .A2(\reg_module/_01939_ ),
    .B1(\reg_module/_01937_ ),
    .Y(\reg_module/_00802_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18804_  (.A(\reg_module/_08968_ ),
    .B(\reg_module/_01750_ ),
    .Y(\reg_module/_01940_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18805_  (.A1(\reg_module/_01275_ ),
    .A2(\reg_module/_01933_ ),
    .B1(net2152),
    .Y(\reg_module/_01941_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18806_  (.A1(\reg_module/_01940_ ),
    .A2(\reg_module/_01941_ ),
    .B1(\reg_module/_01937_ ),
    .Y(\reg_module/_00803_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18807_  (.A(\reg_module/_01408_ ),
    .X(\reg_module/_01942_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18808_  (.A(\reg_module/_08971_ ),
    .B(\reg_module/_01942_ ),
    .Y(\reg_module/_01943_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18809_  (.A(\reg_module/_01254_ ),
    .X(\reg_module/_01944_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18810_  (.A1(\reg_module/_01944_ ),
    .A2(\reg_module/_01933_ ),
    .B1(net1930),
    .Y(\reg_module/_01945_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18811_  (.A1(\reg_module/_01943_ ),
    .A2(\reg_module/_01945_ ),
    .B1(\reg_module/_01937_ ),
    .Y(\reg_module/_00804_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18812_  (.A(\reg_module/_08975_ ),
    .B(\reg_module/_01942_ ),
    .Y(\reg_module/_01946_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18813_  (.A1(\reg_module/_01944_ ),
    .A2(\reg_module/_01933_ ),
    .B1(net1914),
    .Y(\reg_module/_01947_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18814_  (.A1(\reg_module/_01946_ ),
    .A2(\reg_module/_01947_ ),
    .B1(\reg_module/_01937_ ),
    .Y(\reg_module/_00805_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18815_  (.A(\reg_module/_08980_ ),
    .B(\reg_module/_01942_ ),
    .Y(\reg_module/_01948_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18816_  (.A(\reg_module/_01932_ ),
    .X(\reg_module/_01949_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18817_  (.A1(\reg_module/_01944_ ),
    .A2(\reg_module/_01949_ ),
    .B1(net1912),
    .Y(\reg_module/_01950_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18818_  (.A1(\reg_module/_01948_ ),
    .A2(\reg_module/_01950_ ),
    .B1(\reg_module/_01937_ ),
    .Y(\reg_module/_00806_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18819_  (.A(\reg_module/_08984_ ),
    .B(\reg_module/_01942_ ),
    .Y(\reg_module/_01951_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18820_  (.A1(\reg_module/_01944_ ),
    .A2(\reg_module/_01949_ ),
    .B1(net1798),
    .Y(\reg_module/_01952_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18821_  (.A(\reg_module/_01887_ ),
    .X(\reg_module/_01953_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18822_  (.A1(\reg_module/_01951_ ),
    .A2(\reg_module/_01952_ ),
    .B1(\reg_module/_01953_ ),
    .Y(\reg_module/_00807_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18823_  (.A(\reg_module/_08987_ ),
    .B(\reg_module/_01942_ ),
    .Y(\reg_module/_01954_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18824_  (.A1(\reg_module/_01944_ ),
    .A2(\reg_module/_01949_ ),
    .B1(net1795),
    .Y(\reg_module/_01955_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18825_  (.A1(\reg_module/_01954_ ),
    .A2(\reg_module/_01955_ ),
    .B1(\reg_module/_01953_ ),
    .Y(\reg_module/_00808_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18826_  (.A(\reg_module/_08990_ ),
    .B(\reg_module/_01942_ ),
    .Y(\reg_module/_01956_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18827_  (.A1(\reg_module/_01944_ ),
    .A2(\reg_module/_01949_ ),
    .B1(net1911),
    .Y(\reg_module/_01957_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18828_  (.A1(\reg_module/_01956_ ),
    .A2(\reg_module/_01957_ ),
    .B1(\reg_module/_01953_ ),
    .Y(\reg_module/_00809_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18829_  (.A(\reg_module/_01408_ ),
    .X(\reg_module/_01958_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18830_  (.A(\reg_module/_08993_ ),
    .B(\reg_module/_01958_ ),
    .Y(\reg_module/_01959_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18831_  (.A(\reg_module/_01254_ ),
    .X(\reg_module/_01960_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18832_  (.A1(\reg_module/_01960_ ),
    .A2(\reg_module/_01949_ ),
    .B1(net1898),
    .Y(\reg_module/_01961_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18833_  (.A1(\reg_module/_01959_ ),
    .A2(\reg_module/_01961_ ),
    .B1(\reg_module/_01953_ ),
    .Y(\reg_module/_00810_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18834_  (.A(\reg_module/_08998_ ),
    .B(\reg_module/_01958_ ),
    .Y(\reg_module/_01962_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18835_  (.A1(\reg_module/_01960_ ),
    .A2(\reg_module/_01949_ ),
    .B1(net1989),
    .Y(\reg_module/_01963_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18836_  (.A1(\reg_module/_01962_ ),
    .A2(\reg_module/_01963_ ),
    .B1(\reg_module/_01953_ ),
    .Y(\reg_module/_00811_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18837_  (.A(\reg_module/_09003_ ),
    .B(\reg_module/_01958_ ),
    .Y(\reg_module/_01964_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18838_  (.A(\reg_module/_01932_ ),
    .X(\reg_module/_01965_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18839_  (.A1(\reg_module/_01960_ ),
    .A2(\reg_module/_01965_ ),
    .B1(net2128),
    .Y(\reg_module/_01966_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18840_  (.A1(\reg_module/_01964_ ),
    .A2(\reg_module/_01966_ ),
    .B1(\reg_module/_01953_ ),
    .Y(\reg_module/_00812_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18841_  (.A(\reg_module/_09007_ ),
    .B(\reg_module/_01958_ ),
    .Y(\reg_module/_01967_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18842_  (.A1(\reg_module/_01960_ ),
    .A2(\reg_module/_01965_ ),
    .B1(net2141),
    .Y(\reg_module/_01968_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18843_  (.A(\reg_module/_01887_ ),
    .X(\reg_module/_01969_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18844_  (.A1(\reg_module/_01967_ ),
    .A2(\reg_module/_01968_ ),
    .B1(\reg_module/_01969_ ),
    .Y(\reg_module/_00813_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18845_  (.A(\reg_module/_09010_ ),
    .B(\reg_module/_01958_ ),
    .Y(\reg_module/_01970_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18846_  (.A1(\reg_module/_01960_ ),
    .A2(\reg_module/_01965_ ),
    .B1(net2046),
    .Y(\reg_module/_01971_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18847_  (.A1(\reg_module/_01970_ ),
    .A2(\reg_module/_01971_ ),
    .B1(\reg_module/_01969_ ),
    .Y(\reg_module/_00814_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18848_  (.A(\reg_module/_09013_ ),
    .B(\reg_module/_01958_ ),
    .Y(\reg_module/_01972_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18849_  (.A1(\reg_module/_01960_ ),
    .A2(\reg_module/_01965_ ),
    .B1(net2030),
    .Y(\reg_module/_01973_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18850_  (.A1(\reg_module/_01972_ ),
    .A2(\reg_module/_01973_ ),
    .B1(\reg_module/_01969_ ),
    .Y(\reg_module/_00815_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_18851_  (.A(\reg_module/_01381_ ),
    .X(\reg_module/_01974_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18852_  (.A(\reg_module/_01974_ ),
    .X(\reg_module/_01975_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18853_  (.A(\reg_module/_09016_ ),
    .B(\reg_module/_01975_ ),
    .Y(\reg_module/_01976_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18854_  (.A(\reg_module/_01254_ ),
    .X(\reg_module/_01977_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18855_  (.A1(\reg_module/_01977_ ),
    .A2(\reg_module/_01965_ ),
    .B1(net2100),
    .Y(\reg_module/_01978_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18856_  (.A1(\reg_module/_01976_ ),
    .A2(\reg_module/_01978_ ),
    .B1(\reg_module/_01969_ ),
    .Y(\reg_module/_00816_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18857_  (.A(\reg_module/_09020_ ),
    .B(\reg_module/_01975_ ),
    .Y(\reg_module/_01979_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18858_  (.A1(\reg_module/_01977_ ),
    .A2(\reg_module/_01965_ ),
    .B1(net2076),
    .Y(\reg_module/_01980_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18859_  (.A1(\reg_module/_01979_ ),
    .A2(\reg_module/_01980_ ),
    .B1(\reg_module/_01969_ ),
    .Y(\reg_module/_00817_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18860_  (.A(\reg_module/_09025_ ),
    .B(\reg_module/_01975_ ),
    .Y(\reg_module/_01981_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18861_  (.A(\reg_module/_01932_ ),
    .X(\reg_module/_01982_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18862_  (.A1(\reg_module/_01977_ ),
    .A2(\reg_module/_01982_ ),
    .B1(net2047),
    .Y(\reg_module/_01983_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18863_  (.A1(\reg_module/_01981_ ),
    .A2(\reg_module/_01983_ ),
    .B1(\reg_module/_01969_ ),
    .Y(\reg_module/_00818_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18864_  (.A(\reg_module/_09030_ ),
    .B(\reg_module/_01975_ ),
    .Y(\reg_module/_01984_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18865_  (.A1(\reg_module/_01977_ ),
    .A2(\reg_module/_01982_ ),
    .B1(net2044),
    .Y(\reg_module/_01985_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18866_  (.A(\reg_module/_01506_ ),
    .X(\reg_module/_01986_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18867_  (.A(\reg_module/_01986_ ),
    .X(\reg_module/_01987_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18868_  (.A1(\reg_module/_01984_ ),
    .A2(\reg_module/_01985_ ),
    .B1(\reg_module/_01987_ ),
    .Y(\reg_module/_00819_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18869_  (.A(\reg_module/_09033_ ),
    .B(\reg_module/_01975_ ),
    .Y(\reg_module/_01988_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18870_  (.A1(\reg_module/_01977_ ),
    .A2(\reg_module/_01982_ ),
    .B1(net2153),
    .Y(\reg_module/_01989_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18871_  (.A1(\reg_module/_01988_ ),
    .A2(\reg_module/_01989_ ),
    .B1(\reg_module/_01987_ ),
    .Y(\reg_module/_00820_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18872_  (.A(\reg_module/_09036_ ),
    .B(\reg_module/_01975_ ),
    .Y(\reg_module/_01990_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18873_  (.A1(\reg_module/_01977_ ),
    .A2(\reg_module/_01982_ ),
    .B1(net2096),
    .Y(\reg_module/_01991_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18874_  (.A1(\reg_module/_01990_ ),
    .A2(\reg_module/_01991_ ),
    .B1(\reg_module/_01987_ ),
    .Y(\reg_module/_00821_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_18875_  (.A(\reg_module/_01974_ ),
    .X(\reg_module/_01992_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18876_  (.A(\reg_module/_09039_ ),
    .B(\reg_module/_01992_ ),
    .Y(\reg_module/_01993_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18877_  (.A(\reg_module/_01254_ ),
    .X(\reg_module/_01994_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18878_  (.A1(\reg_module/_01994_ ),
    .A2(\reg_module/_01982_ ),
    .B1(net2091),
    .Y(\reg_module/_01995_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18879_  (.A1(\reg_module/_01993_ ),
    .A2(\reg_module/_01995_ ),
    .B1(\reg_module/_01987_ ),
    .Y(\reg_module/_00822_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18880_  (.A(\reg_module/_09043_ ),
    .B(\reg_module/_01992_ ),
    .Y(\reg_module/_01996_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18881_  (.A1(\reg_module/_01994_ ),
    .A2(\reg_module/_01982_ ),
    .B1(net2187),
    .Y(\reg_module/_01997_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18882_  (.A1(\reg_module/_01996_ ),
    .A2(\reg_module/_01997_ ),
    .B1(\reg_module/_01987_ ),
    .Y(\reg_module/_00823_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18883_  (.A(\reg_module/_09049_ ),
    .B(\reg_module/_01992_ ),
    .Y(\reg_module/_01998_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18884_  (.A(\reg_module/_01931_ ),
    .X(\reg_module/_01999_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18885_  (.A1(\reg_module/_01994_ ),
    .A2(\reg_module/_01999_ ),
    .B1(net1760),
    .Y(\reg_module/_02000_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18886_  (.A1(\reg_module/_01998_ ),
    .A2(\reg_module/_02000_ ),
    .B1(\reg_module/_01987_ ),
    .Y(\reg_module/_00824_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18887_  (.A(\reg_module/_09053_ ),
    .B(\reg_module/_01992_ ),
    .Y(\reg_module/_02001_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18888_  (.A1(\reg_module/_01994_ ),
    .A2(\reg_module/_01999_ ),
    .B1(net1673),
    .Y(\reg_module/_02002_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18889_  (.A(\reg_module/_01986_ ),
    .X(\reg_module/_02003_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18890_  (.A1(\reg_module/_02001_ ),
    .A2(\reg_module/_02002_ ),
    .B1(\reg_module/_02003_ ),
    .Y(\reg_module/_00825_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18891_  (.A(\reg_module/_09056_ ),
    .B(\reg_module/_01992_ ),
    .Y(\reg_module/_02004_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18892_  (.A1(\reg_module/_01994_ ),
    .A2(\reg_module/_01999_ ),
    .B1(net1790),
    .Y(\reg_module/_02005_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18893_  (.A1(\reg_module/_02004_ ),
    .A2(\reg_module/_02005_ ),
    .B1(\reg_module/_02003_ ),
    .Y(\reg_module/_00826_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18894_  (.A(\reg_module/_09059_ ),
    .B(\reg_module/_01992_ ),
    .Y(\reg_module/_02006_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18895_  (.A1(\reg_module/_01994_ ),
    .A2(\reg_module/_01999_ ),
    .B1(net1923),
    .Y(\reg_module/_02007_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18896_  (.A1(\reg_module/_02006_ ),
    .A2(\reg_module/_02007_ ),
    .B1(\reg_module/_02003_ ),
    .Y(\reg_module/_00827_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18897_  (.A(\reg_module/_01974_ ),
    .X(\reg_module/_02008_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18898_  (.A(\reg_module/_09062_ ),
    .B(\reg_module/_02008_ ),
    .Y(\reg_module/_02009_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18899_  (.A(\reg_module/_01154_ ),
    .X(\reg_module/_02010_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18900_  (.A(\reg_module/_02010_ ),
    .X(\reg_module/_02011_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18901_  (.A1(\reg_module/_02011_ ),
    .A2(\reg_module/_01999_ ),
    .B1(net1808),
    .Y(\reg_module/_02012_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18902_  (.A1(\reg_module/_02009_ ),
    .A2(\reg_module/_02012_ ),
    .B1(\reg_module/_02003_ ),
    .Y(\reg_module/_00828_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18903_  (.A(\reg_module/_09066_ ),
    .B(\reg_module/_02008_ ),
    .Y(\reg_module/_02013_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18904_  (.A1(\reg_module/_02011_ ),
    .A2(\reg_module/_01999_ ),
    .B1(net1730),
    .Y(\reg_module/_02014_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18905_  (.A1(\reg_module/_02013_ ),
    .A2(\reg_module/_02014_ ),
    .B1(\reg_module/_02003_ ),
    .Y(\reg_module/_00829_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18906_  (.A(\reg_module/_09070_ ),
    .B(\reg_module/_02008_ ),
    .Y(\reg_module/_02015_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18907_  (.A1(\reg_module/_02011_ ),
    .A2(\reg_module/_01932_ ),
    .B1(net1530),
    .Y(\reg_module/_02016_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18908_  (.A1(\reg_module/_02015_ ),
    .A2(\reg_module/_02016_ ),
    .B1(\reg_module/_02003_ ),
    .Y(\reg_module/_00830_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18909_  (.A(\reg_module/_09074_ ),
    .B(\reg_module/_02008_ ),
    .Y(\reg_module/_02017_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18910_  (.A1(\reg_module/_02011_ ),
    .A2(\reg_module/_01932_ ),
    .B1(net1906),
    .Y(\reg_module/_02018_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18911_  (.A(\reg_module/_01986_ ),
    .X(\reg_module/_02019_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18912_  (.A1(\reg_module/_02017_ ),
    .A2(\reg_module/_02018_ ),
    .B1(\reg_module/_02019_ ),
    .Y(\reg_module/_00831_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18913_  (.A(\reg_module/_09081_ ),
    .B(\reg_module/_02008_ ),
    .Y(\reg_module/_02020_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_18914_  (.A(\reg_module/_09076_ ),
    .Y(\reg_module/_02021_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18915_  (.A(\reg_module/_02021_ ),
    .X(\reg_module/_02022_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18916_  (.A(\reg_module/_02022_ ),
    .X(\reg_module/_02023_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18917_  (.A1(\reg_module/_02011_ ),
    .A2(\reg_module/_02023_ ),
    .B1(net1742),
    .Y(\reg_module/_02024_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18918_  (.A1(\reg_module/_02020_ ),
    .A2(\reg_module/_02024_ ),
    .B1(\reg_module/_02019_ ),
    .Y(\reg_module/_00832_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18919_  (.A(\reg_module/_09084_ ),
    .B(\reg_module/_02008_ ),
    .Y(\reg_module/_02025_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18920_  (.A1(\reg_module/_02011_ ),
    .A2(\reg_module/_02023_ ),
    .B1(net2019),
    .Y(\reg_module/_02026_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18921_  (.A1(\reg_module/_02025_ ),
    .A2(\reg_module/_02026_ ),
    .B1(\reg_module/_02019_ ),
    .Y(\reg_module/_00833_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18922_  (.A(\reg_module/_01974_ ),
    .X(\reg_module/_02027_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18923_  (.A(\reg_module/_09087_ ),
    .B(\reg_module/_02027_ ),
    .Y(\reg_module/_02028_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18924_  (.A(\reg_module/_02010_ ),
    .X(\reg_module/_02029_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18925_  (.A1(\reg_module/_02029_ ),
    .A2(\reg_module/_02023_ ),
    .B1(net2057),
    .Y(\reg_module/_02030_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18926_  (.A1(\reg_module/_02028_ ),
    .A2(\reg_module/_02030_ ),
    .B1(\reg_module/_02019_ ),
    .Y(\reg_module/_00834_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18927_  (.A(\reg_module/_09091_ ),
    .B(\reg_module/_02027_ ),
    .Y(\reg_module/_02031_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18928_  (.A1(\reg_module/_02029_ ),
    .A2(\reg_module/_02023_ ),
    .B1(net1701),
    .Y(\reg_module/_02032_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18929_  (.A1(\reg_module/_02031_ ),
    .A2(\reg_module/_02032_ ),
    .B1(\reg_module/_02019_ ),
    .Y(\reg_module/_00835_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18930_  (.A(\reg_module/_09095_ ),
    .B(\reg_module/_02027_ ),
    .Y(\reg_module/_02033_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18931_  (.A1(\reg_module/_02029_ ),
    .A2(\reg_module/_02023_ ),
    .B1(net1929),
    .Y(\reg_module/_02034_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18932_  (.A1(\reg_module/_02033_ ),
    .A2(\reg_module/_02034_ ),
    .B1(\reg_module/_02019_ ),
    .Y(\reg_module/_00836_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18933_  (.A(\reg_module/_09099_ ),
    .B(\reg_module/_02027_ ),
    .Y(\reg_module/_02035_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18934_  (.A1(\reg_module/_02029_ ),
    .A2(\reg_module/_02023_ ),
    .B1(net1957),
    .Y(\reg_module/_02036_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18935_  (.A(\reg_module/_01986_ ),
    .X(\reg_module/_02037_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18936_  (.A1(\reg_module/_02035_ ),
    .A2(\reg_module/_02036_ ),
    .B1(\reg_module/_02037_ ),
    .Y(\reg_module/_00837_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18937_  (.A(\reg_module/_09103_ ),
    .B(\reg_module/_02027_ ),
    .Y(\reg_module/_02038_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18938_  (.A(\reg_module/_02022_ ),
    .X(\reg_module/_02039_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18939_  (.A1(\reg_module/_02029_ ),
    .A2(\reg_module/_02039_ ),
    .B1(net1733),
    .Y(\reg_module/_02040_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18940_  (.A1(\reg_module/_02038_ ),
    .A2(\reg_module/_02040_ ),
    .B1(\reg_module/_02037_ ),
    .Y(\reg_module/_00838_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18941_  (.A(\reg_module/_09106_ ),
    .B(\reg_module/_02027_ ),
    .Y(\reg_module/_02041_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18942_  (.A1(\reg_module/_02029_ ),
    .A2(\reg_module/_02039_ ),
    .B1(net1763),
    .Y(\reg_module/_02042_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18943_  (.A1(\reg_module/_02041_ ),
    .A2(\reg_module/_02042_ ),
    .B1(\reg_module/_02037_ ),
    .Y(\reg_module/_00839_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18944_  (.A(\reg_module/_01974_ ),
    .X(\reg_module/_02043_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18945_  (.A(\reg_module/_09109_ ),
    .B(\reg_module/_02043_ ),
    .Y(\reg_module/_02044_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18946_  (.A(\reg_module/_02010_ ),
    .X(\reg_module/_02045_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18947_  (.A1(\reg_module/_02045_ ),
    .A2(\reg_module/_02039_ ),
    .B1(net1954),
    .Y(\reg_module/_02046_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18948_  (.A1(\reg_module/_02044_ ),
    .A2(\reg_module/_02046_ ),
    .B1(\reg_module/_02037_ ),
    .Y(\reg_module/_00840_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18949_  (.A(\reg_module/_09113_ ),
    .B(\reg_module/_02043_ ),
    .Y(\reg_module/_02047_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18950_  (.A1(\reg_module/_02045_ ),
    .A2(\reg_module/_02039_ ),
    .B1(net1748),
    .Y(\reg_module/_02048_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18951_  (.A1(\reg_module/_02047_ ),
    .A2(\reg_module/_02048_ ),
    .B1(\reg_module/_02037_ ),
    .Y(\reg_module/_00841_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18952_  (.A(\reg_module/_09117_ ),
    .B(\reg_module/_02043_ ),
    .Y(\reg_module/_02049_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18953_  (.A1(\reg_module/_02045_ ),
    .A2(\reg_module/_02039_ ),
    .B1(net1738),
    .Y(\reg_module/_02050_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18954_  (.A1(\reg_module/_02049_ ),
    .A2(\reg_module/_02050_ ),
    .B1(\reg_module/_02037_ ),
    .Y(\reg_module/_00842_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18955_  (.A(\reg_module/_09121_ ),
    .B(\reg_module/_02043_ ),
    .Y(\reg_module/_02051_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18956_  (.A1(\reg_module/_02045_ ),
    .A2(\reg_module/_02039_ ),
    .B1(net1877),
    .Y(\reg_module/_02052_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18957_  (.A(\reg_module/_01986_ ),
    .X(\reg_module/_02053_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18958_  (.A1(\reg_module/_02051_ ),
    .A2(\reg_module/_02052_ ),
    .B1(\reg_module/_02053_ ),
    .Y(\reg_module/_00843_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18959_  (.A(\reg_module/_09125_ ),
    .B(\reg_module/_02043_ ),
    .Y(\reg_module/_02054_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18960_  (.A(\reg_module/_02022_ ),
    .X(\reg_module/_02055_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18961_  (.A1(\reg_module/_02045_ ),
    .A2(\reg_module/_02055_ ),
    .B1(net1843),
    .Y(\reg_module/_02056_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18962_  (.A1(\reg_module/_02054_ ),
    .A2(\reg_module/_02056_ ),
    .B1(\reg_module/_02053_ ),
    .Y(\reg_module/_00844_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18963_  (.A(\reg_module/_09128_ ),
    .B(\reg_module/_02043_ ),
    .Y(\reg_module/_02057_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18964_  (.A1(\reg_module/_02045_ ),
    .A2(\reg_module/_02055_ ),
    .B1(net1942),
    .Y(\reg_module/_02058_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18965_  (.A1(\reg_module/_02057_ ),
    .A2(\reg_module/_02058_ ),
    .B1(\reg_module/_02053_ ),
    .Y(\reg_module/_00845_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18966_  (.A(\reg_module/_01974_ ),
    .X(\reg_module/_02059_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18967_  (.A(\reg_module/_09131_ ),
    .B(\reg_module/_02059_ ),
    .Y(\reg_module/_02060_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18968_  (.A(\reg_module/_02010_ ),
    .X(\reg_module/_02061_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18969_  (.A1(\reg_module/_02061_ ),
    .A2(\reg_module/_02055_ ),
    .B1(net1941),
    .Y(\reg_module/_02062_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18970_  (.A1(\reg_module/_02060_ ),
    .A2(\reg_module/_02062_ ),
    .B1(\reg_module/_02053_ ),
    .Y(\reg_module/_00846_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18971_  (.A(\reg_module/_09136_ ),
    .B(\reg_module/_02059_ ),
    .Y(\reg_module/_02063_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18972_  (.A1(\reg_module/_02061_ ),
    .A2(\reg_module/_02055_ ),
    .B1(net1782),
    .Y(\reg_module/_02064_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18973_  (.A1(\reg_module/_02063_ ),
    .A2(\reg_module/_02064_ ),
    .B1(\reg_module/_02053_ ),
    .Y(\reg_module/_00847_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18974_  (.A(\reg_module/_09140_ ),
    .B(\reg_module/_02059_ ),
    .Y(\reg_module/_02065_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18975_  (.A1(\reg_module/_02061_ ),
    .A2(\reg_module/_02055_ ),
    .B1(net1784),
    .Y(\reg_module/_02066_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18976_  (.A1(\reg_module/_02065_ ),
    .A2(\reg_module/_02066_ ),
    .B1(\reg_module/_02053_ ),
    .Y(\reg_module/_00848_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18977_  (.A(\reg_module/_09144_ ),
    .B(\reg_module/_02059_ ),
    .Y(\reg_module/_02067_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18978_  (.A1(\reg_module/_02061_ ),
    .A2(\reg_module/_02055_ ),
    .B1(net1908),
    .Y(\reg_module/_02068_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18979_  (.A(\reg_module/_01986_ ),
    .X(\reg_module/_02069_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18980_  (.A1(\reg_module/_02067_ ),
    .A2(\reg_module/_02068_ ),
    .B1(\reg_module/_02069_ ),
    .Y(\reg_module/_00849_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18981_  (.A(\reg_module/_09148_ ),
    .B(\reg_module/_02059_ ),
    .Y(\reg_module/_02070_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_18982_  (.A(\reg_module/_02022_ ),
    .X(\reg_module/_02071_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18983_  (.A1(\reg_module/_02061_ ),
    .A2(\reg_module/_02071_ ),
    .B1(net1931),
    .Y(\reg_module/_02072_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18984_  (.A1(\reg_module/_02070_ ),
    .A2(\reg_module/_02072_ ),
    .B1(\reg_module/_02069_ ),
    .Y(\reg_module/_00850_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18985_  (.A(\reg_module/_09151_ ),
    .B(\reg_module/_02059_ ),
    .Y(\reg_module/_02073_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18986_  (.A1(\reg_module/_02061_ ),
    .A2(\reg_module/_02071_ ),
    .B1(net1893),
    .Y(\reg_module/_02074_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18987_  (.A1(\reg_module/_02073_ ),
    .A2(\reg_module/_02074_ ),
    .B1(\reg_module/_02069_ ),
    .Y(\reg_module/_00851_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_18988_  (.A(\reg_module/_01381_ ),
    .X(\reg_module/_02075_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18989_  (.A(\reg_module/_02075_ ),
    .X(\reg_module/_02076_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18990_  (.A(\reg_module/_09154_ ),
    .B(\reg_module/_02076_ ),
    .Y(\reg_module/_02077_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_18991_  (.A(\reg_module/_02010_ ),
    .X(\reg_module/_02078_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18992_  (.A1(\reg_module/_02078_ ),
    .A2(\reg_module/_02071_ ),
    .B1(net1779),
    .Y(\reg_module/_02079_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18993_  (.A1(\reg_module/_02077_ ),
    .A2(\reg_module/_02079_ ),
    .B1(\reg_module/_02069_ ),
    .Y(\reg_module/_00852_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18994_  (.A(\reg_module/_09158_ ),
    .B(\reg_module/_02076_ ),
    .Y(\reg_module/_02080_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18995_  (.A1(\reg_module/_02078_ ),
    .A2(\reg_module/_02071_ ),
    .B1(net1677),
    .Y(\reg_module/_02081_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18996_  (.A1(\reg_module/_02080_ ),
    .A2(\reg_module/_02081_ ),
    .B1(\reg_module/_02069_ ),
    .Y(\reg_module/_00853_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_18997_  (.A(\reg_module/_09162_ ),
    .B(\reg_module/_02076_ ),
    .Y(\reg_module/_02082_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_18998_  (.A1(\reg_module/_02078_ ),
    .A2(\reg_module/_02071_ ),
    .B1(net1918),
    .Y(\reg_module/_02083_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_18999_  (.A1(\reg_module/_02082_ ),
    .A2(\reg_module/_02083_ ),
    .B1(\reg_module/_02069_ ),
    .Y(\reg_module/_00854_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19000_  (.A(\reg_module/_09167_ ),
    .B(\reg_module/_02076_ ),
    .Y(\reg_module/_02084_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19001_  (.A1(\reg_module/_02078_ ),
    .A2(\reg_module/_02071_ ),
    .B1(net1885),
    .Y(\reg_module/_02085_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_19002_  (.A(\reg_module/_01506_ ),
    .X(\reg_module/_02086_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19003_  (.A(\reg_module/_02086_ ),
    .X(\reg_module/_02087_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19004_  (.A1(\reg_module/_02084_ ),
    .A2(\reg_module/_02085_ ),
    .B1(\reg_module/_02087_ ),
    .Y(\reg_module/_00855_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19005_  (.A(\reg_module/_09171_ ),
    .B(\reg_module/_02076_ ),
    .Y(\reg_module/_02088_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19006_  (.A(\reg_module/_02021_ ),
    .X(\reg_module/_02089_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19007_  (.A1(\reg_module/_02078_ ),
    .A2(\reg_module/_02089_ ),
    .B1(net1727),
    .Y(\reg_module/_02090_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19008_  (.A1(\reg_module/_02088_ ),
    .A2(\reg_module/_02090_ ),
    .B1(\reg_module/_02087_ ),
    .Y(\reg_module/_00856_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19009_  (.A(\reg_module/_09174_ ),
    .B(\reg_module/_02076_ ),
    .Y(\reg_module/_02091_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19010_  (.A1(\reg_module/_02078_ ),
    .A2(\reg_module/_02089_ ),
    .B1(net1848),
    .Y(\reg_module/_02092_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19011_  (.A1(\reg_module/_02091_ ),
    .A2(\reg_module/_02092_ ),
    .B1(\reg_module/_02087_ ),
    .Y(\reg_module/_00857_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19012_  (.A(\reg_module/_02075_ ),
    .X(\reg_module/_02093_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19013_  (.A(\reg_module/_09177_ ),
    .B(\reg_module/_02093_ ),
    .Y(\reg_module/_02094_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19014_  (.A(\reg_module/_02010_ ),
    .X(\reg_module/_02095_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19015_  (.A1(\reg_module/_02095_ ),
    .A2(\reg_module/_02089_ ),
    .B1(net1849),
    .Y(\reg_module/_02096_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19016_  (.A1(\reg_module/_02094_ ),
    .A2(\reg_module/_02096_ ),
    .B1(\reg_module/_02087_ ),
    .Y(\reg_module/_00858_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19017_  (.A(\reg_module/_09181_ ),
    .B(\reg_module/_02093_ ),
    .Y(\reg_module/_02097_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19018_  (.A1(\reg_module/_02095_ ),
    .A2(\reg_module/_02089_ ),
    .B1(net1901),
    .Y(\reg_module/_02098_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19019_  (.A1(\reg_module/_02097_ ),
    .A2(\reg_module/_02098_ ),
    .B1(\reg_module/_02087_ ),
    .Y(\reg_module/_00859_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19020_  (.A(\reg_module/_09186_ ),
    .B(\reg_module/_02093_ ),
    .Y(\reg_module/_02099_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19021_  (.A1(\reg_module/_02095_ ),
    .A2(\reg_module/_02089_ ),
    .B1(net1851),
    .Y(\reg_module/_02100_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19022_  (.A1(\reg_module/_02099_ ),
    .A2(\reg_module/_02100_ ),
    .B1(\reg_module/_02087_ ),
    .Y(\reg_module/_00860_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19023_  (.A(\reg_module/_09190_ ),
    .B(\reg_module/_02093_ ),
    .Y(\reg_module/_02101_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19024_  (.A1(\reg_module/_02095_ ),
    .A2(\reg_module/_02089_ ),
    .B1(net1874),
    .Y(\reg_module/_02102_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19025_  (.A(\reg_module/_02086_ ),
    .X(\reg_module/_02103_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19026_  (.A1(\reg_module/_02101_ ),
    .A2(\reg_module/_02102_ ),
    .B1(\reg_module/_02103_ ),
    .Y(\reg_module/_00861_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19027_  (.A(\reg_module/_09193_ ),
    .B(\reg_module/_02093_ ),
    .Y(\reg_module/_02104_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19028_  (.A1(\reg_module/_02095_ ),
    .A2(\reg_module/_02022_ ),
    .B1(net1876),
    .Y(\reg_module/_02105_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19029_  (.A1(\reg_module/_02104_ ),
    .A2(\reg_module/_02105_ ),
    .B1(\reg_module/_02103_ ),
    .Y(\reg_module/_00862_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19030_  (.A(\reg_module/_09196_ ),
    .B(\reg_module/_02093_ ),
    .Y(\reg_module/_02106_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19031_  (.A1(\reg_module/_02095_ ),
    .A2(\reg_module/_02022_ ),
    .B1(net1809),
    .Y(\reg_module/_02107_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19032_  (.A1(\reg_module/_02106_ ),
    .A2(\reg_module/_02107_ ),
    .B1(\reg_module/_02103_ ),
    .Y(\reg_module/_00863_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19033_  (.A(\reg_module/_02075_ ),
    .X(\reg_module/_02108_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19034_  (.A(\reg_module/_09206_ ),
    .B(\reg_module/_02108_ ),
    .Y(\reg_module/_02109_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19035_  (.A(\reg_module/_01300_ ),
    .B(\reg_module/_09199_ ),
    .Y(\reg_module/_02110_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_19036_  (.A(\reg_module/_02110_ ),
    .X(\reg_module/_02111_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19037_  (.A(\reg_module/_02111_ ),
    .X(\reg_module/_02112_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19038_  (.A(\reg_module/_02112_ ),
    .B(net1624),
    .Y(\reg_module/_02113_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19039_  (.A1(\reg_module/_02109_ ),
    .A2(\reg_module/_02113_ ),
    .B1(\reg_module/_02103_ ),
    .Y(\reg_module/_00864_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19040_  (.A(\reg_module/_09209_ ),
    .B(\reg_module/_02108_ ),
    .Y(\reg_module/_02114_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19041_  (.A(\reg_module/_02112_ ),
    .B(net1523),
    .Y(\reg_module/_02115_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19042_  (.A1(\reg_module/_02114_ ),
    .A2(\reg_module/_02115_ ),
    .B1(\reg_module/_02103_ ),
    .Y(\reg_module/_00865_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19043_  (.A(\reg_module/_09212_ ),
    .B(\reg_module/_02108_ ),
    .Y(\reg_module/_02116_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19044_  (.A(\reg_module/_02112_ ),
    .B(net1928),
    .Y(\reg_module/_02117_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19045_  (.A1(\reg_module/_02116_ ),
    .A2(\reg_module/_02117_ ),
    .B1(\reg_module/_02103_ ),
    .Y(\reg_module/_00866_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19046_  (.A(\reg_module/_09216_ ),
    .B(\reg_module/_02108_ ),
    .Y(\reg_module/_02118_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19047_  (.A(\reg_module/_02112_ ),
    .B(net1959),
    .Y(\reg_module/_02119_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19048_  (.A(\reg_module/_02086_ ),
    .X(\reg_module/_02120_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19049_  (.A1(\reg_module/_02118_ ),
    .A2(\reg_module/_02119_ ),
    .B1(\reg_module/_02120_ ),
    .Y(\reg_module/_00867_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19050_  (.A(\reg_module/_09219_ ),
    .B(\reg_module/_02108_ ),
    .Y(\reg_module/_02121_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19051_  (.A(\reg_module/_02112_ ),
    .B(net1938),
    .Y(\reg_module/_02122_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19052_  (.A1(\reg_module/_02121_ ),
    .A2(\reg_module/_02122_ ),
    .B1(\reg_module/_02120_ ),
    .Y(\reg_module/_00868_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19053_  (.A(\reg_module/_09222_ ),
    .B(\reg_module/_02108_ ),
    .Y(\reg_module/_02123_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19054_  (.A(\reg_module/_02112_ ),
    .B(net1872),
    .Y(\reg_module/_02124_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19055_  (.A1(\reg_module/_02123_ ),
    .A2(\reg_module/_02124_ ),
    .B1(\reg_module/_02120_ ),
    .Y(\reg_module/_00869_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19056_  (.A(\reg_module/_02075_ ),
    .X(\reg_module/_02125_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19057_  (.A(\reg_module/_09228_ ),
    .B(\reg_module/_02125_ ),
    .Y(\reg_module/_02126_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19058_  (.A(\reg_module/_02111_ ),
    .X(\reg_module/_02127_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19059_  (.A(\reg_module/_02127_ ),
    .B(net2117),
    .Y(\reg_module/_02128_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19060_  (.A1(\reg_module/_02126_ ),
    .A2(\reg_module/_02128_ ),
    .B1(\reg_module/_02120_ ),
    .Y(\reg_module/_00870_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19061_  (.A(\reg_module/_09231_ ),
    .B(\reg_module/_02125_ ),
    .Y(\reg_module/_02129_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19062_  (.A(\reg_module/_02127_ ),
    .B(net2070),
    .Y(\reg_module/_02130_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19063_  (.A1(\reg_module/_02129_ ),
    .A2(\reg_module/_02130_ ),
    .B1(\reg_module/_02120_ ),
    .Y(\reg_module/_00871_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19064_  (.A(\reg_module/_09234_ ),
    .B(\reg_module/_02125_ ),
    .Y(\reg_module/_02131_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19065_  (.A(\reg_module/_02127_ ),
    .B(net2015),
    .Y(\reg_module/_02132_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19066_  (.A1(\reg_module/_02131_ ),
    .A2(\reg_module/_02132_ ),
    .B1(\reg_module/_02120_ ),
    .Y(\reg_module/_00872_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19067_  (.A(\reg_module/_09238_ ),
    .B(\reg_module/_02125_ ),
    .Y(\reg_module/_02133_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19068_  (.A(\reg_module/_02127_ ),
    .B(net1752),
    .Y(\reg_module/_02134_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19069_  (.A(\reg_module/_02086_ ),
    .X(\reg_module/_02135_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19070_  (.A1(\reg_module/_02133_ ),
    .A2(\reg_module/_02134_ ),
    .B1(\reg_module/_02135_ ),
    .Y(\reg_module/_00873_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19071_  (.A(\reg_module/_09241_ ),
    .B(\reg_module/_02125_ ),
    .Y(\reg_module/_02136_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19072_  (.A(\reg_module/_02127_ ),
    .B(net1805),
    .Y(\reg_module/_02137_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19073_  (.A1(\reg_module/_02136_ ),
    .A2(\reg_module/_02137_ ),
    .B1(\reg_module/_02135_ ),
    .Y(\reg_module/_00874_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19074_  (.A(\reg_module/_09244_ ),
    .B(\reg_module/_02125_ ),
    .Y(\reg_module/_02138_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19075_  (.A(\reg_module/_02127_ ),
    .B(net1995),
    .Y(\reg_module/_02139_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19076_  (.A1(\reg_module/_02138_ ),
    .A2(\reg_module/_02139_ ),
    .B1(\reg_module/_02135_ ),
    .Y(\reg_module/_00875_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19077_  (.A(\reg_module/_02075_ ),
    .X(\reg_module/_02140_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19078_  (.A(\reg_module/_09250_ ),
    .B(\reg_module/_02140_ ),
    .Y(\reg_module/_02141_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19079_  (.A(\reg_module/_02111_ ),
    .X(\reg_module/_02142_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19080_  (.A(\reg_module/_02142_ ),
    .B(net1823),
    .Y(\reg_module/_02143_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19081_  (.A1(\reg_module/_02141_ ),
    .A2(\reg_module/_02143_ ),
    .B1(\reg_module/_02135_ ),
    .Y(\reg_module/_00876_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19082_  (.A(\reg_module/_09253_ ),
    .B(\reg_module/_02140_ ),
    .Y(\reg_module/_02144_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19083_  (.A(\reg_module/_02142_ ),
    .B(net1873),
    .Y(\reg_module/_02145_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19084_  (.A1(\reg_module/_02144_ ),
    .A2(\reg_module/_02145_ ),
    .B1(\reg_module/_02135_ ),
    .Y(\reg_module/_00877_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19085_  (.A(\reg_module/_09256_ ),
    .B(\reg_module/_02140_ ),
    .Y(\reg_module/_02146_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19086_  (.A(\reg_module/_02142_ ),
    .B(net1976),
    .Y(\reg_module/_02147_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19087_  (.A1(\reg_module/_02146_ ),
    .A2(\reg_module/_02147_ ),
    .B1(\reg_module/_02135_ ),
    .Y(\reg_module/_00878_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19088_  (.A(\reg_module/_09260_ ),
    .B(\reg_module/_02140_ ),
    .Y(\reg_module/_02148_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19089_  (.A(\reg_module/_02142_ ),
    .B(net1762),
    .Y(\reg_module/_02149_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_19090_  (.A(\reg_module/_02086_ ),
    .X(\reg_module/_02150_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19091_  (.A1(\reg_module/_02148_ ),
    .A2(\reg_module/_02149_ ),
    .B1(\reg_module/_02150_ ),
    .Y(\reg_module/_00879_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19092_  (.A(\reg_module/_09263_ ),
    .B(\reg_module/_02140_ ),
    .Y(\reg_module/_02151_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19093_  (.A(\reg_module/_02142_ ),
    .B(net1902),
    .Y(\reg_module/_02152_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19094_  (.A1(\reg_module/_02151_ ),
    .A2(\reg_module/_02152_ ),
    .B1(\reg_module/_02150_ ),
    .Y(\reg_module/_00880_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19095_  (.A(\reg_module/_09266_ ),
    .B(\reg_module/_02140_ ),
    .Y(\reg_module/_02153_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19096_  (.A(\reg_module/_02142_ ),
    .B(net2018),
    .Y(\reg_module/_02154_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19097_  (.A1(\reg_module/_02153_ ),
    .A2(\reg_module/_02154_ ),
    .B1(\reg_module/_02150_ ),
    .Y(\reg_module/_00881_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19098_  (.A(\reg_module/_02075_ ),
    .X(\reg_module/_02155_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19099_  (.A(\reg_module/_09273_ ),
    .B(\reg_module/_02155_ ),
    .Y(\reg_module/_02156_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19100_  (.A(\reg_module/_02111_ ),
    .X(\reg_module/_02157_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19101_  (.A(\reg_module/_02157_ ),
    .B(net1951),
    .Y(\reg_module/_02158_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19102_  (.A1(\reg_module/_02156_ ),
    .A2(\reg_module/_02158_ ),
    .B1(\reg_module/_02150_ ),
    .Y(\reg_module/_00882_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19103_  (.A(\reg_module/_09276_ ),
    .B(\reg_module/_02155_ ),
    .Y(\reg_module/_02159_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19104_  (.A(\reg_module/_02157_ ),
    .B(net1882),
    .Y(\reg_module/_02160_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19105_  (.A1(\reg_module/_02159_ ),
    .A2(\reg_module/_02160_ ),
    .B1(\reg_module/_02150_ ),
    .Y(\reg_module/_00883_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19106_  (.A(\reg_module/_09279_ ),
    .B(\reg_module/_02155_ ),
    .Y(\reg_module/_02161_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19107_  (.A(\reg_module/_02157_ ),
    .B(net2008),
    .Y(\reg_module/_02162_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19108_  (.A1(\reg_module/_02161_ ),
    .A2(\reg_module/_02162_ ),
    .B1(\reg_module/_02150_ ),
    .Y(\reg_module/_00884_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19109_  (.A(\reg_module/_09283_ ),
    .B(\reg_module/_02155_ ),
    .Y(\reg_module/_02163_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19110_  (.A(\reg_module/_02157_ ),
    .B(net1966),
    .Y(\reg_module/_02164_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19111_  (.A(\reg_module/_02086_ ),
    .X(\reg_module/_02165_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19112_  (.A1(\reg_module/_02163_ ),
    .A2(\reg_module/_02164_ ),
    .B1(\reg_module/_02165_ ),
    .Y(\reg_module/_00885_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19113_  (.A(\reg_module/_09286_ ),
    .B(\reg_module/_02155_ ),
    .Y(\reg_module/_02166_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19114_  (.A(\reg_module/_02157_ ),
    .B(net1844),
    .Y(\reg_module/_02167_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19115_  (.A1(\reg_module/_02166_ ),
    .A2(\reg_module/_02167_ ),
    .B1(\reg_module/_02165_ ),
    .Y(\reg_module/_00886_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19116_  (.A(\reg_module/_09289_ ),
    .B(\reg_module/_02155_ ),
    .Y(\reg_module/_02168_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19117_  (.A(\reg_module/_02157_ ),
    .B(net2104),
    .Y(\reg_module/_02169_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19118_  (.A1(\reg_module/_02168_ ),
    .A2(\reg_module/_02169_ ),
    .B1(\reg_module/_02165_ ),
    .Y(\reg_module/_00887_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_19119_  (.A(\reg_module/_01381_ ),
    .X(\reg_module/_02170_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19120_  (.A(\reg_module/_02170_ ),
    .X(\reg_module/_02171_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19121_  (.A(\reg_module/_09295_ ),
    .B(\reg_module/_02171_ ),
    .Y(\reg_module/_02172_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19122_  (.A(\reg_module/_02110_ ),
    .X(\reg_module/_02173_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19123_  (.A(\reg_module/_02173_ ),
    .B(net1619),
    .Y(\reg_module/_02174_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19124_  (.A1(\reg_module/_02172_ ),
    .A2(\reg_module/_02174_ ),
    .B1(\reg_module/_02165_ ),
    .Y(\reg_module/_00888_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19125_  (.A(\reg_module/_09298_ ),
    .B(\reg_module/_02171_ ),
    .Y(\reg_module/_02175_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19126_  (.A(\reg_module/_02173_ ),
    .B(net1393),
    .Y(\reg_module/_02176_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19127_  (.A1(\reg_module/_02175_ ),
    .A2(\reg_module/_02176_ ),
    .B1(\reg_module/_02165_ ),
    .Y(\reg_module/_00889_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19128_  (.A(\reg_module/_09301_ ),
    .B(\reg_module/_02171_ ),
    .Y(\reg_module/_02177_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19129_  (.A(\reg_module/_02173_ ),
    .B(net1862),
    .Y(\reg_module/_02178_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19130_  (.A1(\reg_module/_02177_ ),
    .A2(\reg_module/_02178_ ),
    .B1(\reg_module/_02165_ ),
    .Y(\reg_module/_00890_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19131_  (.A(\reg_module/_09307_ ),
    .B(\reg_module/_02171_ ),
    .Y(\reg_module/_02179_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19132_  (.A(\reg_module/_02173_ ),
    .B(net1547),
    .Y(\reg_module/_02180_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19133_  (.A(\reg_module/_01545_ ),
    .X(\reg_module/_02181_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19134_  (.A(\reg_module/_02181_ ),
    .X(\reg_module/_02182_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19135_  (.A1(\reg_module/_02179_ ),
    .A2(\reg_module/_02180_ ),
    .B1(\reg_module/_02182_ ),
    .Y(\reg_module/_00891_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19136_  (.A(\reg_module/_09310_ ),
    .B(\reg_module/_02171_ ),
    .Y(\reg_module/_02183_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19137_  (.A(\reg_module/_02173_ ),
    .B(net1571),
    .Y(\reg_module/_02184_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19138_  (.A1(\reg_module/_02183_ ),
    .A2(\reg_module/_02184_ ),
    .B1(\reg_module/_02182_ ),
    .Y(\reg_module/_00892_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19139_  (.A(\reg_module/_09313_ ),
    .B(\reg_module/_02171_ ),
    .Y(\reg_module/_02185_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19140_  (.A(\reg_module/_02173_ ),
    .B(net1482),
    .Y(\reg_module/_02186_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19141_  (.A1(\reg_module/_02185_ ),
    .A2(\reg_module/_02186_ ),
    .B1(\reg_module/_02182_ ),
    .Y(\reg_module/_00893_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_19142_  (.A(\reg_module/_02170_ ),
    .X(\reg_module/_02187_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19143_  (.A(\reg_module/_09317_ ),
    .B(\reg_module/_02187_ ),
    .Y(\reg_module/_02188_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19144_  (.A(\reg_module/_02111_ ),
    .B(net1531),
    .Y(\reg_module/_02189_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19145_  (.A1(\reg_module/_02188_ ),
    .A2(\reg_module/_02189_ ),
    .B1(\reg_module/_02182_ ),
    .Y(\reg_module/_00894_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19146_  (.A(\reg_module/_09320_ ),
    .B(\reg_module/_02187_ ),
    .Y(\reg_module/_02190_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19147_  (.A(\reg_module/_02111_ ),
    .B(net1697),
    .Y(\reg_module/_02191_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19148_  (.A1(\reg_module/_02190_ ),
    .A2(\reg_module/_02191_ ),
    .B1(\reg_module/_02182_ ),
    .Y(\reg_module/_00895_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_19149_  (.A(\reg_module/_07653_ ),
    .X(\reg_module/_02192_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_19150_  (.A(\reg_module/_02192_ ),
    .X(\reg_module/_02193_ ));
 sky130_fd_sc_hd__nor2_2 \reg_module/_19151_  (.A(\reg_module/_09322_ ),
    .B(\reg_module/_01154_ ),
    .Y(\reg_module/_02194_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_19152_  (.A(\reg_module/_02194_ ),
    .X(\reg_module/_02195_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19153_  (.A(\reg_module/_02195_ ),
    .X(\reg_module/_02196_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19154_  (.A(\reg_module/gprf[896] ),
    .B(\reg_module/_02196_ ),
    .Y(\reg_module/_02197_ ));
 sky130_fd_sc_hd__clkbuf_8 \reg_module/_19155_  (.A(\reg_module/_07635_ ),
    .X(\reg_module/_02198_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19156_  (.A(\reg_module/_02198_ ),
    .X(\reg_module/_02199_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19157_  (.A(\reg_module/_02194_ ),
    .X(\reg_module/_02200_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19158_  (.A1(\reg_module/_07513_ ),
    .A2(\reg_module/_02199_ ),
    .B1(\reg_module/_02200_ ),
    .Y(\reg_module/_02201_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19159_  (.A(\reg_module/_02193_ ),
    .B(\reg_module/_02197_ ),
    .C_N(\reg_module/_02201_ ),
    .Y(\reg_module/_00896_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19160_  (.A(\reg_module/gprf[897] ),
    .B(\reg_module/_02196_ ),
    .Y(\reg_module/_02202_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19161_  (.A1(\reg_module/_07517_ ),
    .A2(\reg_module/_02199_ ),
    .B1(\reg_module/_02200_ ),
    .Y(\reg_module/_02203_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19162_  (.A(\reg_module/_02193_ ),
    .B(\reg_module/_02202_ ),
    .C_N(\reg_module/_02203_ ),
    .Y(\reg_module/_00897_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19163_  (.A(\reg_module/gprf[898] ),
    .B(\reg_module/_02196_ ),
    .Y(\reg_module/_02204_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19164_  (.A1(\reg_module/_07520_ ),
    .A2(\reg_module/_02199_ ),
    .B1(\reg_module/_02200_ ),
    .Y(\reg_module/_02205_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19165_  (.A(\reg_module/_02193_ ),
    .B(\reg_module/_02204_ ),
    .C_N(\reg_module/_02205_ ),
    .Y(\reg_module/_00898_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19166_  (.A(\reg_module/_07654_ ),
    .X(\reg_module/_02206_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19167_  (.A(\reg_module/gprf[899] ),
    .B(\reg_module/_02196_ ),
    .Y(\reg_module/_02207_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19168_  (.A1(\reg_module/_07522_ ),
    .A2(\reg_module/_02199_ ),
    .B1(\reg_module/_02200_ ),
    .Y(\reg_module/_02208_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19169_  (.A(\reg_module/_02206_ ),
    .B(\reg_module/_02207_ ),
    .C_N(\reg_module/_02208_ ),
    .Y(\reg_module/_00899_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19170_  (.A(\reg_module/gprf[900] ),
    .B(\reg_module/_02196_ ),
    .Y(\reg_module/_02209_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_19171_  (.A(\reg_module/_02194_ ),
    .X(\reg_module/_02210_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19172_  (.A(\reg_module/_02210_ ),
    .X(\reg_module/_02211_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19173_  (.A1(\reg_module/_07527_ ),
    .A2(\reg_module/_02199_ ),
    .B1(\reg_module/_02211_ ),
    .Y(\reg_module/_02212_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19174_  (.A(\reg_module/_02206_ ),
    .B(\reg_module/_02209_ ),
    .C_N(\reg_module/_02212_ ),
    .Y(\reg_module/_00900_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19175_  (.A(\reg_module/gprf[901] ),
    .B(\reg_module/_02196_ ),
    .Y(\reg_module/_02213_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19176_  (.A1(\reg_module/_07531_ ),
    .A2(\reg_module/_02199_ ),
    .B1(\reg_module/_02211_ ),
    .Y(\reg_module/_02214_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19177_  (.A(\reg_module/_02206_ ),
    .B(\reg_module/_02213_ ),
    .C_N(\reg_module/_02214_ ),
    .Y(\reg_module/_00901_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19178_  (.A(\reg_module/_02195_ ),
    .X(\reg_module/_02215_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19179_  (.A(net2103),
    .B(\reg_module/_02215_ ),
    .Y(\reg_module/_02216_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19180_  (.A(\reg_module/_02198_ ),
    .X(\reg_module/_02217_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19181_  (.A1(\reg_module/_07534_ ),
    .A2(\reg_module/_02217_ ),
    .B1(\reg_module/_02211_ ),
    .Y(\reg_module/_02218_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19182_  (.A(\reg_module/_02206_ ),
    .B(\reg_module/_02216_ ),
    .C_N(\reg_module/_02218_ ),
    .Y(\reg_module/_00902_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19183_  (.A(net2116),
    .B(\reg_module/_02215_ ),
    .Y(\reg_module/_02219_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19184_  (.A1(\reg_module/_07538_ ),
    .A2(\reg_module/_02217_ ),
    .B1(\reg_module/_02211_ ),
    .Y(\reg_module/_02220_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19185_  (.A(\reg_module/_02206_ ),
    .B(\reg_module/_02219_ ),
    .C_N(\reg_module/_02220_ ),
    .Y(\reg_module/_00903_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19186_  (.A(net2062),
    .B(\reg_module/_02215_ ),
    .Y(\reg_module/_02221_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19187_  (.A1(\reg_module/_07540_ ),
    .A2(\reg_module/_02217_ ),
    .B1(\reg_module/_02211_ ),
    .Y(\reg_module/_02222_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19188_  (.A(\reg_module/_02206_ ),
    .B(\reg_module/_02221_ ),
    .C_N(\reg_module/_02222_ ),
    .Y(\reg_module/_00904_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19189_  (.A(\reg_module/_07654_ ),
    .X(\reg_module/_02223_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19190_  (.A(net2101),
    .B(\reg_module/_02215_ ),
    .Y(\reg_module/_02224_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19191_  (.A1(\reg_module/_07544_ ),
    .A2(\reg_module/_02217_ ),
    .B1(\reg_module/_02211_ ),
    .Y(\reg_module/_02225_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19192_  (.A(\reg_module/_02223_ ),
    .B(\reg_module/_02224_ ),
    .C_N(\reg_module/_02225_ ),
    .Y(\reg_module/_00905_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19193_  (.A(net2111),
    .B(\reg_module/_02215_ ),
    .Y(\reg_module/_02226_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19194_  (.A(\reg_module/_02210_ ),
    .X(\reg_module/_02227_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19195_  (.A1(\reg_module/_07547_ ),
    .A2(\reg_module/_02217_ ),
    .B1(\reg_module/_02227_ ),
    .Y(\reg_module/_02228_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19196_  (.A(\reg_module/_02223_ ),
    .B(\reg_module/_02226_ ),
    .C_N(\reg_module/_02228_ ),
    .Y(\reg_module/_00906_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19197_  (.A(net2084),
    .B(\reg_module/_02215_ ),
    .Y(\reg_module/_02229_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19198_  (.A1(\reg_module/_07551_ ),
    .A2(\reg_module/_02217_ ),
    .B1(\reg_module/_02227_ ),
    .Y(\reg_module/_02230_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19199_  (.A(\reg_module/_02223_ ),
    .B(\reg_module/_02229_ ),
    .C_N(\reg_module/_02230_ ),
    .Y(\reg_module/_00907_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19200_  (.A(\reg_module/_02210_ ),
    .X(\reg_module/_02231_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19201_  (.A(\reg_module/gprf[908] ),
    .B(\reg_module/_02231_ ),
    .Y(\reg_module/_02232_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19202_  (.A(\reg_module/_02198_ ),
    .X(\reg_module/_02233_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19203_  (.A1(\reg_module/_07554_ ),
    .A2(\reg_module/_02233_ ),
    .B1(\reg_module/_02227_ ),
    .Y(\reg_module/_02234_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19204_  (.A(\reg_module/_02223_ ),
    .B(\reg_module/_02232_ ),
    .C_N(\reg_module/_02234_ ),
    .Y(\reg_module/_00908_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19205_  (.A(net2208),
    .B(\reg_module/_02231_ ),
    .Y(\reg_module/_02235_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19206_  (.A1(\reg_module/_07557_ ),
    .A2(\reg_module/_02233_ ),
    .B1(\reg_module/_02227_ ),
    .Y(\reg_module/_02236_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19207_  (.A(\reg_module/_02223_ ),
    .B(\reg_module/_02235_ ),
    .C_N(\reg_module/_02236_ ),
    .Y(\reg_module/_00909_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19208_  (.A(net2195),
    .B(\reg_module/_02231_ ),
    .Y(\reg_module/_02237_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19209_  (.A1(\reg_module/_07560_ ),
    .A2(\reg_module/_02233_ ),
    .B1(\reg_module/_02227_ ),
    .Y(\reg_module/_02238_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19210_  (.A(\reg_module/_02223_ ),
    .B(\reg_module/_02237_ ),
    .C_N(\reg_module/_02238_ ),
    .Y(\reg_module/_00910_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19211_  (.A(\reg_module/_07654_ ),
    .X(\reg_module/_02239_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19212_  (.A(net2198),
    .B(\reg_module/_02231_ ),
    .Y(\reg_module/_02240_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19213_  (.A1(\reg_module/_07564_ ),
    .A2(\reg_module/_02233_ ),
    .B1(\reg_module/_02227_ ),
    .Y(\reg_module/_02241_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19214_  (.A(\reg_module/_02239_ ),
    .B(\reg_module/_02240_ ),
    .C_N(\reg_module/_02241_ ),
    .Y(\reg_module/_00911_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19215_  (.A(net2163),
    .B(\reg_module/_02231_ ),
    .Y(\reg_module/_02242_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19216_  (.A(\reg_module/_02210_ ),
    .X(\reg_module/_02243_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19217_  (.A1(\reg_module/_07567_ ),
    .A2(\reg_module/_02233_ ),
    .B1(\reg_module/_02243_ ),
    .Y(\reg_module/_02244_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19218_  (.A(\reg_module/_02239_ ),
    .B(\reg_module/_02242_ ),
    .C_N(\reg_module/_02244_ ),
    .Y(\reg_module/_00912_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19219_  (.A(net2093),
    .B(\reg_module/_02231_ ),
    .Y(\reg_module/_02245_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19220_  (.A1(\reg_module/_07571_ ),
    .A2(\reg_module/_02233_ ),
    .B1(\reg_module/_02243_ ),
    .Y(\reg_module/_02246_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19221_  (.A(\reg_module/_02239_ ),
    .B(\reg_module/_02245_ ),
    .C_N(\reg_module/_02246_ ),
    .Y(\reg_module/_00913_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19222_  (.A(\reg_module/_02210_ ),
    .X(\reg_module/_02247_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19223_  (.A(net2145),
    .B(\reg_module/_02247_ ),
    .Y(\reg_module/_02248_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19224_  (.A(\reg_module/_02198_ ),
    .X(\reg_module/_02249_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19225_  (.A1(\reg_module/_07574_ ),
    .A2(\reg_module/_02249_ ),
    .B1(\reg_module/_02243_ ),
    .Y(\reg_module/_02250_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19226_  (.A(\reg_module/_02239_ ),
    .B(\reg_module/_02248_ ),
    .C_N(\reg_module/_02250_ ),
    .Y(\reg_module/_00914_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19227_  (.A(net2085),
    .B(\reg_module/_02247_ ),
    .Y(\reg_module/_02251_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19228_  (.A1(\reg_module/_07578_ ),
    .A2(\reg_module/_02249_ ),
    .B1(\reg_module/_02243_ ),
    .Y(\reg_module/_02252_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19229_  (.A(\reg_module/_02239_ ),
    .B(\reg_module/_02251_ ),
    .C_N(\reg_module/_02252_ ),
    .Y(\reg_module/_00915_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19230_  (.A(net2082),
    .B(\reg_module/_02247_ ),
    .Y(\reg_module/_02253_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19231_  (.A1(\reg_module/_07580_ ),
    .A2(\reg_module/_02249_ ),
    .B1(\reg_module/_02243_ ),
    .Y(\reg_module/_02254_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19232_  (.A(\reg_module/_02239_ ),
    .B(\reg_module/_02253_ ),
    .C_N(\reg_module/_02254_ ),
    .Y(\reg_module/_00916_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_19233_  (.A(\reg_module/_07654_ ),
    .X(\reg_module/_02255_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19234_  (.A(net2060),
    .B(\reg_module/_02247_ ),
    .Y(\reg_module/_02256_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19235_  (.A1(\reg_module/_07584_ ),
    .A2(\reg_module/_02249_ ),
    .B1(\reg_module/_02243_ ),
    .Y(\reg_module/_02257_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19236_  (.A(\reg_module/_02255_ ),
    .B(\reg_module/_02256_ ),
    .C_N(\reg_module/_02257_ ),
    .Y(\reg_module/_00917_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19237_  (.A(net2068),
    .B(\reg_module/_02247_ ),
    .Y(\reg_module/_02258_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19238_  (.A(\reg_module/_02194_ ),
    .X(\reg_module/_02259_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19239_  (.A1(\reg_module/_07587_ ),
    .A2(\reg_module/_02249_ ),
    .B1(\reg_module/_02259_ ),
    .Y(\reg_module/_02260_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19240_  (.A(\reg_module/_02255_ ),
    .B(\reg_module/_02258_ ),
    .C_N(\reg_module/_02260_ ),
    .Y(\reg_module/_00918_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19241_  (.A(net2125),
    .B(\reg_module/_02247_ ),
    .Y(\reg_module/_02261_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19242_  (.A1(\reg_module/_07590_ ),
    .A2(\reg_module/_02249_ ),
    .B1(\reg_module/_02259_ ),
    .Y(\reg_module/_02262_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19243_  (.A(\reg_module/_02255_ ),
    .B(\reg_module/_02261_ ),
    .C_N(\reg_module/_02262_ ),
    .Y(\reg_module/_00919_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19244_  (.A(\reg_module/_02210_ ),
    .X(\reg_module/_02263_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19245_  (.A(net2071),
    .B(\reg_module/_02263_ ),
    .Y(\reg_module/_02264_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19246_  (.A(\reg_module/_07635_ ),
    .X(\reg_module/_02265_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19247_  (.A1(\reg_module/_07594_ ),
    .A2(\reg_module/_02265_ ),
    .B1(\reg_module/_02259_ ),
    .Y(\reg_module/_02266_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19248_  (.A(\reg_module/_02255_ ),
    .B(\reg_module/_02264_ ),
    .C_N(\reg_module/_02266_ ),
    .Y(\reg_module/_00920_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19249_  (.A(net2049),
    .B(\reg_module/_02263_ ),
    .Y(\reg_module/_02267_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19250_  (.A1(\reg_module/_07598_ ),
    .A2(\reg_module/_02265_ ),
    .B1(\reg_module/_02259_ ),
    .Y(\reg_module/_02268_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19251_  (.A(\reg_module/_02255_ ),
    .B(\reg_module/_02267_ ),
    .C_N(\reg_module/_02268_ ),
    .Y(\reg_module/_00921_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19252_  (.A(net2136),
    .B(\reg_module/_02263_ ),
    .Y(\reg_module/_02269_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19253_  (.A1(\reg_module/_07601_ ),
    .A2(\reg_module/_02265_ ),
    .B1(\reg_module/_02259_ ),
    .Y(\reg_module/_02270_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19254_  (.A(\reg_module/_02255_ ),
    .B(\reg_module/_02269_ ),
    .C_N(\reg_module/_02270_ ),
    .Y(\reg_module/_00922_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19255_  (.A(net2090),
    .B(\reg_module/_02263_ ),
    .Y(\reg_module/_02271_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19256_  (.A1(\reg_module/_07604_ ),
    .A2(\reg_module/_02265_ ),
    .B1(\reg_module/_02259_ ),
    .Y(\reg_module/_02272_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19257_  (.A(\reg_module/_01546_ ),
    .B(\reg_module/_02271_ ),
    .C_N(\reg_module/_02272_ ),
    .Y(\reg_module/_00923_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19258_  (.A(net2122),
    .B(\reg_module/_02263_ ),
    .Y(\reg_module/_02273_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19259_  (.A1(\reg_module/_07606_ ),
    .A2(\reg_module/_02265_ ),
    .B1(\reg_module/_02195_ ),
    .Y(\reg_module/_02274_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19260_  (.A(\reg_module/_01546_ ),
    .B(\reg_module/_02273_ ),
    .C_N(\reg_module/_02274_ ),
    .Y(\reg_module/_00924_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19261_  (.A(net2137),
    .B(\reg_module/_02263_ ),
    .Y(\reg_module/_02275_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19262_  (.A1(\reg_module/_07610_ ),
    .A2(\reg_module/_02265_ ),
    .B1(\reg_module/_02195_ ),
    .Y(\reg_module/_02276_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19263_  (.A(\reg_module/_01546_ ),
    .B(\reg_module/_02275_ ),
    .C_N(\reg_module/_02276_ ),
    .Y(\reg_module/_00925_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19264_  (.A(net2126),
    .B(\reg_module/_02200_ ),
    .Y(\reg_module/_02277_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19265_  (.A1(\reg_module/_07612_ ),
    .A2(\reg_module/_02198_ ),
    .B1(\reg_module/_02195_ ),
    .Y(\reg_module/_02278_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19266_  (.A(\reg_module/_01546_ ),
    .B(\reg_module/_02277_ ),
    .C_N(\reg_module/_02278_ ),
    .Y(\reg_module/_00926_ ));
 sky130_fd_sc_hd__nor2_1 \reg_module/_19267_  (.A(net2077),
    .B(\reg_module/_02200_ ),
    .Y(\reg_module/_02279_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19268_  (.A1(\reg_module/_07616_ ),
    .A2(\reg_module/_02198_ ),
    .B1(\reg_module/_02195_ ),
    .Y(\reg_module/_02280_ ));
 sky130_fd_sc_hd__nor3b_1 \reg_module/_19269_  (.A(\reg_module/_01546_ ),
    .B(\reg_module/_02279_ ),
    .C_N(\reg_module/_02280_ ),
    .Y(\reg_module/_00927_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19270_  (.A(\reg_module/_09507_ ),
    .B(\reg_module/_02187_ ),
    .Y(\reg_module/_02281_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19271_  (.A(\reg_module/_01155_ ),
    .X(\reg_module/_02282_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19272_  (.A(\reg_module/_08366_ ),
    .B(\reg_module/_07626_ ),
    .Y(\reg_module/_02283_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_19273_  (.A(\reg_module/_02283_ ),
    .X(\reg_module/_02284_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19274_  (.A(\reg_module/_02284_ ),
    .X(\reg_module/_02285_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19275_  (.A1(\reg_module/_02282_ ),
    .A2(\reg_module/_02285_ ),
    .B1(net1818),
    .Y(\reg_module/_02286_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19276_  (.A1(\reg_module/_02281_ ),
    .A2(\reg_module/_02286_ ),
    .B1(\reg_module/_02182_ ),
    .Y(\reg_module/_00928_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19277_  (.A(\reg_module/_09512_ ),
    .B(\reg_module/_02187_ ),
    .Y(\reg_module/_02287_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19278_  (.A1(\reg_module/_02282_ ),
    .A2(\reg_module/_02285_ ),
    .B1(net1935),
    .Y(\reg_module/_02288_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19279_  (.A(\reg_module/_02181_ ),
    .X(\reg_module/_02289_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19280_  (.A1(\reg_module/_02287_ ),
    .A2(\reg_module/_02288_ ),
    .B1(\reg_module/_02289_ ),
    .Y(\reg_module/_00929_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19281_  (.A(\reg_module/_09516_ ),
    .B(\reg_module/_02187_ ),
    .Y(\reg_module/_02290_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19282_  (.A1(\reg_module/_02282_ ),
    .A2(\reg_module/_02285_ ),
    .B1(net1662),
    .Y(\reg_module/_02291_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19283_  (.A1(\reg_module/_02290_ ),
    .A2(\reg_module/_02291_ ),
    .B1(\reg_module/_02289_ ),
    .Y(\reg_module/_00930_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19284_  (.A(\reg_module/_09519_ ),
    .B(\reg_module/_02187_ ),
    .Y(\reg_module/_02292_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19285_  (.A1(\reg_module/_02282_ ),
    .A2(\reg_module/_02285_ ),
    .B1(net1865),
    .Y(\reg_module/_02293_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19286_  (.A1(\reg_module/_02292_ ),
    .A2(\reg_module/_02293_ ),
    .B1(\reg_module/_02289_ ),
    .Y(\reg_module/_00931_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19287_  (.A(\reg_module/_02170_ ),
    .X(\reg_module/_02294_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19288_  (.A(\reg_module/_09522_ ),
    .B(\reg_module/_02294_ ),
    .Y(\reg_module/_02295_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19289_  (.A1(\reg_module/_02282_ ),
    .A2(\reg_module/_02285_ ),
    .B1(net2025),
    .Y(\reg_module/_02296_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19290_  (.A1(\reg_module/_02295_ ),
    .A2(\reg_module/_02296_ ),
    .B1(\reg_module/_02289_ ),
    .Y(\reg_module/_00932_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19291_  (.A(\reg_module/_09525_ ),
    .B(\reg_module/_02294_ ),
    .Y(\reg_module/_02297_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19292_  (.A1(\reg_module/_02282_ ),
    .A2(\reg_module/_02285_ ),
    .B1(net2010),
    .Y(\reg_module/_02298_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19293_  (.A1(\reg_module/_02297_ ),
    .A2(\reg_module/_02298_ ),
    .B1(\reg_module/_02289_ ),
    .Y(\reg_module/_00933_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19294_  (.A(\reg_module/_09529_ ),
    .B(\reg_module/_02294_ ),
    .Y(\reg_module/_02299_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19295_  (.A(\reg_module/_01155_ ),
    .X(\reg_module/_02300_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19296_  (.A(\reg_module/_02284_ ),
    .X(\reg_module/_02301_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19297_  (.A1(\reg_module/_02300_ ),
    .A2(\reg_module/_02301_ ),
    .B1(net2148),
    .Y(\reg_module/_02302_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19298_  (.A1(\reg_module/_02299_ ),
    .A2(\reg_module/_02302_ ),
    .B1(\reg_module/_02289_ ),
    .Y(\reg_module/_00934_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19299_  (.A(\reg_module/_09534_ ),
    .B(\reg_module/_02294_ ),
    .Y(\reg_module/_02303_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19300_  (.A1(\reg_module/_02300_ ),
    .A2(\reg_module/_02301_ ),
    .B1(net2080),
    .Y(\reg_module/_02304_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19301_  (.A(\reg_module/_02181_ ),
    .X(\reg_module/_02305_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19302_  (.A1(\reg_module/_02303_ ),
    .A2(\reg_module/_02304_ ),
    .B1(\reg_module/_02305_ ),
    .Y(\reg_module/_00935_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19303_  (.A(\reg_module/_09538_ ),
    .B(\reg_module/_02294_ ),
    .Y(\reg_module/_02306_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19304_  (.A1(\reg_module/_02300_ ),
    .A2(\reg_module/_02301_ ),
    .B1(net2123),
    .Y(\reg_module/_02307_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19305_  (.A1(\reg_module/_02306_ ),
    .A2(\reg_module/_02307_ ),
    .B1(\reg_module/_02305_ ),
    .Y(\reg_module/_00936_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19306_  (.A(\reg_module/_09541_ ),
    .B(\reg_module/_02294_ ),
    .Y(\reg_module/_02308_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19307_  (.A1(\reg_module/_02300_ ),
    .A2(\reg_module/_02301_ ),
    .B1(net2051),
    .Y(\reg_module/_02309_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19308_  (.A1(\reg_module/_02308_ ),
    .A2(\reg_module/_02309_ ),
    .B1(\reg_module/_02305_ ),
    .Y(\reg_module/_00937_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19309_  (.A(\reg_module/_02170_ ),
    .X(\reg_module/_02310_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19310_  (.A(\reg_module/_09544_ ),
    .B(\reg_module/_02310_ ),
    .Y(\reg_module/_02311_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19311_  (.A1(\reg_module/_02300_ ),
    .A2(\reg_module/_02301_ ),
    .B1(net2024),
    .Y(\reg_module/_02312_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19312_  (.A1(\reg_module/_02311_ ),
    .A2(\reg_module/_02312_ ),
    .B1(\reg_module/_02305_ ),
    .Y(\reg_module/_00938_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19313_  (.A(\reg_module/_09547_ ),
    .B(\reg_module/_02310_ ),
    .Y(\reg_module/_02313_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19314_  (.A1(\reg_module/_02300_ ),
    .A2(\reg_module/_02301_ ),
    .B1(net2038),
    .Y(\reg_module/_02314_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19315_  (.A1(\reg_module/_02313_ ),
    .A2(\reg_module/_02314_ ),
    .B1(\reg_module/_02305_ ),
    .Y(\reg_module/_00939_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19316_  (.A(\reg_module/_09551_ ),
    .B(\reg_module/_02310_ ),
    .Y(\reg_module/_02315_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19317_  (.A(\reg_module/_01155_ ),
    .X(\reg_module/_02316_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19318_  (.A(\reg_module/_02284_ ),
    .X(\reg_module/_02317_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19319_  (.A1(\reg_module/_02316_ ),
    .A2(\reg_module/_02317_ ),
    .B1(net2108),
    .Y(\reg_module/_02318_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19320_  (.A1(\reg_module/_02315_ ),
    .A2(\reg_module/_02318_ ),
    .B1(\reg_module/_02305_ ),
    .Y(\reg_module/_00940_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19321_  (.A(\reg_module/_09556_ ),
    .B(\reg_module/_02310_ ),
    .Y(\reg_module/_02319_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19322_  (.A1(\reg_module/_02316_ ),
    .A2(\reg_module/_02317_ ),
    .B1(net1993),
    .Y(\reg_module/_02320_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19323_  (.A(\reg_module/_02181_ ),
    .X(\reg_module/_02321_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19324_  (.A1(\reg_module/_02319_ ),
    .A2(\reg_module/_02320_ ),
    .B1(\reg_module/_02321_ ),
    .Y(\reg_module/_00941_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19325_  (.A(\reg_module/_09560_ ),
    .B(\reg_module/_02310_ ),
    .Y(\reg_module/_02322_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19326_  (.A1(\reg_module/_02316_ ),
    .A2(\reg_module/_02317_ ),
    .B1(net2032),
    .Y(\reg_module/_02323_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19327_  (.A1(\reg_module/_02322_ ),
    .A2(\reg_module/_02323_ ),
    .B1(\reg_module/_02321_ ),
    .Y(\reg_module/_00942_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19328_  (.A(\reg_module/_09563_ ),
    .B(\reg_module/_02310_ ),
    .Y(\reg_module/_02324_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19329_  (.A1(\reg_module/_02316_ ),
    .A2(\reg_module/_02317_ ),
    .B1(net2028),
    .Y(\reg_module/_02325_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19330_  (.A1(\reg_module/_02324_ ),
    .A2(\reg_module/_02325_ ),
    .B1(\reg_module/_02321_ ),
    .Y(\reg_module/_00943_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19331_  (.A(\reg_module/_02170_ ),
    .X(\reg_module/_02326_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19332_  (.A(\reg_module/_09566_ ),
    .B(\reg_module/_02326_ ),
    .Y(\reg_module/_02327_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19333_  (.A1(\reg_module/_02316_ ),
    .A2(\reg_module/_02317_ ),
    .B1(net1927),
    .Y(\reg_module/_02328_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19334_  (.A1(\reg_module/_02327_ ),
    .A2(\reg_module/_02328_ ),
    .B1(\reg_module/_02321_ ),
    .Y(\reg_module/_00944_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19335_  (.A(\reg_module/_09569_ ),
    .B(\reg_module/_02326_ ),
    .Y(\reg_module/_02329_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19336_  (.A1(\reg_module/_02316_ ),
    .A2(\reg_module/_02317_ ),
    .B1(net2139),
    .Y(\reg_module/_02330_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19337_  (.A1(\reg_module/_02329_ ),
    .A2(\reg_module/_02330_ ),
    .B1(\reg_module/_02321_ ),
    .Y(\reg_module/_00945_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19338_  (.A(\reg_module/_09573_ ),
    .B(\reg_module/_02326_ ),
    .Y(\reg_module/_02331_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19339_  (.A(\reg_module/_01155_ ),
    .X(\reg_module/_02332_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19340_  (.A(\reg_module/_02284_ ),
    .X(\reg_module/_02333_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19341_  (.A1(\reg_module/_02332_ ),
    .A2(\reg_module/_02333_ ),
    .B1(net1803),
    .Y(\reg_module/_02334_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19342_  (.A1(\reg_module/_02331_ ),
    .A2(\reg_module/_02334_ ),
    .B1(\reg_module/_02321_ ),
    .Y(\reg_module/_00946_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19343_  (.A(\reg_module/_09578_ ),
    .B(\reg_module/_02326_ ),
    .Y(\reg_module/_02335_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19344_  (.A1(\reg_module/_02332_ ),
    .A2(\reg_module/_02333_ ),
    .B1(net1644),
    .Y(\reg_module/_02336_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19345_  (.A(\reg_module/_02181_ ),
    .X(\reg_module/_02337_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19346_  (.A1(\reg_module/_02335_ ),
    .A2(\reg_module/_02336_ ),
    .B1(\reg_module/_02337_ ),
    .Y(\reg_module/_00947_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19347_  (.A(\reg_module/_09582_ ),
    .B(\reg_module/_02326_ ),
    .Y(\reg_module/_02338_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19348_  (.A1(\reg_module/_02332_ ),
    .A2(\reg_module/_02333_ ),
    .B1(net1881),
    .Y(\reg_module/_02339_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19349_  (.A1(\reg_module/_02338_ ),
    .A2(\reg_module/_02339_ ),
    .B1(\reg_module/_02337_ ),
    .Y(\reg_module/_00948_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19350_  (.A(\reg_module/_09585_ ),
    .B(\reg_module/_02326_ ),
    .Y(\reg_module/_02340_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19351_  (.A1(\reg_module/_02332_ ),
    .A2(\reg_module/_02333_ ),
    .B1(net1765),
    .Y(\reg_module/_02341_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19352_  (.A1(\reg_module/_02340_ ),
    .A2(\reg_module/_02341_ ),
    .B1(\reg_module/_02337_ ),
    .Y(\reg_module/_00949_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19353_  (.A(\reg_module/_02170_ ),
    .X(\reg_module/_02342_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19354_  (.A(\reg_module/_09588_ ),
    .B(\reg_module/_02342_ ),
    .Y(\reg_module/_02343_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19355_  (.A1(\reg_module/_02332_ ),
    .A2(\reg_module/_02333_ ),
    .B1(net1949),
    .Y(\reg_module/_02344_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19356_  (.A1(\reg_module/_02343_ ),
    .A2(\reg_module/_02344_ ),
    .B1(\reg_module/_02337_ ),
    .Y(\reg_module/_00950_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19357_  (.A(\reg_module/_09591_ ),
    .B(\reg_module/_02342_ ),
    .Y(\reg_module/_02345_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19358_  (.A1(\reg_module/_02332_ ),
    .A2(\reg_module/_02333_ ),
    .B1(net2074),
    .Y(\reg_module/_02346_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19359_  (.A1(\reg_module/_02345_ ),
    .A2(\reg_module/_02346_ ),
    .B1(\reg_module/_02337_ ),
    .Y(\reg_module/_00951_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19360_  (.A(\reg_module/_09595_ ),
    .B(\reg_module/_02342_ ),
    .Y(\reg_module/_02347_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19361_  (.A(\reg_module/_01155_ ),
    .X(\reg_module/_02348_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19362_  (.A(\reg_module/_02283_ ),
    .X(\reg_module/_02349_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19363_  (.A1(\reg_module/_02348_ ),
    .A2(\reg_module/_02349_ ),
    .B1(net1984),
    .Y(\reg_module/_02350_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19364_  (.A1(\reg_module/_02347_ ),
    .A2(\reg_module/_02350_ ),
    .B1(\reg_module/_02337_ ),
    .Y(\reg_module/_00952_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19365_  (.A(\reg_module/_09600_ ),
    .B(\reg_module/_02342_ ),
    .Y(\reg_module/_02351_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19366_  (.A1(\reg_module/_02348_ ),
    .A2(\reg_module/_02349_ ),
    .B1(net1867),
    .Y(\reg_module/_02352_ ));
 sky130_fd_sc_hd__clkbuf_4 \reg_module/_19367_  (.A(\reg_module/_02181_ ),
    .X(\reg_module/_02353_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19368_  (.A1(\reg_module/_02351_ ),
    .A2(\reg_module/_02352_ ),
    .B1(\reg_module/_02353_ ),
    .Y(\reg_module/_00953_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19369_  (.A(\reg_module/_09604_ ),
    .B(\reg_module/_02342_ ),
    .Y(\reg_module/_02354_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19370_  (.A1(\reg_module/_02348_ ),
    .A2(\reg_module/_02349_ ),
    .B1(net2079),
    .Y(\reg_module/_02355_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19371_  (.A1(\reg_module/_02354_ ),
    .A2(\reg_module/_02355_ ),
    .B1(\reg_module/_02353_ ),
    .Y(\reg_module/_00954_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19372_  (.A(\reg_module/_09607_ ),
    .B(\reg_module/_02342_ ),
    .Y(\reg_module/_02356_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19373_  (.A1(\reg_module/_02348_ ),
    .A2(\reg_module/_02349_ ),
    .B1(net1945),
    .Y(\reg_module/_02357_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19374_  (.A1(\reg_module/_02356_ ),
    .A2(\reg_module/_02357_ ),
    .B1(\reg_module/_02353_ ),
    .Y(\reg_module/_00955_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19375_  (.A(\reg_module/_09610_ ),
    .B(\reg_module/_01382_ ),
    .Y(\reg_module/_02358_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19376_  (.A1(\reg_module/_02348_ ),
    .A2(\reg_module/_02349_ ),
    .B1(net1819),
    .Y(\reg_module/_02359_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19377_  (.A1(\reg_module/_02358_ ),
    .A2(\reg_module/_02359_ ),
    .B1(\reg_module/_02353_ ),
    .Y(\reg_module/_00956_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19378_  (.A(\reg_module/_09613_ ),
    .B(\reg_module/_01382_ ),
    .Y(\reg_module/_02360_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19379_  (.A1(\reg_module/_02348_ ),
    .A2(\reg_module/_02349_ ),
    .B1(net2052),
    .Y(\reg_module/_02361_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19380_  (.A1(\reg_module/_02360_ ),
    .A2(\reg_module/_02361_ ),
    .B1(\reg_module/_02353_ ),
    .Y(\reg_module/_00957_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19381_  (.A(\reg_module/_09616_ ),
    .B(\reg_module/_01382_ ),
    .Y(\reg_module/_02362_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19382_  (.A1(\reg_module/_01156_ ),
    .A2(\reg_module/_02284_ ),
    .B1(net2035),
    .Y(\reg_module/_02363_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19383_  (.A1(\reg_module/_02362_ ),
    .A2(\reg_module/_02363_ ),
    .B1(\reg_module/_02353_ ),
    .Y(\reg_module/_00958_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19384_  (.A(\reg_module/_09621_ ),
    .B(\reg_module/_01382_ ),
    .Y(\reg_module/_02364_ ));
 sky130_fd_sc_hd__o21ai_1 \reg_module/_19385_  (.A1(\reg_module/_01156_ ),
    .A2(\reg_module/_02284_ ),
    .B1(net2012),
    .Y(\reg_module/_02365_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19386_  (.A(\reg_module/_02192_ ),
    .X(\reg_module/_02366_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19387_  (.A1(\reg_module/_02364_ ),
    .A2(\reg_module/_02365_ ),
    .B1(\reg_module/_02366_ ),
    .Y(\reg_module/_00959_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19388_  (.A(\reg_module/_01300_ ),
    .B(\reg_module/_09623_ ),
    .Y(\reg_module/_02367_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_19389_  (.A(\reg_module/_02367_ ),
    .X(\reg_module/_02368_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19390_  (.A(\reg_module/_02368_ ),
    .X(\reg_module/_02369_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19391_  (.A(\reg_module/_02369_ ),
    .B(net1758),
    .Y(\reg_module/_02370_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19392_  (.A(\reg_module/_01919_ ),
    .B(\reg_module/_09628_ ),
    .Y(\reg_module/_02371_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19393_  (.A1(\reg_module/_02370_ ),
    .A2(\reg_module/_02371_ ),
    .B1(\reg_module/_02366_ ),
    .Y(\reg_module/_00960_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19394_  (.A(\reg_module/_02369_ ),
    .B(net1360),
    .Y(\reg_module/_02372_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19395_  (.A(\reg_module/_01868_ ),
    .X(\reg_module/_02373_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19396_  (.A(\reg_module/_02373_ ),
    .B(\reg_module/_09631_ ),
    .Y(\reg_module/_02374_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19397_  (.A1(\reg_module/_02372_ ),
    .A2(\reg_module/_02374_ ),
    .B1(\reg_module/_02366_ ),
    .Y(\reg_module/_00961_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19398_  (.A(\reg_module/_02369_ ),
    .B(net1591),
    .Y(\reg_module/_02375_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19399_  (.A(\reg_module/_02373_ ),
    .B(\reg_module/_09634_ ),
    .Y(\reg_module/_02376_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19400_  (.A1(\reg_module/_02375_ ),
    .A2(\reg_module/_02376_ ),
    .B1(\reg_module/_02366_ ),
    .Y(\reg_module/_00962_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19401_  (.A(\reg_module/_02369_ ),
    .B(net1870),
    .Y(\reg_module/_02377_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19402_  (.A(\reg_module/_02373_ ),
    .B(\reg_module/_09637_ ),
    .Y(\reg_module/_02378_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19403_  (.A1(\reg_module/_02377_ ),
    .A2(\reg_module/_02378_ ),
    .B1(\reg_module/_02366_ ),
    .Y(\reg_module/_00963_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19404_  (.A(\reg_module/_02369_ ),
    .B(net1630),
    .Y(\reg_module/_02379_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19405_  (.A(\reg_module/_02373_ ),
    .B(\reg_module/_09641_ ),
    .Y(\reg_module/_02380_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19406_  (.A1(\reg_module/_02379_ ),
    .A2(\reg_module/_02380_ ),
    .B1(\reg_module/_02366_ ),
    .Y(\reg_module/_00964_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19407_  (.A(\reg_module/_02369_ ),
    .B(net1785),
    .Y(\reg_module/_02381_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19408_  (.A(\reg_module/_02373_ ),
    .B(\reg_module/_09645_ ),
    .Y(\reg_module/_02382_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19409_  (.A(\reg_module/_02192_ ),
    .X(\reg_module/_02383_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19410_  (.A1(\reg_module/_02381_ ),
    .A2(\reg_module/_02382_ ),
    .B1(\reg_module/_02383_ ),
    .Y(\reg_module/_00965_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19411_  (.A(\reg_module/_02368_ ),
    .X(\reg_module/_02384_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19412_  (.A(\reg_module/_02384_ ),
    .B(net1542),
    .Y(\reg_module/_02385_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19413_  (.A(\reg_module/_02373_ ),
    .B(\reg_module/_09649_ ),
    .Y(\reg_module/_02386_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19414_  (.A1(\reg_module/_02385_ ),
    .A2(\reg_module/_02386_ ),
    .B1(\reg_module/_02383_ ),
    .Y(\reg_module/_00966_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19415_  (.A(\reg_module/_02384_ ),
    .B(net1603),
    .Y(\reg_module/_02387_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19416_  (.A(\reg_module/_01868_ ),
    .X(\reg_module/_02388_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19417_  (.A(\reg_module/_02388_ ),
    .B(\reg_module/_09652_ ),
    .Y(\reg_module/_02389_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19418_  (.A1(\reg_module/_02387_ ),
    .A2(\reg_module/_02389_ ),
    .B1(\reg_module/_02383_ ),
    .Y(\reg_module/_00967_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19419_  (.A(\reg_module/_02384_ ),
    .B(net1835),
    .Y(\reg_module/_02390_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19420_  (.A(\reg_module/_02388_ ),
    .B(\reg_module/_09655_ ),
    .Y(\reg_module/_02391_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19421_  (.A1(\reg_module/_02390_ ),
    .A2(\reg_module/_02391_ ),
    .B1(\reg_module/_02383_ ),
    .Y(\reg_module/_00968_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19422_  (.A(\reg_module/_02384_ ),
    .B(net1627),
    .Y(\reg_module/_02392_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19423_  (.A(\reg_module/_02388_ ),
    .B(\reg_module/_09658_ ),
    .Y(\reg_module/_02393_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19424_  (.A1(\reg_module/_02392_ ),
    .A2(\reg_module/_02393_ ),
    .B1(\reg_module/_02383_ ),
    .Y(\reg_module/_00969_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19425_  (.A(\reg_module/_02384_ ),
    .B(net1457),
    .Y(\reg_module/_02394_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19426_  (.A(\reg_module/_02388_ ),
    .B(\reg_module/_09662_ ),
    .Y(\reg_module/_02395_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19427_  (.A1(\reg_module/_02394_ ),
    .A2(\reg_module/_02395_ ),
    .B1(\reg_module/_02383_ ),
    .Y(\reg_module/_00970_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19428_  (.A(\reg_module/_02384_ ),
    .B(net1913),
    .Y(\reg_module/_02396_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19429_  (.A(\reg_module/_02388_ ),
    .B(\reg_module/_09666_ ),
    .Y(\reg_module/_02397_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19430_  (.A(\reg_module/_02192_ ),
    .X(\reg_module/_02398_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19431_  (.A1(\reg_module/_02396_ ),
    .A2(\reg_module/_02397_ ),
    .B1(\reg_module/_02398_ ),
    .Y(\reg_module/_00971_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19432_  (.A(\reg_module/_02368_ ),
    .X(\reg_module/_02399_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19433_  (.A(\reg_module/_02399_ ),
    .B(net1576),
    .Y(\reg_module/_02400_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19434_  (.A(\reg_module/_02388_ ),
    .B(\reg_module/_09670_ ),
    .Y(\reg_module/_02401_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19435_  (.A1(\reg_module/_02400_ ),
    .A2(\reg_module/_02401_ ),
    .B1(\reg_module/_02398_ ),
    .Y(\reg_module/_00972_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19436_  (.A(\reg_module/_02399_ ),
    .B(net1608),
    .Y(\reg_module/_02402_ ));
 sky130_fd_sc_hd__clkbuf_2 \reg_module/_19437_  (.A(\reg_module/_01301_ ),
    .X(\reg_module/_02403_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19438_  (.A(\reg_module/_02403_ ),
    .B(\reg_module/_09673_ ),
    .Y(\reg_module/_02404_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19439_  (.A1(\reg_module/_02402_ ),
    .A2(\reg_module/_02404_ ),
    .B1(\reg_module/_02398_ ),
    .Y(\reg_module/_00973_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19440_  (.A(\reg_module/_02399_ ),
    .B(net1562),
    .Y(\reg_module/_02405_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19441_  (.A(\reg_module/_02403_ ),
    .B(\reg_module/_09676_ ),
    .Y(\reg_module/_02406_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19442_  (.A1(\reg_module/_02405_ ),
    .A2(\reg_module/_02406_ ),
    .B1(\reg_module/_02398_ ),
    .Y(\reg_module/_00974_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19443_  (.A(\reg_module/_02399_ ),
    .B(net1525),
    .Y(\reg_module/_02407_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19444_  (.A(\reg_module/_02403_ ),
    .B(\reg_module/_09679_ ),
    .Y(\reg_module/_02408_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19445_  (.A1(\reg_module/_02407_ ),
    .A2(\reg_module/_02408_ ),
    .B1(\reg_module/_02398_ ),
    .Y(\reg_module/_00975_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19446_  (.A(\reg_module/_02399_ ),
    .B(net1462),
    .Y(\reg_module/_02409_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19447_  (.A(\reg_module/_02403_ ),
    .B(\reg_module/_09683_ ),
    .Y(\reg_module/_02410_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19448_  (.A1(\reg_module/_02409_ ),
    .A2(\reg_module/_02410_ ),
    .B1(\reg_module/_02398_ ),
    .Y(\reg_module/_00976_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19449_  (.A(\reg_module/_02399_ ),
    .B(net1458),
    .Y(\reg_module/_02411_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19450_  (.A(\reg_module/_02403_ ),
    .B(net280),
    .Y(\reg_module/_02412_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19451_  (.A(\reg_module/_02192_ ),
    .X(\reg_module/_02413_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19452_  (.A1(\reg_module/_02411_ ),
    .A2(\reg_module/_02412_ ),
    .B1(\reg_module/_02413_ ),
    .Y(\reg_module/_00977_ ));
 sky130_fd_sc_hd__buf_4 \reg_module/_19453_  (.A(\reg_module/_02368_ ),
    .X(\reg_module/_02414_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19454_  (.A(\reg_module/_02414_ ),
    .B(net1415),
    .Y(\reg_module/_02415_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19455_  (.A(\reg_module/_02403_ ),
    .B(\reg_module/_09691_ ),
    .Y(\reg_module/_02416_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19456_  (.A1(\reg_module/_02415_ ),
    .A2(\reg_module/_02416_ ),
    .B1(\reg_module/_02413_ ),
    .Y(\reg_module/_00978_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19457_  (.A(\reg_module/_02414_ ),
    .B(net1228),
    .Y(\reg_module/_02417_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19458_  (.A(\reg_module/_01301_ ),
    .X(\reg_module/_02418_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19459_  (.A(\reg_module/_02418_ ),
    .B(\reg_module/_09694_ ),
    .Y(\reg_module/_02419_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19460_  (.A1(\reg_module/_02417_ ),
    .A2(\reg_module/_02419_ ),
    .B1(\reg_module/_02413_ ),
    .Y(\reg_module/_00979_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19461_  (.A(\reg_module/_02414_ ),
    .B(net1423),
    .Y(\reg_module/_02420_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19462_  (.A(\reg_module/_02418_ ),
    .B(\reg_module/_09697_ ),
    .Y(\reg_module/_02421_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19463_  (.A1(\reg_module/_02420_ ),
    .A2(\reg_module/_02421_ ),
    .B1(\reg_module/_02413_ ),
    .Y(\reg_module/_00980_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19464_  (.A(\reg_module/_02414_ ),
    .B(net1276),
    .Y(\reg_module/_02422_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19465_  (.A(\reg_module/_02418_ ),
    .B(\reg_module/_09700_ ),
    .Y(\reg_module/_02423_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19466_  (.A1(\reg_module/_02422_ ),
    .A2(\reg_module/_02423_ ),
    .B1(\reg_module/_02413_ ),
    .Y(\reg_module/_00981_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19467_  (.A(\reg_module/_02414_ ),
    .B(net1438),
    .Y(\reg_module/_02424_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19468_  (.A(\reg_module/_02418_ ),
    .B(\reg_module/_09705_ ),
    .Y(\reg_module/_02425_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19469_  (.A1(\reg_module/_02424_ ),
    .A2(\reg_module/_02425_ ),
    .B1(\reg_module/_02413_ ),
    .Y(\reg_module/_00982_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19470_  (.A(\reg_module/_02414_ ),
    .B(net1755),
    .Y(\reg_module/_02426_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19471_  (.A(\reg_module/_02418_ ),
    .B(\reg_module/_09709_ ),
    .Y(\reg_module/_02427_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19472_  (.A(\reg_module/_02192_ ),
    .X(\reg_module/_02428_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19473_  (.A1(\reg_module/_02426_ ),
    .A2(\reg_module/_02427_ ),
    .B1(\reg_module/_02428_ ),
    .Y(\reg_module/_00983_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19474_  (.A(\reg_module/_02367_ ),
    .X(\reg_module/_02429_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19475_  (.A(\reg_module/_02429_ ),
    .B(net1336),
    .Y(\reg_module/_02430_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19476_  (.A(\reg_module/_02418_ ),
    .B(\reg_module/_09713_ ),
    .Y(\reg_module/_02431_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19477_  (.A1(\reg_module/_02430_ ),
    .A2(\reg_module/_02431_ ),
    .B1(\reg_module/_02428_ ),
    .Y(\reg_module/_00984_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19478_  (.A(\reg_module/_02429_ ),
    .B(net1255),
    .Y(\reg_module/_02432_ ));
 sky130_fd_sc_hd__buf_2 \reg_module/_19479_  (.A(\reg_module/_01301_ ),
    .X(\reg_module/_02433_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19480_  (.A(\reg_module/_02433_ ),
    .B(\reg_module/_09716_ ),
    .Y(\reg_module/_02434_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19481_  (.A1(\reg_module/_02432_ ),
    .A2(\reg_module/_02434_ ),
    .B1(\reg_module/_02428_ ),
    .Y(\reg_module/_00985_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19482_  (.A(\reg_module/_02429_ ),
    .B(net1925),
    .Y(\reg_module/_02435_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19483_  (.A(\reg_module/_02433_ ),
    .B(\reg_module/_09719_ ),
    .Y(\reg_module/_02436_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19484_  (.A1(\reg_module/_02435_ ),
    .A2(\reg_module/_02436_ ),
    .B1(\reg_module/_02428_ ),
    .Y(\reg_module/_00986_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19485_  (.A(\reg_module/_02429_ ),
    .B(net1386),
    .Y(\reg_module/_02437_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19486_  (.A(\reg_module/_02433_ ),
    .B(\reg_module/_09722_ ),
    .Y(\reg_module/_02438_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19487_  (.A1(\reg_module/_02437_ ),
    .A2(\reg_module/_02438_ ),
    .B1(\reg_module/_02428_ ),
    .Y(\reg_module/_00987_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19488_  (.A(\reg_module/_02429_ ),
    .B(net1317),
    .Y(\reg_module/_02439_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19489_  (.A(\reg_module/_02433_ ),
    .B(\reg_module/_09726_ ),
    .Y(\reg_module/_02440_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19490_  (.A1(\reg_module/_02439_ ),
    .A2(\reg_module/_02440_ ),
    .B1(\reg_module/_02428_ ),
    .Y(\reg_module/_00988_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19491_  (.A(\reg_module/_02429_ ),
    .B(net1745),
    .Y(\reg_module/_02441_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19492_  (.A(\reg_module/_02433_ ),
    .B(\reg_module/_09730_ ),
    .Y(\reg_module/_02442_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19493_  (.A1(\reg_module/_02441_ ),
    .A2(\reg_module/_02442_ ),
    .B1(\reg_module/_02193_ ),
    .Y(\reg_module/_00989_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19494_  (.A(\reg_module/_02368_ ),
    .B(net1384),
    .Y(\reg_module/_02443_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19495_  (.A(\reg_module/_02433_ ),
    .B(\reg_module/_09733_ ),
    .Y(\reg_module/_02444_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19496_  (.A1(\reg_module/_02443_ ),
    .A2(\reg_module/_02444_ ),
    .B1(\reg_module/_02193_ ),
    .Y(\reg_module/_00990_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19497_  (.A(\reg_module/_02368_ ),
    .B(net1477),
    .Y(\reg_module/_02445_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19498_  (.A(\reg_module/_01288_ ),
    .B(\reg_module/_09736_ ),
    .Y(\reg_module/_02446_ ));
 sky130_fd_sc_hd__a21oi_1 \reg_module/_19499_  (.A1(\reg_module/_02445_ ),
    .A2(\reg_module/_02446_ ),
    .B1(\reg_module/_02193_ ),
    .Y(\reg_module/_00991_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19500_  (.A(net1628),
    .B(net1032),
    .Y(\reg_module/_02447_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19501_  (.A(\reg_module/_02447_ ),
    .Y(\reg_module/_00992_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19502_  (.A(net1193),
    .B(net1034),
    .Y(\reg_module/_02448_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19503_  (.A(\reg_module/_02448_ ),
    .Y(\reg_module/_00993_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19504_  (.A(net1219),
    .B(net1037),
    .Y(\reg_module/_02449_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19505_  (.A(\reg_module/_02449_ ),
    .Y(\reg_module/_00994_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19506_  (.A(net1226),
    .B(net1036),
    .Y(\reg_module/_02450_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19507_  (.A(\reg_module/_02450_ ),
    .Y(\reg_module/_00995_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19508_  (.A(net1210),
    .B(net1037),
    .Y(\reg_module/_02451_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19509_  (.A(\reg_module/_02451_ ),
    .Y(\reg_module/_00996_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19510_  (.A(net1218),
    .B(net1052),
    .Y(\reg_module/_02452_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19511_  (.A(\reg_module/_02452_ ),
    .Y(\reg_module/_00997_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19512_  (.A(net1202),
    .B(net1042),
    .Y(\reg_module/_02453_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19513_  (.A(\reg_module/_02453_ ),
    .Y(\reg_module/_00998_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19514_  (.A(net1215),
    .B(net1043),
    .Y(\reg_module/_02454_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19515_  (.A(\reg_module/_02454_ ),
    .Y(\reg_module/_00999_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19516_  (.A(net1213),
    .B(net1053),
    .Y(\reg_module/_02455_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19517_  (.A(\reg_module/_02455_ ),
    .Y(\reg_module/_01000_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19518_  (.A(net1217),
    .B(net1044),
    .Y(\reg_module/_02456_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19519_  (.A(\reg_module/_02456_ ),
    .Y(\reg_module/_01001_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19520_  (.A(net1221),
    .B(net1044),
    .Y(\reg_module/_02457_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19521_  (.A(\reg_module/_02457_ ),
    .Y(\reg_module/_01002_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19522_  (.A(net1207),
    .B(net1056),
    .Y(\reg_module/_02458_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19523_  (.A(\reg_module/_02458_ ),
    .Y(\reg_module/_01003_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19524_  (.A(net1200),
    .B(net1045),
    .Y(\reg_module/_02459_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19525_  (.A(\reg_module/_02459_ ),
    .Y(\reg_module/_01004_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19526_  (.A(net1220),
    .B(net1066),
    .Y(\reg_module/_02460_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19527_  (.A(\reg_module/_02460_ ),
    .Y(\reg_module/_01005_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19528_  (.A(net1208),
    .B(net1061),
    .Y(\reg_module/_02461_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19529_  (.A(\reg_module/_02461_ ),
    .Y(\reg_module/_01006_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19530_  (.A(net1224),
    .B(net1066),
    .Y(\reg_module/_02462_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19531_  (.A(\reg_module/_02462_ ),
    .Y(\reg_module/_01007_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19532_  (.A(net1211),
    .B(net1061),
    .Y(\reg_module/_02463_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19533_  (.A(\reg_module/_02463_ ),
    .Y(\reg_module/_01008_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19534_  (.A(net1269),
    .B(net1059),
    .Y(\reg_module/_02464_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19535_  (.A(\reg_module/_02464_ ),
    .Y(\reg_module/_01009_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19536_  (.A(net1209),
    .B(net1058),
    .Y(\reg_module/_02465_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19537_  (.A(\reg_module/_02465_ ),
    .Y(\reg_module/_01010_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19538_  (.A(net1212),
    .B(net1058),
    .Y(\reg_module/_02466_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19539_  (.A(\reg_module/_02466_ ),
    .Y(\reg_module/_01011_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19540_  (.A(net1198),
    .B(net1026),
    .Y(\reg_module/_02467_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19541_  (.A(\reg_module/_02467_ ),
    .Y(\reg_module/_01012_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19542_  (.A(net1205),
    .B(net1026),
    .Y(\reg_module/_02468_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19543_  (.A(\reg_module/_02468_ ),
    .Y(\reg_module/_01013_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19544_  (.A(net1195),
    .B(net1026),
    .Y(\reg_module/_02469_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19545_  (.A(\reg_module/_02469_ ),
    .Y(\reg_module/_01014_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19546_  (.A(net1204),
    .B(net1026),
    .Y(\reg_module/_02470_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19547_  (.A(\reg_module/_02470_ ),
    .Y(\reg_module/_01015_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19548_  (.A(net1194),
    .B(net1014),
    .Y(\reg_module/_02471_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19549_  (.A(\reg_module/_02471_ ),
    .Y(\reg_module/_01016_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19550_  (.A(net1197),
    .B(net1014),
    .Y(\reg_module/_02472_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19551_  (.A(\reg_module/_02472_ ),
    .Y(\reg_module/_01017_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19552_  (.A(net1196),
    .B(net1014),
    .Y(\reg_module/_02473_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19553_  (.A(\reg_module/_02473_ ),
    .Y(\reg_module/_01018_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19554_  (.A(net1216),
    .B(net1014),
    .Y(\reg_module/_02474_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19555_  (.A(\reg_module/_02474_ ),
    .Y(\reg_module/_01019_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19556_  (.A(net1199),
    .B(net1012),
    .Y(\reg_module/_02475_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19557_  (.A(\reg_module/_02475_ ),
    .Y(\reg_module/_01020_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19558_  (.A(net1206),
    .B(net1013),
    .Y(\reg_module/_02476_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19559_  (.A(\reg_module/_02476_ ),
    .Y(\reg_module/_01021_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19560_  (.A(net1223),
    .B(net1012),
    .Y(\reg_module/_02477_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19561_  (.A(\reg_module/_02477_ ),
    .Y(\reg_module/_01022_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19562_  (.A(net1222),
    .B(net1012),
    .Y(\reg_module/_02478_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19563_  (.A(\reg_module/_02478_ ),
    .Y(\reg_module/_01023_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19564_  (.A(net1016),
    .B(\wReg_s1_out[0] ),
    .Y(\reg_module/_02479_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19565_  (.A(\reg_module/_02479_ ),
    .Y(\reg_module/_01024_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19566_  (.A(net1023),
    .B(\wReg_s1_out[1] ),
    .Y(\reg_module/_02480_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19567_  (.A(\reg_module/_02480_ ),
    .Y(\reg_module/_01025_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19568_  (.A(net1016),
    .B(\wReg_s1_out[2] ),
    .Y(\reg_module/_02481_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19569_  (.A(\reg_module/_02481_ ),
    .Y(\reg_module/_01026_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19570_  (.A(net1023),
    .B(\wReg_s1_out[3] ),
    .Y(\reg_module/_02482_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19571_  (.A(\reg_module/_02482_ ),
    .Y(\reg_module/_01027_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19572_  (.A(net1029),
    .B(\wReg_s1_out[4] ),
    .Y(\reg_module/_02483_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19573_  (.A(\reg_module/_02483_ ),
    .Y(\reg_module/_01028_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19574_  (.A(net1016),
    .B(\wReg_s2_out[0] ),
    .Y(\reg_module/_02484_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19575_  (.A(\reg_module/_02484_ ),
    .Y(\reg_module/_01029_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19576_  (.A(net1023),
    .B(\wReg_s2_out[1] ),
    .Y(\reg_module/_02485_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19577_  (.A(\reg_module/_02485_ ),
    .Y(\reg_module/_01030_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19578_  (.A(net1023),
    .B(\wReg_s2_out[2] ),
    .Y(\reg_module/_02486_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19579_  (.A(\reg_module/_02486_ ),
    .Y(\reg_module/_01031_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19580_  (.A(net1023),
    .B(\wReg_s2_out[3] ),
    .Y(\reg_module/_02487_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19581_  (.A(\reg_module/_02487_ ),
    .Y(\reg_module/_01032_ ));
 sky130_fd_sc_hd__nand2_1 \reg_module/_19582_  (.A(net1023),
    .B(\wReg_s2_out[4] ),
    .Y(\reg_module/_02488_ ));
 sky130_fd_sc_hd__inv_2 \reg_module/_19583_  (.A(\reg_module/_02488_ ),
    .Y(\reg_module/_01033_ ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19584_  (.CLK(clknet_leaf_176_clk),
    .D(\reg_module/_00000_ ),
    .Q(\reg_module/gprf[0] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19585_  (.CLK(clknet_leaf_175_clk),
    .D(\reg_module/_00001_ ),
    .Q(\reg_module/gprf[1] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19586_  (.CLK(clknet_leaf_172_clk),
    .D(\reg_module/_00002_ ),
    .Q(\reg_module/gprf[2] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19587_  (.CLK(clknet_leaf_171_clk),
    .D(\reg_module/_00003_ ),
    .Q(\reg_module/gprf[3] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19588_  (.CLK(clknet_leaf_159_clk),
    .D(\reg_module/_00004_ ),
    .Q(\reg_module/gprf[4] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19589_  (.CLK(clknet_leaf_159_clk),
    .D(\reg_module/_00005_ ),
    .Q(\reg_module/gprf[5] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19590_  (.CLK(clknet_leaf_149_clk),
    .D(\reg_module/_00006_ ),
    .Q(\reg_module/gprf[6] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19591_  (.CLK(clknet_leaf_148_clk),
    .D(\reg_module/_00007_ ),
    .Q(\reg_module/gprf[7] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19592_  (.CLK(clknet_leaf_148_clk),
    .D(\reg_module/_00008_ ),
    .Q(\reg_module/gprf[8] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19593_  (.CLK(clknet_leaf_148_clk),
    .D(\reg_module/_00009_ ),
    .Q(\reg_module/gprf[9] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19594_  (.CLK(clknet_leaf_144_clk),
    .D(\reg_module/_00010_ ),
    .Q(\reg_module/gprf[10] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19595_  (.CLK(clknet_leaf_144_clk),
    .D(\reg_module/_00011_ ),
    .Q(\reg_module/gprf[11] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19596_  (.CLK(clknet_leaf_100_clk),
    .D(\reg_module/_00012_ ),
    .Q(\reg_module/gprf[12] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19597_  (.CLK(clknet_leaf_100_clk),
    .D(\reg_module/_00013_ ),
    .Q(\reg_module/gprf[13] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19598_  (.CLK(clknet_leaf_100_clk),
    .D(\reg_module/_00014_ ),
    .Q(\reg_module/gprf[14] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19599_  (.CLK(clknet_leaf_100_clk),
    .D(\reg_module/_00015_ ),
    .Q(\reg_module/gprf[15] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19600_  (.CLK(clknet_leaf_99_clk),
    .D(\reg_module/_00016_ ),
    .Q(\reg_module/gprf[16] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19601_  (.CLK(clknet_leaf_99_clk),
    .D(\reg_module/_00017_ ),
    .Q(\reg_module/gprf[17] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19602_  (.CLK(clknet_leaf_80_clk),
    .D(\reg_module/_00018_ ),
    .Q(\reg_module/gprf[18] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19603_  (.CLK(clknet_leaf_80_clk),
    .D(\reg_module/_00019_ ),
    .Q(\reg_module/gprf[19] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19604_  (.CLK(clknet_leaf_80_clk),
    .D(\reg_module/_00020_ ),
    .Q(\reg_module/gprf[20] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19605_  (.CLK(clknet_leaf_80_clk),
    .D(\reg_module/_00021_ ),
    .Q(\reg_module/gprf[21] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19606_  (.CLK(clknet_leaf_19_clk),
    .D(\reg_module/_00022_ ),
    .Q(\reg_module/gprf[22] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19607_  (.CLK(clknet_leaf_18_clk),
    .D(\reg_module/_00023_ ),
    .Q(\reg_module/gprf[23] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19608_  (.CLK(clknet_leaf_222_clk),
    .D(\reg_module/_00024_ ),
    .Q(\reg_module/gprf[24] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19609_  (.CLK(clknet_leaf_222_clk),
    .D(\reg_module/_00025_ ),
    .Q(\reg_module/gprf[25] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19610_  (.CLK(clknet_leaf_223_clk),
    .D(\reg_module/_00026_ ),
    .Q(\reg_module/gprf[26] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19611_  (.CLK(clknet_leaf_1_clk),
    .D(\reg_module/_00027_ ),
    .Q(\reg_module/gprf[27] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19612_  (.CLK(clknet_leaf_220_clk),
    .D(\reg_module/_00028_ ),
    .Q(\reg_module/gprf[28] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19613_  (.CLK(clknet_leaf_220_clk),
    .D(\reg_module/_00029_ ),
    .Q(\reg_module/gprf[29] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19614_  (.CLK(clknet_leaf_218_clk),
    .D(\reg_module/_00030_ ),
    .Q(\reg_module/gprf[30] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19615_  (.CLK(clknet_leaf_218_clk),
    .D(\reg_module/_00031_ ),
    .Q(\reg_module/gprf[31] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19616_  (.CLK(clknet_leaf_174_clk),
    .D(\reg_module/_00032_ ),
    .Q(\reg_module/gprf[32] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19617_  (.CLK(clknet_leaf_174_clk),
    .D(\reg_module/_00033_ ),
    .Q(\reg_module/gprf[33] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19618_  (.CLK(clknet_leaf_173_clk),
    .D(\reg_module/_00034_ ),
    .Q(\reg_module/gprf[34] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19619_  (.CLK(clknet_leaf_173_clk),
    .D(\reg_module/_00035_ ),
    .Q(\reg_module/gprf[35] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19620_  (.CLK(clknet_leaf_163_clk),
    .D(\reg_module/_00036_ ),
    .Q(\reg_module/gprf[36] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19621_  (.CLK(clknet_leaf_163_clk),
    .D(\reg_module/_00037_ ),
    .Q(\reg_module/gprf[37] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19622_  (.CLK(clknet_leaf_147_clk),
    .D(\reg_module/_00038_ ),
    .Q(\reg_module/gprf[38] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19623_  (.CLK(clknet_leaf_148_clk),
    .D(\reg_module/_00039_ ),
    .Q(\reg_module/gprf[39] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19624_  (.CLK(clknet_leaf_147_clk),
    .D(\reg_module/_00040_ ),
    .Q(\reg_module/gprf[40] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19625_  (.CLK(clknet_leaf_147_clk),
    .D(\reg_module/_00041_ ),
    .Q(\reg_module/gprf[41] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19626_  (.CLK(clknet_leaf_144_clk),
    .D(\reg_module/_00042_ ),
    .Q(\reg_module/gprf[42] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19627_  (.CLK(clknet_leaf_142_clk),
    .D(\reg_module/_00043_ ),
    .Q(\reg_module/gprf[43] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19628_  (.CLK(clknet_leaf_99_clk),
    .D(\reg_module/_00044_ ),
    .Q(\reg_module/gprf[44] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19629_  (.CLK(clknet_leaf_99_clk),
    .D(\reg_module/_00045_ ),
    .Q(\reg_module/gprf[45] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19630_  (.CLK(clknet_leaf_99_clk),
    .D(\reg_module/_00046_ ),
    .Q(\reg_module/gprf[46] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19631_  (.CLK(clknet_leaf_99_clk),
    .D(\reg_module/_00047_ ),
    .Q(\reg_module/gprf[47] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19632_  (.CLK(clknet_leaf_98_clk),
    .D(\reg_module/_00048_ ),
    .Q(\reg_module/gprf[48] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19633_  (.CLK(clknet_leaf_98_clk),
    .D(\reg_module/_00049_ ),
    .Q(\reg_module/gprf[49] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19634_  (.CLK(clknet_leaf_78_clk),
    .D(\reg_module/_00050_ ),
    .Q(\reg_module/gprf[50] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19635_  (.CLK(clknet_leaf_78_clk),
    .D(\reg_module/_00051_ ),
    .Q(\reg_module/gprf[51] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19636_  (.CLK(clknet_leaf_69_clk),
    .D(\reg_module/_00052_ ),
    .Q(\reg_module/gprf[52] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19637_  (.CLK(clknet_leaf_68_clk),
    .D(\reg_module/_00053_ ),
    .Q(\reg_module/gprf[53] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19638_  (.CLK(clknet_leaf_67_clk),
    .D(\reg_module/_00054_ ),
    .Q(\reg_module/gprf[54] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19639_  (.CLK(clknet_leaf_67_clk),
    .D(\reg_module/_00055_ ),
    .Q(\reg_module/gprf[55] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19640_  (.CLK(clknet_leaf_222_clk),
    .D(\reg_module/_00056_ ),
    .Q(\reg_module/gprf[56] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19641_  (.CLK(clknet_leaf_5_clk),
    .D(\reg_module/_00057_ ),
    .Q(\reg_module/gprf[57] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19642_  (.CLK(clknet_leaf_223_clk),
    .D(\reg_module/_00058_ ),
    .Q(\reg_module/gprf[58] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19643_  (.CLK(clknet_leaf_1_clk),
    .D(\reg_module/_00059_ ),
    .Q(\reg_module/gprf[59] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19644_  (.CLK(clknet_leaf_2_clk),
    .D(\reg_module/_00060_ ),
    .Q(\reg_module/gprf[60] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19645_  (.CLK(clknet_leaf_2_clk),
    .D(\reg_module/_00061_ ),
    .Q(\reg_module/gprf[61] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19646_  (.CLK(clknet_leaf_213_clk),
    .D(\reg_module/_00062_ ),
    .Q(\reg_module/gprf[62] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19647_  (.CLK(clknet_leaf_213_clk),
    .D(\reg_module/_00063_ ),
    .Q(\reg_module/gprf[63] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19648_  (.CLK(clknet_leaf_176_clk),
    .D(\reg_module/_00064_ ),
    .Q(\reg_module/gprf[64] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19649_  (.CLK(clknet_leaf_215_clk),
    .D(\reg_module/_00065_ ),
    .Q(\reg_module/gprf[65] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19650_  (.CLK(clknet_leaf_173_clk),
    .D(\reg_module/_00066_ ),
    .Q(\reg_module/gprf[66] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19651_  (.CLK(clknet_leaf_174_clk),
    .D(\reg_module/_00067_ ),
    .Q(\reg_module/gprf[67] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19652_  (.CLK(clknet_leaf_155_clk),
    .D(\reg_module/_00068_ ),
    .Q(\reg_module/gprf[68] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19653_  (.CLK(clknet_leaf_155_clk),
    .D(\reg_module/_00069_ ),
    .Q(\reg_module/gprf[69] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19654_  (.CLK(clknet_leaf_148_clk),
    .D(\reg_module/_00070_ ),
    .Q(\reg_module/gprf[70] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19655_  (.CLK(clknet_leaf_148_clk),
    .D(\reg_module/_00071_ ),
    .Q(\reg_module/gprf[71] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19656_  (.CLK(clknet_leaf_148_clk),
    .D(\reg_module/_00072_ ),
    .Q(\reg_module/gprf[72] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19657_  (.CLK(clknet_leaf_145_clk),
    .D(\reg_module/_00073_ ),
    .Q(\reg_module/gprf[73] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19658_  (.CLK(clknet_leaf_143_clk),
    .D(\reg_module/_00074_ ),
    .Q(\reg_module/gprf[74] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19659_  (.CLK(clknet_leaf_143_clk),
    .D(\reg_module/_00075_ ),
    .Q(\reg_module/gprf[75] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19660_  (.CLK(clknet_leaf_104_clk),
    .D(\reg_module/_00076_ ),
    .Q(\reg_module/gprf[76] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19661_  (.CLK(clknet_leaf_104_clk),
    .D(\reg_module/_00077_ ),
    .Q(\reg_module/gprf[77] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19662_  (.CLK(clknet_leaf_100_clk),
    .D(\reg_module/_00078_ ),
    .Q(\reg_module/gprf[78] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19663_  (.CLK(clknet_leaf_104_clk),
    .D(\reg_module/_00079_ ),
    .Q(\reg_module/gprf[79] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19664_  (.CLK(clknet_leaf_103_clk),
    .D(\reg_module/_00080_ ),
    .Q(\reg_module/gprf[80] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19665_  (.CLK(clknet_leaf_101_clk),
    .D(\reg_module/_00081_ ),
    .Q(\reg_module/gprf[81] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19666_  (.CLK(clknet_leaf_75_clk),
    .D(\reg_module/_00082_ ),
    .Q(\reg_module/gprf[82] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19667_  (.CLK(clknet_leaf_81_clk),
    .D(\reg_module/_00083_ ),
    .Q(\reg_module/gprf[83] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19668_  (.CLK(clknet_leaf_76_clk),
    .D(\reg_module/_00084_ ),
    .Q(\reg_module/gprf[84] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19669_  (.CLK(clknet_leaf_76_clk),
    .D(\reg_module/_00085_ ),
    .Q(\reg_module/gprf[85] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19670_  (.CLK(clknet_leaf_17_clk),
    .D(\reg_module/_00086_ ),
    .Q(\reg_module/gprf[86] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19671_  (.CLK(clknet_leaf_17_clk),
    .D(\reg_module/_00087_ ),
    .Q(\reg_module/gprf[87] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19672_  (.CLK(clknet_leaf_6_clk),
    .D(\reg_module/_00088_ ),
    .Q(\reg_module/gprf[88] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19673_  (.CLK(clknet_leaf_6_clk),
    .D(\reg_module/_00089_ ),
    .Q(\reg_module/gprf[89] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19674_  (.CLK(clknet_leaf_5_clk),
    .D(\reg_module/_00090_ ),
    .Q(\reg_module/gprf[90] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19675_  (.CLK(clknet_leaf_5_clk),
    .D(\reg_module/_00091_ ),
    .Q(\reg_module/gprf[91] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19676_  (.CLK(clknet_leaf_206_clk),
    .D(\reg_module/_00092_ ),
    .Q(\reg_module/gprf[92] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19677_  (.CLK(clknet_leaf_219_clk),
    .D(\reg_module/_00093_ ),
    .Q(\reg_module/gprf[93] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19678_  (.CLK(clknet_leaf_218_clk),
    .D(\reg_module/_00094_ ),
    .Q(\reg_module/gprf[94] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19679_  (.CLK(clknet_leaf_213_clk),
    .D(\reg_module/_00095_ ),
    .Q(\reg_module/gprf[95] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19680_  (.CLK(clknet_leaf_215_clk),
    .D(\reg_module/_00096_ ),
    .Q(\reg_module/gprf[96] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19681_  (.CLK(clknet_leaf_215_clk),
    .D(\reg_module/_00097_ ),
    .Q(\reg_module/gprf[97] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19682_  (.CLK(clknet_leaf_162_clk),
    .D(\reg_module/_00098_ ),
    .Q(\reg_module/gprf[98] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19683_  (.CLK(clknet_leaf_162_clk),
    .D(\reg_module/_00099_ ),
    .Q(\reg_module/gprf[99] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19684_  (.CLK(clknet_leaf_163_clk),
    .D(\reg_module/_00100_ ),
    .Q(\reg_module/gprf[100] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19685_  (.CLK(clknet_leaf_155_clk),
    .D(\reg_module/_00101_ ),
    .Q(\reg_module/gprf[101] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19686_  (.CLK(clknet_leaf_150_clk),
    .D(\reg_module/_00102_ ),
    .Q(\reg_module/gprf[102] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19687_  (.CLK(clknet_leaf_150_clk),
    .D(\reg_module/_00103_ ),
    .Q(\reg_module/gprf[103] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19688_  (.CLK(clknet_leaf_145_clk),
    .D(\reg_module/_00104_ ),
    .Q(\reg_module/gprf[104] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19689_  (.CLK(clknet_leaf_145_clk),
    .D(\reg_module/_00105_ ),
    .Q(\reg_module/gprf[105] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19690_  (.CLK(clknet_leaf_145_clk),
    .D(\reg_module/_00106_ ),
    .Q(\reg_module/gprf[106] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19691_  (.CLK(clknet_leaf_146_clk),
    .D(\reg_module/_00107_ ),
    .Q(\reg_module/gprf[107] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19692_  (.CLK(clknet_leaf_103_clk),
    .D(\reg_module/_00108_ ),
    .Q(\reg_module/gprf[108] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19693_  (.CLK(clknet_leaf_103_clk),
    .D(\reg_module/_00109_ ),
    .Q(\reg_module/gprf[109] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19694_  (.CLK(clknet_leaf_101_clk),
    .D(\reg_module/_00110_ ),
    .Q(\reg_module/gprf[110] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19695_  (.CLK(clknet_leaf_101_clk),
    .D(\reg_module/_00111_ ),
    .Q(\reg_module/gprf[111] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19696_  (.CLK(clknet_leaf_101_clk),
    .D(\reg_module/_00112_ ),
    .Q(\reg_module/gprf[112] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19697_  (.CLK(clknet_leaf_101_clk),
    .D(\reg_module/_00113_ ),
    .Q(\reg_module/gprf[113] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19698_  (.CLK(clknet_leaf_81_clk),
    .D(\reg_module/_00114_ ),
    .Q(\reg_module/gprf[114] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19699_  (.CLK(clknet_leaf_81_clk),
    .D(\reg_module/_00115_ ),
    .Q(\reg_module/gprf[115] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19700_  (.CLK(clknet_leaf_70_clk),
    .D(\reg_module/_00116_ ),
    .Q(\reg_module/gprf[116] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19701_  (.CLK(clknet_leaf_66_clk),
    .D(\reg_module/_00117_ ),
    .Q(\reg_module/gprf[117] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19702_  (.CLK(clknet_leaf_19_clk),
    .D(\reg_module/_00118_ ),
    .Q(\reg_module/gprf[118] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19703_  (.CLK(clknet_leaf_19_clk),
    .D(\reg_module/_00119_ ),
    .Q(\reg_module/gprf[119] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19704_  (.CLK(clknet_leaf_16_clk),
    .D(\reg_module/_00120_ ),
    .Q(\reg_module/gprf[120] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19705_  (.CLK(clknet_leaf_16_clk),
    .D(\reg_module/_00121_ ),
    .Q(\reg_module/gprf[121] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19706_  (.CLK(clknet_leaf_3_clk),
    .D(\reg_module/_00122_ ),
    .Q(\reg_module/gprf[122] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19707_  (.CLK(clknet_leaf_2_clk),
    .D(\reg_module/_00123_ ),
    .Q(\reg_module/gprf[123] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19708_  (.CLK(clknet_leaf_220_clk),
    .D(\reg_module/_00124_ ),
    .Q(\reg_module/gprf[124] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19709_  (.CLK(clknet_leaf_219_clk),
    .D(\reg_module/_00125_ ),
    .Q(\reg_module/gprf[125] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19710_  (.CLK(clknet_leaf_219_clk),
    .D(\reg_module/_00126_ ),
    .Q(\reg_module/gprf[126] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19711_  (.CLK(clknet_leaf_208_clk),
    .D(\reg_module/_00127_ ),
    .Q(\reg_module/gprf[127] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19712_  (.CLK(clknet_leaf_175_clk),
    .D(\reg_module/_00128_ ),
    .Q(\reg_module/gprf[128] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19713_  (.CLK(clknet_leaf_175_clk),
    .D(\reg_module/_00129_ ),
    .Q(\reg_module/gprf[129] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19714_  (.CLK(clknet_leaf_171_clk),
    .D(\reg_module/_00130_ ),
    .Q(\reg_module/gprf[130] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19715_  (.CLK(clknet_leaf_170_clk),
    .D(\reg_module/_00131_ ),
    .Q(\reg_module/gprf[131] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19716_  (.CLK(clknet_leaf_160_clk),
    .D(\reg_module/_00132_ ),
    .Q(\reg_module/gprf[132] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19717_  (.CLK(clknet_leaf_160_clk),
    .D(\reg_module/_00133_ ),
    .Q(\reg_module/gprf[133] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19718_  (.CLK(clknet_leaf_157_clk),
    .D(\reg_module/_00134_ ),
    .Q(\reg_module/gprf[134] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19719_  (.CLK(clknet_leaf_158_clk),
    .D(\reg_module/_00135_ ),
    .Q(\reg_module/gprf[135] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19720_  (.CLK(clknet_leaf_157_clk),
    .D(\reg_module/_00136_ ),
    .Q(\reg_module/gprf[136] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19721_  (.CLK(clknet_leaf_157_clk),
    .D(\reg_module/_00137_ ),
    .Q(\reg_module/gprf[137] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19722_  (.CLK(clknet_leaf_149_clk),
    .D(\reg_module/_00138_ ),
    .Q(\reg_module/gprf[138] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19723_  (.CLK(clknet_leaf_157_clk),
    .D(\reg_module/_00139_ ),
    .Q(\reg_module/gprf[139] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19724_  (.CLK(clknet_leaf_105_clk),
    .D(\reg_module/_00140_ ),
    .Q(\reg_module/gprf[140] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19725_  (.CLK(clknet_leaf_104_clk),
    .D(\reg_module/_00141_ ),
    .Q(\reg_module/gprf[141] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19726_  (.CLK(clknet_leaf_104_clk),
    .D(\reg_module/_00142_ ),
    .Q(\reg_module/gprf[142] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19727_  (.CLK(clknet_leaf_105_clk),
    .D(\reg_module/_00143_ ),
    .Q(\reg_module/gprf[143] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19728_  (.CLK(clknet_leaf_143_clk),
    .D(\reg_module/_00144_ ),
    .Q(\reg_module/gprf[144] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19729_  (.CLK(clknet_leaf_143_clk),
    .D(\reg_module/_00145_ ),
    .Q(\reg_module/gprf[145] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19730_  (.CLK(clknet_leaf_193_clk),
    .D(\reg_module/_00146_ ),
    .Q(\reg_module/gprf[146] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19731_  (.CLK(clknet_leaf_193_clk),
    .D(\reg_module/_00147_ ),
    .Q(\reg_module/gprf[147] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19732_  (.CLK(clknet_leaf_193_clk),
    .D(\reg_module/_00148_ ),
    .Q(\reg_module/gprf[148] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19733_  (.CLK(clknet_leaf_193_clk),
    .D(\reg_module/_00149_ ),
    .Q(\reg_module/gprf[149] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19734_  (.CLK(clknet_leaf_193_clk),
    .D(\reg_module/_00150_ ),
    .Q(\reg_module/gprf[150] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19735_  (.CLK(clknet_leaf_192_clk),
    .D(\reg_module/_00151_ ),
    .Q(\reg_module/gprf[151] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19736_  (.CLK(clknet_leaf_0_clk),
    .D(\reg_module/_00152_ ),
    .Q(\reg_module/gprf[152] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19737_  (.CLK(clknet_leaf_0_clk),
    .D(\reg_module/_00153_ ),
    .Q(\reg_module/gprf[153] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19738_  (.CLK(clknet_leaf_0_clk),
    .D(\reg_module/_00154_ ),
    .Q(\reg_module/gprf[154] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19739_  (.CLK(clknet_leaf_1_clk),
    .D(\reg_module/_00155_ ),
    .Q(\reg_module/gprf[155] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19740_  (.CLK(clknet_leaf_221_clk),
    .D(\reg_module/_00156_ ),
    .Q(\reg_module/gprf[156] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19741_  (.CLK(clknet_leaf_221_clk),
    .D(\reg_module/_00157_ ),
    .Q(\reg_module/gprf[157] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19742_  (.CLK(clknet_leaf_217_clk),
    .D(\reg_module/_00158_ ),
    .Q(\reg_module/gprf[158] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19743_  (.CLK(clknet_leaf_217_clk),
    .D(\reg_module/_00159_ ),
    .Q(\reg_module/gprf[159] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19744_  (.CLK(clknet_leaf_174_clk),
    .D(\reg_module/_00160_ ),
    .Q(\reg_module/gprf[160] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19745_  (.CLK(clknet_leaf_174_clk),
    .D(\reg_module/_00161_ ),
    .Q(\reg_module/gprf[161] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19746_  (.CLK(clknet_leaf_172_clk),
    .D(\reg_module/_00162_ ),
    .Q(\reg_module/gprf[162] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19747_  (.CLK(clknet_leaf_171_clk),
    .D(\reg_module/_00163_ ),
    .Q(\reg_module/gprf[163] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19748_  (.CLK(clknet_leaf_169_clk),
    .D(\reg_module/_00164_ ),
    .Q(\reg_module/gprf[164] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19749_  (.CLK(clknet_leaf_170_clk),
    .D(\reg_module/_00165_ ),
    .Q(\reg_module/gprf[165] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19750_  (.CLK(clknet_leaf_155_clk),
    .D(\reg_module/_00166_ ),
    .Q(\reg_module/gprf[166] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19751_  (.CLK(clknet_leaf_155_clk),
    .D(\reg_module/_00167_ ),
    .Q(\reg_module/gprf[167] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19752_  (.CLK(clknet_leaf_156_clk),
    .D(\reg_module/_00168_ ),
    .Q(\reg_module/gprf[168] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19753_  (.CLK(clknet_leaf_156_clk),
    .D(\reg_module/_00169_ ),
    .Q(\reg_module/gprf[169] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19754_  (.CLK(clknet_leaf_150_clk),
    .D(\reg_module/_00170_ ),
    .Q(\reg_module/gprf[170] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19755_  (.CLK(clknet_leaf_156_clk),
    .D(\reg_module/_00171_ ),
    .Q(\reg_module/gprf[171] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19756_  (.CLK(clknet_leaf_106_clk),
    .D(\reg_module/_00172_ ),
    .Q(\reg_module/gprf[172] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19757_  (.CLK(clknet_leaf_106_clk),
    .D(\reg_module/_00173_ ),
    .Q(\reg_module/gprf[173] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19758_  (.CLK(clknet_leaf_106_clk),
    .D(\reg_module/_00174_ ),
    .Q(\reg_module/gprf[174] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19759_  (.CLK(clknet_leaf_106_clk),
    .D(\reg_module/_00175_ ),
    .Q(\reg_module/gprf[175] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19760_  (.CLK(clknet_leaf_141_clk),
    .D(\reg_module/_00176_ ),
    .Q(\reg_module/gprf[176] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19761_  (.CLK(clknet_leaf_141_clk),
    .D(\reg_module/_00177_ ),
    .Q(\reg_module/gprf[177] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19762_  (.CLK(clknet_leaf_123_clk),
    .D(\reg_module/_00178_ ),
    .Q(\reg_module/gprf[178] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19763_  (.CLK(clknet_leaf_124_clk),
    .D(\reg_module/_00179_ ),
    .Q(\reg_module/gprf[179] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19764_  (.CLK(clknet_leaf_123_clk),
    .D(\reg_module/_00180_ ),
    .Q(\reg_module/gprf[180] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19765_  (.CLK(clknet_leaf_195_clk),
    .D(\reg_module/_00181_ ),
    .Q(\reg_module/gprf[181] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19766_  (.CLK(clknet_leaf_195_clk),
    .D(\reg_module/_00182_ ),
    .Q(\reg_module/gprf[182] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19767_  (.CLK(clknet_leaf_123_clk),
    .D(\reg_module/_00183_ ),
    .Q(\reg_module/gprf[183] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19768_  (.CLK(clknet_leaf_222_clk),
    .D(\reg_module/_00184_ ),
    .Q(\reg_module/gprf[184] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19769_  (.CLK(clknet_leaf_223_clk),
    .D(\reg_module/_00185_ ),
    .Q(\reg_module/gprf[185] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19770_  (.CLK(clknet_leaf_223_clk),
    .D(\reg_module/_00186_ ),
    .Q(\reg_module/gprf[186] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19771_  (.CLK(clknet_leaf_1_clk),
    .D(\reg_module/_00187_ ),
    .Q(\reg_module/gprf[187] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19772_  (.CLK(clknet_leaf_2_clk),
    .D(\reg_module/_00188_ ),
    .Q(\reg_module/gprf[188] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19773_  (.CLK(clknet_leaf_221_clk),
    .D(\reg_module/_00189_ ),
    .Q(\reg_module/gprf[189] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19774_  (.CLK(clknet_leaf_217_clk),
    .D(\reg_module/_00190_ ),
    .Q(\reg_module/gprf[190] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19775_  (.CLK(clknet_leaf_217_clk),
    .D(\reg_module/_00191_ ),
    .Q(\reg_module/gprf[191] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19776_  (.CLK(clknet_leaf_176_clk),
    .D(\reg_module/_00192_ ),
    .Q(\reg_module/gprf[192] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19777_  (.CLK(clknet_leaf_175_clk),
    .D(\reg_module/_00193_ ),
    .Q(\reg_module/gprf[193] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19778_  (.CLK(clknet_leaf_172_clk),
    .D(\reg_module/_00194_ ),
    .Q(\reg_module/gprf[194] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19779_  (.CLK(clknet_leaf_172_clk),
    .D(\reg_module/_00195_ ),
    .Q(\reg_module/gprf[195] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19780_  (.CLK(clknet_leaf_159_clk),
    .D(\reg_module/_00196_ ),
    .Q(\reg_module/gprf[196] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19781_  (.CLK(clknet_leaf_159_clk),
    .D(\reg_module/_00197_ ),
    .Q(\reg_module/gprf[197] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19782_  (.CLK(clknet_leaf_155_clk),
    .D(\reg_module/_00198_ ),
    .Q(\reg_module/gprf[198] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19783_  (.CLK(clknet_leaf_155_clk),
    .D(\reg_module/_00199_ ),
    .Q(\reg_module/gprf[199] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19784_  (.CLK(clknet_leaf_156_clk),
    .D(\reg_module/_00200_ ),
    .Q(\reg_module/gprf[200] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19785_  (.CLK(clknet_leaf_156_clk),
    .D(\reg_module/_00201_ ),
    .Q(\reg_module/gprf[201] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19786_  (.CLK(clknet_leaf_150_clk),
    .D(\reg_module/_00202_ ),
    .Q(\reg_module/gprf[202] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19787_  (.CLK(clknet_leaf_150_clk),
    .D(\reg_module/_00203_ ),
    .Q(\reg_module/gprf[203] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19788_  (.CLK(clknet_leaf_106_clk),
    .D(\reg_module/_00204_ ),
    .Q(\reg_module/gprf[204] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19789_  (.CLK(clknet_leaf_106_clk),
    .D(\reg_module/_00205_ ),
    .Q(\reg_module/gprf[205] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19790_  (.CLK(clknet_leaf_106_clk),
    .D(\reg_module/_00206_ ),
    .Q(\reg_module/gprf[206] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19791_  (.CLK(clknet_leaf_106_clk),
    .D(\reg_module/_00207_ ),
    .Q(\reg_module/gprf[207] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19792_  (.CLK(clknet_leaf_141_clk),
    .D(\reg_module/_00208_ ),
    .Q(\reg_module/gprf[208] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19793_  (.CLK(clknet_leaf_141_clk),
    .D(\reg_module/_00209_ ),
    .Q(\reg_module/gprf[209] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19794_  (.CLK(clknet_leaf_124_clk),
    .D(\reg_module/_00210_ ),
    .Q(\reg_module/gprf[210] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19795_  (.CLK(clknet_leaf_124_clk),
    .D(\reg_module/_00211_ ),
    .Q(\reg_module/gprf[211] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19796_  (.CLK(clknet_leaf_124_clk),
    .D(\reg_module/_00212_ ),
    .Q(\reg_module/gprf[212] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19797_  (.CLK(clknet_leaf_124_clk),
    .D(\reg_module/_00213_ ),
    .Q(\reg_module/gprf[213] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19798_  (.CLK(clknet_leaf_195_clk),
    .D(\reg_module/_00214_ ),
    .Q(\reg_module/gprf[214] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19799_  (.CLK(clknet_leaf_195_clk),
    .D(\reg_module/_00215_ ),
    .Q(\reg_module/gprf[215] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19800_  (.CLK(clknet_leaf_222_clk),
    .D(\reg_module/_00216_ ),
    .Q(\reg_module/gprf[216] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19801_  (.CLK(clknet_leaf_222_clk),
    .D(\reg_module/_00217_ ),
    .Q(\reg_module/gprf[217] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19802_  (.CLK(clknet_leaf_223_clk),
    .D(\reg_module/_00218_ ),
    .Q(\reg_module/gprf[218] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19803_  (.CLK(clknet_leaf_1_clk),
    .D(\reg_module/_00219_ ),
    .Q(\reg_module/gprf[219] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19804_  (.CLK(clknet_leaf_221_clk),
    .D(\reg_module/_00220_ ),
    .Q(\reg_module/gprf[220] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19805_  (.CLK(clknet_leaf_221_clk),
    .D(\reg_module/_00221_ ),
    .Q(\reg_module/gprf[221] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19806_  (.CLK(clknet_leaf_218_clk),
    .D(\reg_module/_00222_ ),
    .Q(\reg_module/gprf[222] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19807_  (.CLK(clknet_leaf_217_clk),
    .D(\reg_module/_00223_ ),
    .Q(\reg_module/gprf[223] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19808_  (.CLK(clknet_leaf_175_clk),
    .D(\reg_module/_00224_ ),
    .Q(\reg_module/gprf[224] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19809_  (.CLK(clknet_leaf_175_clk),
    .D(\reg_module/_00225_ ),
    .Q(\reg_module/gprf[225] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19810_  (.CLK(clknet_leaf_171_clk),
    .D(\reg_module/_00226_ ),
    .Q(\reg_module/gprf[226] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19811_  (.CLK(clknet_leaf_170_clk),
    .D(\reg_module/_00227_ ),
    .Q(\reg_module/gprf[227] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19812_  (.CLK(clknet_leaf_160_clk),
    .D(\reg_module/_00228_ ),
    .Q(\reg_module/gprf[228] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19813_  (.CLK(clknet_leaf_160_clk),
    .D(\reg_module/_00229_ ),
    .Q(\reg_module/gprf[229] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19814_  (.CLK(clknet_leaf_158_clk),
    .D(\reg_module/_00230_ ),
    .Q(\reg_module/gprf[230] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19815_  (.CLK(clknet_leaf_158_clk),
    .D(\reg_module/_00231_ ),
    .Q(\reg_module/gprf[231] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19816_  (.CLK(clknet_leaf_157_clk),
    .D(\reg_module/_00232_ ),
    .Q(\reg_module/gprf[232] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19817_  (.CLK(clknet_leaf_157_clk),
    .D(\reg_module/_00233_ ),
    .Q(\reg_module/gprf[233] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19818_  (.CLK(clknet_leaf_157_clk),
    .D(\reg_module/_00234_ ),
    .Q(\reg_module/gprf[234] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19819_  (.CLK(clknet_leaf_157_clk),
    .D(\reg_module/_00235_ ),
    .Q(\reg_module/gprf[235] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19820_  (.CLK(clknet_leaf_105_clk),
    .D(\reg_module/_00236_ ),
    .Q(\reg_module/gprf[236] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19821_  (.CLK(clknet_leaf_105_clk),
    .D(\reg_module/_00237_ ),
    .Q(\reg_module/gprf[237] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19822_  (.CLK(clknet_leaf_105_clk),
    .D(\reg_module/_00238_ ),
    .Q(\reg_module/gprf[238] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19823_  (.CLK(clknet_leaf_105_clk),
    .D(\reg_module/_00239_ ),
    .Q(\reg_module/gprf[239] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19824_  (.CLK(clknet_leaf_143_clk),
    .D(\reg_module/_00240_ ),
    .Q(\reg_module/gprf[240] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19825_  (.CLK(clknet_leaf_142_clk),
    .D(\reg_module/_00241_ ),
    .Q(\reg_module/gprf[241] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19826_  (.CLK(clknet_leaf_193_clk),
    .D(\reg_module/_00242_ ),
    .Q(\reg_module/gprf[242] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19827_  (.CLK(clknet_leaf_193_clk),
    .D(\reg_module/_00243_ ),
    .Q(\reg_module/gprf[243] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19828_  (.CLK(clknet_leaf_193_clk),
    .D(\reg_module/_00244_ ),
    .Q(\reg_module/gprf[244] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19829_  (.CLK(clknet_leaf_193_clk),
    .D(\reg_module/_00245_ ),
    .Q(\reg_module/gprf[245] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19830_  (.CLK(clknet_leaf_194_clk),
    .D(\reg_module/_00246_ ),
    .Q(\reg_module/gprf[246] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19831_  (.CLK(clknet_leaf_192_clk),
    .D(\reg_module/_00247_ ),
    .Q(\reg_module/gprf[247] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19832_  (.CLK(clknet_leaf_223_clk),
    .D(\reg_module/_00248_ ),
    .Q(\reg_module/gprf[248] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19833_  (.CLK(clknet_leaf_0_clk),
    .D(\reg_module/_00249_ ),
    .Q(\reg_module/gprf[249] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19834_  (.CLK(clknet_leaf_1_clk),
    .D(\reg_module/_00250_ ),
    .Q(\reg_module/gprf[250] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19835_  (.CLK(clknet_leaf_1_clk),
    .D(\reg_module/_00251_ ),
    .Q(\reg_module/gprf[251] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19836_  (.CLK(clknet_leaf_221_clk),
    .D(\reg_module/_00252_ ),
    .Q(\reg_module/gprf[252] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19837_  (.CLK(clknet_leaf_221_clk),
    .D(\reg_module/_00253_ ),
    .Q(\reg_module/gprf[253] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19838_  (.CLK(clknet_leaf_218_clk),
    .D(\reg_module/_00254_ ),
    .Q(\reg_module/gprf[254] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19839_  (.CLK(clknet_leaf_217_clk),
    .D(\reg_module/_00255_ ),
    .Q(\reg_module/gprf[255] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19840_  (.CLK(clknet_leaf_190_clk),
    .D(\reg_module/_00256_ ),
    .Q(\reg_module/gprf[256] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19841_  (.CLK(clknet_leaf_189_clk),
    .D(\reg_module/_00257_ ),
    .Q(\reg_module/gprf[257] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19842_  (.CLK(clknet_leaf_184_clk),
    .D(\reg_module/_00258_ ),
    .Q(\reg_module/gprf[258] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19843_  (.CLK(clknet_leaf_186_clk),
    .D(\reg_module/_00259_ ),
    .Q(\reg_module/gprf[259] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19844_  (.CLK(clknet_leaf_156_clk),
    .D(\reg_module/_00260_ ),
    .Q(\reg_module/gprf[260] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19845_  (.CLK(clknet_leaf_155_clk),
    .D(\reg_module/_00261_ ),
    .Q(\reg_module/gprf[261] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19846_  (.CLK(clknet_leaf_154_clk),
    .D(\reg_module/_00262_ ),
    .Q(\reg_module/gprf[262] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19847_  (.CLK(clknet_leaf_156_clk),
    .D(\reg_module/_00263_ ),
    .Q(\reg_module/gprf[263] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19848_  (.CLK(clknet_leaf_150_clk),
    .D(\reg_module/_00264_ ),
    .Q(\reg_module/gprf[264] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19849_  (.CLK(clknet_leaf_150_clk),
    .D(\reg_module/_00265_ ),
    .Q(\reg_module/gprf[265] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19850_  (.CLK(clknet_leaf_108_clk),
    .D(\reg_module/_00266_ ),
    .Q(\reg_module/gprf[266] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19851_  (.CLK(clknet_leaf_96_clk),
    .D(\reg_module/_00267_ ),
    .Q(\reg_module/gprf[267] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19852_  (.CLK(clknet_leaf_96_clk),
    .D(\reg_module/_00268_ ),
    .Q(\reg_module/gprf[268] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19853_  (.CLK(clknet_leaf_111_clk),
    .D(\reg_module/_00269_ ),
    .Q(\reg_module/gprf[269] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19854_  (.CLK(clknet_leaf_95_clk),
    .D(\reg_module/_00270_ ),
    .Q(\reg_module/gprf[270] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19855_  (.CLK(clknet_leaf_96_clk),
    .D(\reg_module/_00271_ ),
    .Q(\reg_module/gprf[271] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19856_  (.CLK(clknet_leaf_113_clk),
    .D(\reg_module/_00272_ ),
    .Q(\reg_module/gprf[272] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19857_  (.CLK(clknet_leaf_83_clk),
    .D(\reg_module/_00273_ ),
    .Q(\reg_module/gprf[273] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19858_  (.CLK(clknet_leaf_82_clk),
    .D(\reg_module/_00274_ ),
    .Q(\reg_module/gprf[274] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19859_  (.CLK(clknet_leaf_67_clk),
    .D(\reg_module/_00275_ ),
    .Q(\reg_module/gprf[275] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19860_  (.CLK(clknet_leaf_67_clk),
    .D(\reg_module/_00276_ ),
    .Q(\reg_module/gprf[276] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19861_  (.CLK(clknet_leaf_67_clk),
    .D(\reg_module/_00277_ ),
    .Q(\reg_module/gprf[277] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19862_  (.CLK(clknet_leaf_66_clk),
    .D(\reg_module/_00278_ ),
    .Q(\reg_module/gprf[278] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19863_  (.CLK(clknet_leaf_66_clk),
    .D(\reg_module/_00279_ ),
    .Q(\reg_module/gprf[279] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19864_  (.CLK(clknet_leaf_6_clk),
    .D(\reg_module/_00280_ ),
    .Q(\reg_module/gprf[280] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19865_  (.CLK(clknet_leaf_6_clk),
    .D(\reg_module/_00281_ ),
    .Q(\reg_module/gprf[281] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19866_  (.CLK(clknet_leaf_3_clk),
    .D(\reg_module/_00282_ ),
    .Q(\reg_module/gprf[282] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19867_  (.CLK(clknet_leaf_205_clk),
    .D(\reg_module/_00283_ ),
    .Q(\reg_module/gprf[283] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19868_  (.CLK(clknet_leaf_204_clk),
    .D(\reg_module/_00284_ ),
    .Q(\reg_module/gprf[284] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19869_  (.CLK(clknet_leaf_205_clk),
    .D(\reg_module/_00285_ ),
    .Q(\reg_module/gprf[285] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19870_  (.CLK(clknet_leaf_209_clk),
    .D(\reg_module/_00286_ ),
    .Q(\reg_module/gprf[286] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19871_  (.CLK(clknet_leaf_209_clk),
    .D(\reg_module/_00287_ ),
    .Q(\reg_module/gprf[287] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19872_  (.CLK(clknet_leaf_189_clk),
    .D(\reg_module/_00288_ ),
    .Q(\reg_module/gprf[288] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19873_  (.CLK(clknet_leaf_189_clk),
    .D(\reg_module/_00289_ ),
    .Q(\reg_module/gprf[289] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19874_  (.CLK(clknet_leaf_187_clk),
    .D(\reg_module/_00290_ ),
    .Q(\reg_module/gprf[290] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19875_  (.CLK(clknet_leaf_187_clk),
    .D(\reg_module/_00291_ ),
    .Q(\reg_module/gprf[291] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19876_  (.CLK(clknet_leaf_154_clk),
    .D(\reg_module/_00292_ ),
    .Q(\reg_module/gprf[292] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19877_  (.CLK(clknet_leaf_154_clk),
    .D(\reg_module/_00293_ ),
    .Q(\reg_module/gprf[293] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19878_  (.CLK(clknet_leaf_152_clk),
    .D(\reg_module/_00294_ ),
    .Q(\reg_module/gprf[294] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19879_  (.CLK(clknet_leaf_152_clk),
    .D(\reg_module/_00295_ ),
    .Q(\reg_module/gprf[295] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19880_  (.CLK(clknet_leaf_151_clk),
    .D(\reg_module/_00296_ ),
    .Q(\reg_module/gprf[296] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19881_  (.CLK(clknet_leaf_151_clk),
    .D(\reg_module/_00297_ ),
    .Q(\reg_module/gprf[297] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19882_  (.CLK(clknet_leaf_108_clk),
    .D(\reg_module/_00298_ ),
    .Q(\reg_module/gprf[298] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19883_  (.CLK(clknet_leaf_108_clk),
    .D(\reg_module/_00299_ ),
    .Q(\reg_module/gprf[299] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19884_  (.CLK(clknet_leaf_96_clk),
    .D(\reg_module/_00300_ ),
    .Q(\reg_module/gprf[300] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19885_  (.CLK(clknet_leaf_95_clk),
    .D(\reg_module/_00301_ ),
    .Q(\reg_module/gprf[301] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19886_  (.CLK(clknet_leaf_95_clk),
    .D(\reg_module/_00302_ ),
    .Q(\reg_module/gprf[302] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19887_  (.CLK(clknet_leaf_95_clk),
    .D(\reg_module/_00303_ ),
    .Q(\reg_module/gprf[303] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19888_  (.CLK(clknet_leaf_83_clk),
    .D(\reg_module/_00304_ ),
    .Q(\reg_module/gprf[304] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19889_  (.CLK(clknet_leaf_83_clk),
    .D(\reg_module/_00305_ ),
    .Q(\reg_module/gprf[305] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19890_  (.CLK(clknet_leaf_79_clk),
    .D(\reg_module/_00306_ ),
    .Q(\reg_module/gprf[306] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19891_  (.CLK(clknet_leaf_78_clk),
    .D(\reg_module/_00307_ ),
    .Q(\reg_module/gprf[307] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19892_  (.CLK(clknet_leaf_69_clk),
    .D(\reg_module/_00308_ ),
    .Q(\reg_module/gprf[308] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19893_  (.CLK(clknet_leaf_68_clk),
    .D(\reg_module/_00309_ ),
    .Q(\reg_module/gprf[309] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19894_  (.CLK(clknet_leaf_65_clk),
    .D(\reg_module/_00310_ ),
    .Q(\reg_module/gprf[310] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19895_  (.CLK(clknet_leaf_67_clk),
    .D(\reg_module/_00311_ ),
    .Q(\reg_module/gprf[311] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19896_  (.CLK(clknet_leaf_8_clk),
    .D(\reg_module/_00312_ ),
    .Q(\reg_module/gprf[312] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19897_  (.CLK(clknet_leaf_5_clk),
    .D(\reg_module/_00313_ ),
    .Q(\reg_module/gprf[313] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19898_  (.CLK(clknet_leaf_4_clk),
    .D(\reg_module/_00314_ ),
    .Q(\reg_module/gprf[314] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19899_  (.CLK(clknet_leaf_4_clk),
    .D(\reg_module/_00315_ ),
    .Q(\reg_module/gprf[315] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19900_  (.CLK(clknet_leaf_204_clk),
    .D(\reg_module/_00316_ ),
    .Q(\reg_module/gprf[316] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19901_  (.CLK(clknet_leaf_204_clk),
    .D(\reg_module/_00317_ ),
    .Q(\reg_module/gprf[317] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19902_  (.CLK(clknet_leaf_209_clk),
    .D(\reg_module/_00318_ ),
    .Q(\reg_module/gprf[318] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19903_  (.CLK(clknet_leaf_211_clk),
    .D(\reg_module/_00319_ ),
    .Q(\reg_module/gprf[319] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19904_  (.CLK(clknet_leaf_181_clk),
    .D(\reg_module/_00320_ ),
    .Q(\reg_module/gprf[320] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19905_  (.CLK(clknet_leaf_181_clk),
    .D(\reg_module/_00321_ ),
    .Q(\reg_module/gprf[321] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19906_  (.CLK(clknet_leaf_185_clk),
    .D(\reg_module/_00322_ ),
    .Q(\reg_module/gprf[322] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19907_  (.CLK(clknet_leaf_185_clk),
    .D(\reg_module/_00323_ ),
    .Q(\reg_module/gprf[323] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19908_  (.CLK(clknet_leaf_154_clk),
    .D(\reg_module/_00324_ ),
    .Q(\reg_module/gprf[324] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19909_  (.CLK(clknet_leaf_154_clk),
    .D(\reg_module/_00325_ ),
    .Q(\reg_module/gprf[325] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19910_  (.CLK(clknet_leaf_152_clk),
    .D(\reg_module/_00326_ ),
    .Q(\reg_module/gprf[326] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19911_  (.CLK(clknet_leaf_152_clk),
    .D(\reg_module/_00327_ ),
    .Q(\reg_module/gprf[327] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19912_  (.CLK(clknet_leaf_136_clk),
    .D(\reg_module/_00328_ ),
    .Q(\reg_module/gprf[328] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19913_  (.CLK(clknet_leaf_136_clk),
    .D(\reg_module/_00329_ ),
    .Q(\reg_module/gprf[329] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19914_  (.CLK(clknet_leaf_108_clk),
    .D(\reg_module/_00330_ ),
    .Q(\reg_module/gprf[330] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19915_  (.CLK(clknet_leaf_139_clk),
    .D(\reg_module/_00331_ ),
    .Q(\reg_module/gprf[331] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19916_  (.CLK(clknet_leaf_111_clk),
    .D(\reg_module/_00332_ ),
    .Q(\reg_module/gprf[332] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19917_  (.CLK(clknet_leaf_111_clk),
    .D(\reg_module/_00333_ ),
    .Q(\reg_module/gprf[333] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19918_  (.CLK(clknet_leaf_96_clk),
    .D(\reg_module/_00334_ ),
    .Q(\reg_module/gprf[334] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19919_  (.CLK(clknet_leaf_96_clk),
    .D(\reg_module/_00335_ ),
    .Q(\reg_module/gprf[335] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19920_  (.CLK(clknet_leaf_95_clk),
    .D(\reg_module/_00336_ ),
    .Q(\reg_module/gprf[336] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19921_  (.CLK(clknet_leaf_112_clk),
    .D(\reg_module/_00337_ ),
    .Q(\reg_module/gprf[337] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19922_  (.CLK(clknet_leaf_82_clk),
    .D(\reg_module/_00338_ ),
    .Q(\reg_module/gprf[338] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19923_  (.CLK(clknet_leaf_80_clk),
    .D(\reg_module/_00339_ ),
    .Q(\reg_module/gprf[339] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19924_  (.CLK(clknet_leaf_69_clk),
    .D(\reg_module/_00340_ ),
    .Q(\reg_module/gprf[340] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19925_  (.CLK(clknet_leaf_69_clk),
    .D(\reg_module/_00341_ ),
    .Q(\reg_module/gprf[341] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19926_  (.CLK(clknet_leaf_66_clk),
    .D(\reg_module/_00342_ ),
    .Q(\reg_module/gprf[342] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19927_  (.CLK(clknet_leaf_66_clk),
    .D(\reg_module/_00343_ ),
    .Q(\reg_module/gprf[343] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19928_  (.CLK(clknet_leaf_6_clk),
    .D(\reg_module/_00344_ ),
    .Q(\reg_module/gprf[344] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19929_  (.CLK(clknet_leaf_6_clk),
    .D(\reg_module/_00345_ ),
    .Q(\reg_module/gprf[345] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19930_  (.CLK(clknet_leaf_8_clk),
    .D(\reg_module/_00346_ ),
    .Q(\reg_module/gprf[346] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19931_  (.CLK(clknet_leaf_4_clk),
    .D(\reg_module/_00347_ ),
    .Q(\reg_module/gprf[347] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19932_  (.CLK(clknet_leaf_206_clk),
    .D(\reg_module/_00348_ ),
    .Q(\reg_module/gprf[348] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19933_  (.CLK(clknet_leaf_206_clk),
    .D(\reg_module/_00349_ ),
    .Q(\reg_module/gprf[349] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19934_  (.CLK(clknet_leaf_206_clk),
    .D(\reg_module/_00350_ ),
    .Q(\reg_module/gprf[350] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19935_  (.CLK(clknet_leaf_207_clk),
    .D(\reg_module/_00351_ ),
    .Q(\reg_module/gprf[351] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19936_  (.CLK(clknet_leaf_189_clk),
    .D(\reg_module/_00352_ ),
    .Q(\reg_module/gprf[352] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19937_  (.CLK(clknet_leaf_182_clk),
    .D(\reg_module/_00353_ ),
    .Q(\reg_module/gprf[353] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19938_  (.CLK(clknet_leaf_185_clk),
    .D(\reg_module/_00354_ ),
    .Q(\reg_module/gprf[354] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19939_  (.CLK(clknet_leaf_164_clk),
    .D(\reg_module/_00355_ ),
    .Q(\reg_module/gprf[355] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19940_  (.CLK(clknet_leaf_154_clk),
    .D(\reg_module/_00356_ ),
    .Q(\reg_module/gprf[356] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19941_  (.CLK(clknet_leaf_155_clk),
    .D(\reg_module/_00357_ ),
    .Q(\reg_module/gprf[357] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19942_  (.CLK(clknet_leaf_150_clk),
    .D(\reg_module/_00358_ ),
    .Q(\reg_module/gprf[358] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19943_  (.CLK(clknet_leaf_150_clk),
    .D(\reg_module/_00359_ ),
    .Q(\reg_module/gprf[359] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19944_  (.CLK(clknet_leaf_140_clk),
    .D(\reg_module/_00360_ ),
    .Q(\reg_module/gprf[360] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19945_  (.CLK(clknet_leaf_140_clk),
    .D(\reg_module/_00361_ ),
    .Q(\reg_module/gprf[361] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19946_  (.CLK(clknet_leaf_141_clk),
    .D(\reg_module/_00362_ ),
    .Q(\reg_module/gprf[362] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19947_  (.CLK(clknet_leaf_141_clk),
    .D(\reg_module/_00363_ ),
    .Q(\reg_module/gprf[363] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19948_  (.CLK(clknet_leaf_97_clk),
    .D(\reg_module/_00364_ ),
    .Q(\reg_module/gprf[364] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19949_  (.CLK(clknet_leaf_97_clk),
    .D(\reg_module/_00365_ ),
    .Q(\reg_module/gprf[365] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19950_  (.CLK(clknet_leaf_97_clk),
    .D(\reg_module/_00366_ ),
    .Q(\reg_module/gprf[366] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19951_  (.CLK(clknet_leaf_98_clk),
    .D(\reg_module/_00367_ ),
    .Q(\reg_module/gprf[367] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19952_  (.CLK(clknet_leaf_98_clk),
    .D(\reg_module/_00368_ ),
    .Q(\reg_module/gprf[368] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19953_  (.CLK(clknet_leaf_98_clk),
    .D(\reg_module/_00369_ ),
    .Q(\reg_module/gprf[369] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19954_  (.CLK(clknet_leaf_78_clk),
    .D(\reg_module/_00370_ ),
    .Q(\reg_module/gprf[370] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19955_  (.CLK(clknet_leaf_78_clk),
    .D(\reg_module/_00371_ ),
    .Q(\reg_module/gprf[371] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19956_  (.CLK(clknet_leaf_69_clk),
    .D(\reg_module/_00372_ ),
    .Q(\reg_module/gprf[372] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19957_  (.CLK(clknet_leaf_68_clk),
    .D(\reg_module/_00373_ ),
    .Q(\reg_module/gprf[373] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19958_  (.CLK(clknet_leaf_65_clk),
    .D(\reg_module/_00374_ ),
    .Q(\reg_module/gprf[374] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19959_  (.CLK(clknet_leaf_65_clk),
    .D(\reg_module/_00375_ ),
    .Q(\reg_module/gprf[375] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19960_  (.CLK(clknet_leaf_6_clk),
    .D(\reg_module/_00376_ ),
    .Q(\reg_module/gprf[376] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19961_  (.CLK(clknet_leaf_5_clk),
    .D(\reg_module/_00377_ ),
    .Q(\reg_module/gprf[377] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19962_  (.CLK(clknet_leaf_5_clk),
    .D(\reg_module/_00378_ ),
    .Q(\reg_module/gprf[378] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19963_  (.CLK(clknet_leaf_5_clk),
    .D(\reg_module/_00379_ ),
    .Q(\reg_module/gprf[379] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19964_  (.CLK(clknet_leaf_206_clk),
    .D(\reg_module/_00380_ ),
    .Q(\reg_module/gprf[380] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19965_  (.CLK(clknet_leaf_205_clk),
    .D(\reg_module/_00381_ ),
    .Q(\reg_module/gprf[381] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19966_  (.CLK(clknet_leaf_219_clk),
    .D(\reg_module/_00382_ ),
    .Q(\reg_module/gprf[382] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19967_  (.CLK(clknet_leaf_219_clk),
    .D(\reg_module/_00383_ ),
    .Q(\reg_module/gprf[383] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19968_  (.CLK(clknet_leaf_176_clk),
    .D(\reg_module/_00384_ ),
    .Q(\reg_module/gprf[384] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19969_  (.CLK(clknet_leaf_175_clk),
    .D(\reg_module/_00385_ ),
    .Q(\reg_module/gprf[385] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19970_  (.CLK(clknet_leaf_172_clk),
    .D(\reg_module/_00386_ ),
    .Q(\reg_module/gprf[386] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19971_  (.CLK(clknet_leaf_171_clk),
    .D(\reg_module/_00387_ ),
    .Q(\reg_module/gprf[387] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19972_  (.CLK(clknet_leaf_171_clk),
    .D(\reg_module/_00388_ ),
    .Q(\reg_module/gprf[388] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19973_  (.CLK(clknet_leaf_171_clk),
    .D(\reg_module/_00389_ ),
    .Q(\reg_module/gprf[389] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19974_  (.CLK(clknet_leaf_186_clk),
    .D(\reg_module/_00390_ ),
    .Q(\reg_module/gprf[390] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19975_  (.CLK(clknet_leaf_134_clk),
    .D(\reg_module/_00391_ ),
    .Q(\reg_module/gprf[391] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19976_  (.CLK(clknet_leaf_133_clk),
    .D(\reg_module/_00392_ ),
    .Q(\reg_module/gprf[392] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19977_  (.CLK(clknet_leaf_133_clk),
    .D(\reg_module/_00393_ ),
    .Q(\reg_module/gprf[393] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19978_  (.CLK(clknet_leaf_131_clk),
    .D(\reg_module/_00394_ ),
    .Q(\reg_module/gprf[394] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19979_  (.CLK(clknet_leaf_130_clk),
    .D(\reg_module/_00395_ ),
    .Q(\reg_module/gprf[395] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19980_  (.CLK(clknet_leaf_114_clk),
    .D(\reg_module/_00396_ ),
    .Q(\reg_module/gprf[396] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19981_  (.CLK(clknet_leaf_113_clk),
    .D(\reg_module/_00397_ ),
    .Q(\reg_module/gprf[397] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19982_  (.CLK(clknet_leaf_83_clk),
    .D(\reg_module/_00398_ ),
    .Q(\reg_module/gprf[398] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19983_  (.CLK(clknet_leaf_113_clk),
    .D(\reg_module/_00399_ ),
    .Q(\reg_module/gprf[399] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19984_  (.CLK(clknet_leaf_83_clk),
    .D(\reg_module/_00400_ ),
    .Q(\reg_module/gprf[400] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19985_  (.CLK(clknet_leaf_83_clk),
    .D(\reg_module/_00401_ ),
    .Q(\reg_module/gprf[401] ));
 sky130_fd_sc_hd__dfxtp_2 \reg_module/_19986_  (.CLK(clknet_leaf_18_clk),
    .D(\reg_module/_00402_ ),
    .Q(\reg_module/gprf[402] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19987_  (.CLK(clknet_leaf_18_clk),
    .D(\reg_module/_00403_ ),
    .Q(\reg_module/gprf[403] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19988_  (.CLK(clknet_leaf_18_clk),
    .D(\reg_module/_00404_ ),
    .Q(\reg_module/gprf[404] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19989_  (.CLK(clknet_leaf_18_clk),
    .D(\reg_module/_00405_ ),
    .Q(\reg_module/gprf[405] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19990_  (.CLK(clknet_leaf_17_clk),
    .D(\reg_module/_00406_ ),
    .Q(\reg_module/gprf[406] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19991_  (.CLK(clknet_leaf_17_clk),
    .D(\reg_module/_00407_ ),
    .Q(\reg_module/gprf[407] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19992_  (.CLK(clknet_leaf_222_clk),
    .D(\reg_module/_00408_ ),
    .Q(\reg_module/gprf[408] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19993_  (.CLK(clknet_leaf_222_clk),
    .D(\reg_module/_00409_ ),
    .Q(\reg_module/gprf[409] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19994_  (.CLK(clknet_leaf_1_clk),
    .D(\reg_module/_00410_ ),
    .Q(\reg_module/gprf[410] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19995_  (.CLK(clknet_leaf_1_clk),
    .D(\reg_module/_00411_ ),
    .Q(\reg_module/gprf[411] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19996_  (.CLK(clknet_leaf_2_clk),
    .D(\reg_module/_00412_ ),
    .Q(\reg_module/gprf[412] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19997_  (.CLK(clknet_leaf_2_clk),
    .D(\reg_module/_00413_ ),
    .Q(\reg_module/gprf[413] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19998_  (.CLK(clknet_leaf_218_clk),
    .D(\reg_module/_00414_ ),
    .Q(\reg_module/gprf[414] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_19999_  (.CLK(clknet_leaf_218_clk),
    .D(\reg_module/_00415_ ),
    .Q(\reg_module/gprf[415] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20000_  (.CLK(clknet_leaf_179_clk),
    .D(\reg_module/_00416_ ),
    .Q(\reg_module/gprf[416] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20001_  (.CLK(clknet_leaf_177_clk),
    .D(\reg_module/_00417_ ),
    .Q(\reg_module/gprf[417] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20002_  (.CLK(clknet_leaf_173_clk),
    .D(\reg_module/_00418_ ),
    .Q(\reg_module/gprf[418] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20003_  (.CLK(clknet_leaf_168_clk),
    .D(\reg_module/_00419_ ),
    .Q(\reg_module/gprf[419] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20004_  (.CLK(clknet_leaf_168_clk),
    .D(\reg_module/_00420_ ),
    .Q(\reg_module/gprf[420] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20005_  (.CLK(clknet_leaf_168_clk),
    .D(\reg_module/_00421_ ),
    .Q(\reg_module/gprf[421] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20006_  (.CLK(clknet_leaf_187_clk),
    .D(\reg_module/_00422_ ),
    .Q(\reg_module/gprf[422] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20007_  (.CLK(clknet_leaf_187_clk),
    .D(\reg_module/_00423_ ),
    .Q(\reg_module/gprf[423] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20008_  (.CLK(clknet_leaf_132_clk),
    .D(\reg_module/_00424_ ),
    .Q(\reg_module/gprf[424] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20009_  (.CLK(clknet_leaf_131_clk),
    .D(\reg_module/_00425_ ),
    .Q(\reg_module/gprf[425] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20010_  (.CLK(clknet_leaf_131_clk),
    .D(\reg_module/_00426_ ),
    .Q(\reg_module/gprf[426] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20011_  (.CLK(clknet_leaf_125_clk),
    .D(\reg_module/_00427_ ),
    .Q(\reg_module/gprf[427] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20012_  (.CLK(clknet_leaf_115_clk),
    .D(\reg_module/_00428_ ),
    .Q(\reg_module/gprf[428] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20013_  (.CLK(clknet_leaf_81_clk),
    .D(\reg_module/_00429_ ),
    .Q(\reg_module/gprf[429] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20014_  (.CLK(clknet_leaf_82_clk),
    .D(\reg_module/_00430_ ),
    .Q(\reg_module/gprf[430] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20015_  (.CLK(clknet_leaf_82_clk),
    .D(\reg_module/_00431_ ),
    .Q(\reg_module/gprf[431] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20016_  (.CLK(clknet_leaf_82_clk),
    .D(\reg_module/_00432_ ),
    .Q(\reg_module/gprf[432] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20017_  (.CLK(clknet_leaf_81_clk),
    .D(\reg_module/_00433_ ),
    .Q(\reg_module/gprf[433] ));
 sky130_fd_sc_hd__dfxtp_2 \reg_module/_20018_  (.CLK(clknet_leaf_14_clk),
    .D(\reg_module/_00434_ ),
    .Q(\reg_module/gprf[434] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20019_  (.CLK(clknet_leaf_13_clk),
    .D(\reg_module/_00435_ ),
    .Q(\reg_module/gprf[435] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20020_  (.CLK(clknet_leaf_13_clk),
    .D(\reg_module/_00436_ ),
    .Q(\reg_module/gprf[436] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20021_  (.CLK(clknet_leaf_13_clk),
    .D(\reg_module/_00437_ ),
    .Q(\reg_module/gprf[437] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20022_  (.CLK(clknet_leaf_17_clk),
    .D(\reg_module/_00438_ ),
    .Q(\reg_module/gprf[438] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20023_  (.CLK(clknet_leaf_14_clk),
    .D(\reg_module/_00439_ ),
    .Q(\reg_module/gprf[439] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20024_  (.CLK(clknet_leaf_5_clk),
    .D(\reg_module/_00440_ ),
    .Q(\reg_module/gprf[440] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20025_  (.CLK(clknet_leaf_5_clk),
    .D(\reg_module/_00441_ ),
    .Q(\reg_module/gprf[441] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20026_  (.CLK(clknet_leaf_3_clk),
    .D(\reg_module/_00442_ ),
    .Q(\reg_module/gprf[442] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20027_  (.CLK(clknet_leaf_3_clk),
    .D(\reg_module/_00443_ ),
    .Q(\reg_module/gprf[443] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20028_  (.CLK(clknet_leaf_2_clk),
    .D(\reg_module/_00444_ ),
    .Q(\reg_module/gprf[444] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20029_  (.CLK(clknet_leaf_2_clk),
    .D(\reg_module/_00445_ ),
    .Q(\reg_module/gprf[445] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20030_  (.CLK(clknet_leaf_218_clk),
    .D(\reg_module/_00446_ ),
    .Q(\reg_module/gprf[446] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20031_  (.CLK(clknet_leaf_218_clk),
    .D(\reg_module/_00447_ ),
    .Q(\reg_module/gprf[447] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20032_  (.CLK(clknet_leaf_180_clk),
    .D(\reg_module/_00448_ ),
    .Q(\reg_module/gprf[448] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20033_  (.CLK(clknet_leaf_180_clk),
    .D(\reg_module/_00449_ ),
    .Q(\reg_module/gprf[449] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20034_  (.CLK(clknet_leaf_178_clk),
    .D(\reg_module/_00450_ ),
    .Q(\reg_module/gprf[450] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20035_  (.CLK(clknet_leaf_182_clk),
    .D(\reg_module/_00451_ ),
    .Q(\reg_module/gprf[451] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20036_  (.CLK(clknet_leaf_167_clk),
    .D(\reg_module/_00452_ ),
    .Q(\reg_module/gprf[452] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20037_  (.CLK(clknet_leaf_185_clk),
    .D(\reg_module/_00453_ ),
    .Q(\reg_module/gprf[453] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20038_  (.CLK(clknet_leaf_187_clk),
    .D(\reg_module/_00454_ ),
    .Q(\reg_module/gprf[454] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20039_  (.CLK(clknet_leaf_132_clk),
    .D(\reg_module/_00455_ ),
    .Q(\reg_module/gprf[455] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20040_  (.CLK(clknet_leaf_132_clk),
    .D(\reg_module/_00456_ ),
    .Q(\reg_module/gprf[456] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20041_  (.CLK(clknet_leaf_187_clk),
    .D(\reg_module/_00457_ ),
    .Q(\reg_module/gprf[457] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20042_  (.CLK(clknet_leaf_126_clk),
    .D(\reg_module/_00458_ ),
    .Q(\reg_module/gprf[458] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20043_  (.CLK(clknet_leaf_126_clk),
    .D(\reg_module/_00459_ ),
    .Q(\reg_module/gprf[459] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20044_  (.CLK(clknet_leaf_119_clk),
    .D(\reg_module/_00460_ ),
    .Q(\reg_module/gprf[460] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20045_  (.CLK(clknet_leaf_115_clk),
    .D(\reg_module/_00461_ ),
    .Q(\reg_module/gprf[461] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20046_  (.CLK(clknet_leaf_115_clk),
    .D(\reg_module/_00462_ ),
    .Q(\reg_module/gprf[462] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20047_  (.CLK(clknet_leaf_116_clk),
    .D(\reg_module/_00463_ ),
    .Q(\reg_module/gprf[463] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20048_  (.CLK(clknet_leaf_115_clk),
    .D(\reg_module/_00464_ ),
    .Q(\reg_module/gprf[464] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20049_  (.CLK(clknet_leaf_115_clk),
    .D(\reg_module/_00465_ ),
    .Q(\reg_module/gprf[465] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20050_  (.CLK(clknet_leaf_120_clk),
    .D(\reg_module/_00466_ ),
    .Q(\reg_module/gprf[466] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20051_  (.CLK(clknet_leaf_120_clk),
    .D(\reg_module/_00467_ ),
    .Q(\reg_module/gprf[467] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20052_  (.CLK(clknet_leaf_13_clk),
    .D(\reg_module/_00468_ ),
    .Q(\reg_module/gprf[468] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20053_  (.CLK(clknet_leaf_13_clk),
    .D(\reg_module/_00469_ ),
    .Q(\reg_module/gprf[469] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20054_  (.CLK(clknet_leaf_15_clk),
    .D(\reg_module/_00470_ ),
    .Q(\reg_module/gprf[470] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20055_  (.CLK(clknet_leaf_15_clk),
    .D(\reg_module/_00471_ ),
    .Q(\reg_module/gprf[471] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20056_  (.CLK(clknet_leaf_15_clk),
    .D(\reg_module/_00472_ ),
    .Q(\reg_module/gprf[472] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20057_  (.CLK(clknet_leaf_15_clk),
    .D(\reg_module/_00473_ ),
    .Q(\reg_module/gprf[473] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20058_  (.CLK(clknet_leaf_4_clk),
    .D(\reg_module/_00474_ ),
    .Q(\reg_module/gprf[474] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20059_  (.CLK(clknet_leaf_4_clk),
    .D(\reg_module/_00475_ ),
    .Q(\reg_module/gprf[475] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20060_  (.CLK(clknet_leaf_206_clk),
    .D(\reg_module/_00476_ ),
    .Q(\reg_module/gprf[476] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20061_  (.CLK(clknet_leaf_206_clk),
    .D(\reg_module/_00477_ ),
    .Q(\reg_module/gprf[477] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20062_  (.CLK(clknet_leaf_219_clk),
    .D(\reg_module/_00478_ ),
    .Q(\reg_module/gprf[478] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20063_  (.CLK(clknet_leaf_218_clk),
    .D(\reg_module/_00479_ ),
    .Q(\reg_module/gprf[479] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20064_  (.CLK(clknet_leaf_180_clk),
    .D(\reg_module/_00480_ ),
    .Q(\reg_module/gprf[480] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20065_  (.CLK(clknet_leaf_181_clk),
    .D(\reg_module/_00481_ ),
    .Q(\reg_module/gprf[481] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20066_  (.CLK(clknet_leaf_182_clk),
    .D(\reg_module/_00482_ ),
    .Q(\reg_module/gprf[482] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20067_  (.CLK(clknet_leaf_182_clk),
    .D(\reg_module/_00483_ ),
    .Q(\reg_module/gprf[483] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20068_  (.CLK(clknet_leaf_184_clk),
    .D(\reg_module/_00484_ ),
    .Q(\reg_module/gprf[484] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20069_  (.CLK(clknet_leaf_184_clk),
    .D(\reg_module/_00485_ ),
    .Q(\reg_module/gprf[485] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20070_  (.CLK(clknet_leaf_187_clk),
    .D(\reg_module/_00486_ ),
    .Q(\reg_module/gprf[486] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20071_  (.CLK(clknet_leaf_188_clk),
    .D(\reg_module/_00487_ ),
    .Q(\reg_module/gprf[487] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20072_  (.CLK(clknet_leaf_188_clk),
    .D(\reg_module/_00488_ ),
    .Q(\reg_module/gprf[488] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20073_  (.CLK(clknet_leaf_193_clk),
    .D(\reg_module/_00489_ ),
    .Q(\reg_module/gprf[489] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20074_  (.CLK(clknet_leaf_125_clk),
    .D(\reg_module/_00490_ ),
    .Q(\reg_module/gprf[490] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20075_  (.CLK(clknet_leaf_125_clk),
    .D(\reg_module/_00491_ ),
    .Q(\reg_module/gprf[491] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20076_  (.CLK(clknet_leaf_119_clk),
    .D(\reg_module/_00492_ ),
    .Q(\reg_module/gprf[492] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20077_  (.CLK(clknet_leaf_119_clk),
    .D(\reg_module/_00493_ ),
    .Q(\reg_module/gprf[493] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20078_  (.CLK(clknet_leaf_119_clk),
    .D(\reg_module/_00494_ ),
    .Q(\reg_module/gprf[494] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20079_  (.CLK(clknet_leaf_115_clk),
    .D(\reg_module/_00495_ ),
    .Q(\reg_module/gprf[495] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20080_  (.CLK(clknet_leaf_115_clk),
    .D(\reg_module/_00496_ ),
    .Q(\reg_module/gprf[496] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20081_  (.CLK(clknet_leaf_120_clk),
    .D(\reg_module/_00497_ ),
    .Q(\reg_module/gprf[497] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20082_  (.CLK(clknet_leaf_120_clk),
    .D(\reg_module/_00498_ ),
    .Q(\reg_module/gprf[498] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20083_  (.CLK(clknet_leaf_120_clk),
    .D(\reg_module/_00499_ ),
    .Q(\reg_module/gprf[499] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20084_  (.CLK(clknet_leaf_14_clk),
    .D(\reg_module/_00500_ ),
    .Q(\reg_module/gprf[500] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20085_  (.CLK(clknet_leaf_15_clk),
    .D(\reg_module/_00501_ ),
    .Q(\reg_module/gprf[501] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20086_  (.CLK(clknet_leaf_17_clk),
    .D(\reg_module/_00502_ ),
    .Q(\reg_module/gprf[502] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20087_  (.CLK(clknet_leaf_16_clk),
    .D(\reg_module/_00503_ ),
    .Q(\reg_module/gprf[503] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20088_  (.CLK(clknet_leaf_16_clk),
    .D(\reg_module/_00504_ ),
    .Q(\reg_module/gprf[504] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20089_  (.CLK(clknet_leaf_15_clk),
    .D(\reg_module/_00505_ ),
    .Q(\reg_module/gprf[505] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20090_  (.CLK(clknet_leaf_3_clk),
    .D(\reg_module/_00506_ ),
    .Q(\reg_module/gprf[506] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20091_  (.CLK(clknet_leaf_3_clk),
    .D(\reg_module/_00507_ ),
    .Q(\reg_module/gprf[507] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20092_  (.CLK(clknet_leaf_205_clk),
    .D(\reg_module/_00508_ ),
    .Q(\reg_module/gprf[508] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20093_  (.CLK(clknet_leaf_2_clk),
    .D(\reg_module/_00509_ ),
    .Q(\reg_module/gprf[509] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20094_  (.CLK(clknet_leaf_219_clk),
    .D(\reg_module/_00510_ ),
    .Q(\reg_module/gprf[510] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20095_  (.CLK(clknet_leaf_208_clk),
    .D(\reg_module/_00511_ ),
    .Q(\reg_module/gprf[511] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20096_  (.CLK(clknet_leaf_161_clk),
    .D(\reg_module/_00512_ ),
    .Q(\reg_module/gprf[512] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20097_  (.CLK(clknet_leaf_161_clk),
    .D(\reg_module/_00513_ ),
    .Q(\reg_module/gprf[513] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20098_  (.CLK(clknet_leaf_161_clk),
    .D(\reg_module/_00514_ ),
    .Q(\reg_module/gprf[514] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20099_  (.CLK(clknet_leaf_161_clk),
    .D(\reg_module/_00515_ ),
    .Q(\reg_module/gprf[515] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20100_  (.CLK(clknet_leaf_161_clk),
    .D(\reg_module/_00516_ ),
    .Q(\reg_module/gprf[516] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20101_  (.CLK(clknet_leaf_161_clk),
    .D(\reg_module/_00517_ ),
    .Q(\reg_module/gprf[517] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20102_  (.CLK(clknet_leaf_147_clk),
    .D(\reg_module/_00518_ ),
    .Q(\reg_module/gprf[518] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20103_  (.CLK(clknet_leaf_147_clk),
    .D(\reg_module/_00519_ ),
    .Q(\reg_module/gprf[519] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20104_  (.CLK(clknet_leaf_147_clk),
    .D(\reg_module/_00520_ ),
    .Q(\reg_module/gprf[520] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20105_  (.CLK(clknet_leaf_146_clk),
    .D(\reg_module/_00521_ ),
    .Q(\reg_module/gprf[521] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20106_  (.CLK(clknet_leaf_145_clk),
    .D(\reg_module/_00522_ ),
    .Q(\reg_module/gprf[522] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20107_  (.CLK(clknet_leaf_146_clk),
    .D(\reg_module/_00523_ ),
    .Q(\reg_module/gprf[523] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20108_  (.CLK(clknet_leaf_97_clk),
    .D(\reg_module/_00524_ ),
    .Q(\reg_module/gprf[524] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20109_  (.CLK(clknet_leaf_97_clk),
    .D(\reg_module/_00525_ ),
    .Q(\reg_module/gprf[525] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20110_  (.CLK(clknet_leaf_97_clk),
    .D(\reg_module/_00526_ ),
    .Q(\reg_module/gprf[526] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20111_  (.CLK(clknet_leaf_97_clk),
    .D(\reg_module/_00527_ ),
    .Q(\reg_module/gprf[527] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20112_  (.CLK(clknet_leaf_101_clk),
    .D(\reg_module/_00528_ ),
    .Q(\reg_module/gprf[528] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20113_  (.CLK(clknet_leaf_98_clk),
    .D(\reg_module/_00529_ ),
    .Q(\reg_module/gprf[529] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20114_  (.CLK(clknet_leaf_13_clk),
    .D(\reg_module/_00530_ ),
    .Q(\reg_module/gprf[530] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20115_  (.CLK(clknet_leaf_71_clk),
    .D(\reg_module/_00531_ ),
    .Q(\reg_module/gprf[531] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20116_  (.CLK(clknet_leaf_66_clk),
    .D(\reg_module/_00532_ ),
    .Q(\reg_module/gprf[532] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20117_  (.CLK(clknet_leaf_71_clk),
    .D(\reg_module/_00533_ ),
    .Q(\reg_module/gprf[533] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20118_  (.CLK(clknet_leaf_13_clk),
    .D(\reg_module/_00534_ ),
    .Q(\reg_module/gprf[534] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20119_  (.CLK(clknet_leaf_66_clk),
    .D(\reg_module/_00535_ ),
    .Q(\reg_module/gprf[535] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20120_  (.CLK(clknet_leaf_200_clk),
    .D(\reg_module/_00536_ ),
    .Q(\reg_module/gprf[536] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20121_  (.CLK(clknet_leaf_200_clk),
    .D(\reg_module/_00537_ ),
    .Q(\reg_module/gprf[537] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20122_  (.CLK(clknet_leaf_200_clk),
    .D(\reg_module/_00538_ ),
    .Q(\reg_module/gprf[538] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20123_  (.CLK(clknet_leaf_201_clk),
    .D(\reg_module/_00539_ ),
    .Q(\reg_module/gprf[539] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20124_  (.CLK(clknet_leaf_200_clk),
    .D(\reg_module/_00540_ ),
    .Q(\reg_module/gprf[540] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20125_  (.CLK(clknet_leaf_200_clk),
    .D(\reg_module/_00541_ ),
    .Q(\reg_module/gprf[541] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20126_  (.CLK(clknet_leaf_214_clk),
    .D(\reg_module/_00542_ ),
    .Q(\reg_module/gprf[542] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20127_  (.CLK(clknet_leaf_215_clk),
    .D(\reg_module/_00543_ ),
    .Q(\reg_module/gprf[543] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20128_  (.CLK(clknet_leaf_174_clk),
    .D(\reg_module/_00544_ ),
    .Q(\reg_module/gprf[544] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20129_  (.CLK(clknet_leaf_173_clk),
    .D(\reg_module/_00545_ ),
    .Q(\reg_module/gprf[545] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20130_  (.CLK(clknet_leaf_173_clk),
    .D(\reg_module/_00546_ ),
    .Q(\reg_module/gprf[546] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20131_  (.CLK(clknet_leaf_168_clk),
    .D(\reg_module/_00547_ ),
    .Q(\reg_module/gprf[547] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20132_  (.CLK(clknet_leaf_163_clk),
    .D(\reg_module/_00548_ ),
    .Q(\reg_module/gprf[548] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20133_  (.CLK(clknet_leaf_163_clk),
    .D(\reg_module/_00549_ ),
    .Q(\reg_module/gprf[549] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20134_  (.CLK(clknet_leaf_150_clk),
    .D(\reg_module/_00550_ ),
    .Q(\reg_module/gprf[550] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20135_  (.CLK(clknet_leaf_150_clk),
    .D(\reg_module/_00551_ ),
    .Q(\reg_module/gprf[551] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20136_  (.CLK(clknet_leaf_151_clk),
    .D(\reg_module/_00552_ ),
    .Q(\reg_module/gprf[552] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20137_  (.CLK(clknet_leaf_147_clk),
    .D(\reg_module/_00553_ ),
    .Q(\reg_module/gprf[553] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20138_  (.CLK(clknet_leaf_141_clk),
    .D(\reg_module/_00554_ ),
    .Q(\reg_module/gprf[554] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20139_  (.CLK(clknet_leaf_141_clk),
    .D(\reg_module/_00555_ ),
    .Q(\reg_module/gprf[555] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20140_  (.CLK(clknet_leaf_98_clk),
    .D(\reg_module/_00556_ ),
    .Q(\reg_module/gprf[556] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20141_  (.CLK(clknet_leaf_98_clk),
    .D(\reg_module/_00557_ ),
    .Q(\reg_module/gprf[557] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20142_  (.CLK(clknet_leaf_98_clk),
    .D(\reg_module/_00558_ ),
    .Q(\reg_module/gprf[558] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20143_  (.CLK(clknet_leaf_98_clk),
    .D(\reg_module/_00559_ ),
    .Q(\reg_module/gprf[559] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20144_  (.CLK(clknet_leaf_98_clk),
    .D(\reg_module/_00560_ ),
    .Q(\reg_module/gprf[560] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20145_  (.CLK(clknet_leaf_98_clk),
    .D(\reg_module/_00561_ ),
    .Q(\reg_module/gprf[561] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20146_  (.CLK(clknet_leaf_78_clk),
    .D(\reg_module/_00562_ ),
    .Q(\reg_module/gprf[562] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20147_  (.CLK(clknet_leaf_78_clk),
    .D(\reg_module/_00563_ ),
    .Q(\reg_module/gprf[563] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20148_  (.CLK(clknet_leaf_78_clk),
    .D(\reg_module/_00564_ ),
    .Q(\reg_module/gprf[564] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20149_  (.CLK(clknet_leaf_68_clk),
    .D(\reg_module/_00565_ ),
    .Q(\reg_module/gprf[565] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20150_  (.CLK(clknet_leaf_67_clk),
    .D(\reg_module/_00566_ ),
    .Q(\reg_module/gprf[566] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20151_  (.CLK(clknet_leaf_66_clk),
    .D(\reg_module/_00567_ ),
    .Q(\reg_module/gprf[567] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20152_  (.CLK(clknet_leaf_9_clk),
    .D(\reg_module/_00568_ ),
    .Q(\reg_module/gprf[568] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20153_  (.CLK(clknet_leaf_198_clk),
    .D(\reg_module/_00569_ ),
    .Q(\reg_module/gprf[569] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20154_  (.CLK(clknet_leaf_198_clk),
    .D(\reg_module/_00570_ ),
    .Q(\reg_module/gprf[570] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20155_  (.CLK(clknet_leaf_199_clk),
    .D(\reg_module/_00571_ ),
    .Q(\reg_module/gprf[571] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20156_  (.CLK(clknet_leaf_202_clk),
    .D(\reg_module/_00572_ ),
    .Q(\reg_module/gprf[572] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20157_  (.CLK(clknet_leaf_202_clk),
    .D(\reg_module/_00573_ ),
    .Q(\reg_module/gprf[573] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20158_  (.CLK(clknet_leaf_214_clk),
    .D(\reg_module/_00574_ ),
    .Q(\reg_module/gprf[574] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20159_  (.CLK(clknet_leaf_212_clk),
    .D(\reg_module/_00575_ ),
    .Q(\reg_module/gprf[575] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20160_  (.CLK(clknet_leaf_177_clk),
    .D(\reg_module/_00576_ ),
    .Q(\reg_module/gprf[576] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20161_  (.CLK(clknet_leaf_180_clk),
    .D(\reg_module/_00577_ ),
    .Q(\reg_module/gprf[577] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20162_  (.CLK(clknet_leaf_169_clk),
    .D(\reg_module/_00578_ ),
    .Q(\reg_module/gprf[578] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20163_  (.CLK(clknet_leaf_164_clk),
    .D(\reg_module/_00579_ ),
    .Q(\reg_module/gprf[579] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20164_  (.CLK(clknet_leaf_155_clk),
    .D(\reg_module/_00580_ ),
    .Q(\reg_module/gprf[580] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20165_  (.CLK(clknet_leaf_155_clk),
    .D(\reg_module/_00581_ ),
    .Q(\reg_module/gprf[581] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20166_  (.CLK(clknet_leaf_148_clk),
    .D(\reg_module/_00582_ ),
    .Q(\reg_module/gprf[582] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20167_  (.CLK(clknet_leaf_148_clk),
    .D(\reg_module/_00583_ ),
    .Q(\reg_module/gprf[583] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20168_  (.CLK(clknet_leaf_144_clk),
    .D(\reg_module/_00584_ ),
    .Q(\reg_module/gprf[584] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20169_  (.CLK(clknet_leaf_145_clk),
    .D(\reg_module/_00585_ ),
    .Q(\reg_module/gprf[585] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20170_  (.CLK(clknet_leaf_144_clk),
    .D(\reg_module/_00586_ ),
    .Q(\reg_module/gprf[586] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20171_  (.CLK(clknet_leaf_144_clk),
    .D(\reg_module/_00587_ ),
    .Q(\reg_module/gprf[587] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20172_  (.CLK(clknet_leaf_106_clk),
    .D(\reg_module/_00588_ ),
    .Q(\reg_module/gprf[588] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20173_  (.CLK(clknet_leaf_106_clk),
    .D(\reg_module/_00589_ ),
    .Q(\reg_module/gprf[589] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20174_  (.CLK(clknet_leaf_103_clk),
    .D(\reg_module/_00590_ ),
    .Q(\reg_module/gprf[590] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20175_  (.CLK(clknet_leaf_103_clk),
    .D(\reg_module/_00591_ ),
    .Q(\reg_module/gprf[591] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20176_  (.CLK(clknet_leaf_103_clk),
    .D(\reg_module/_00592_ ),
    .Q(\reg_module/gprf[592] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20177_  (.CLK(clknet_leaf_102_clk),
    .D(\reg_module/_00593_ ),
    .Q(\reg_module/gprf[593] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20178_  (.CLK(clknet_leaf_75_clk),
    .D(\reg_module/_00594_ ),
    .Q(\reg_module/gprf[594] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20179_  (.CLK(clknet_leaf_75_clk),
    .D(\reg_module/_00595_ ),
    .Q(\reg_module/gprf[595] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20180_  (.CLK(clknet_leaf_74_clk),
    .D(\reg_module/_00596_ ),
    .Q(\reg_module/gprf[596] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20181_  (.CLK(clknet_leaf_13_clk),
    .D(\reg_module/_00597_ ),
    .Q(\reg_module/gprf[597] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20182_  (.CLK(clknet_leaf_13_clk),
    .D(\reg_module/_00598_ ),
    .Q(\reg_module/gprf[598] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20183_  (.CLK(clknet_leaf_71_clk),
    .D(\reg_module/_00599_ ),
    .Q(\reg_module/gprf[599] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20184_  (.CLK(clknet_leaf_10_clk),
    .D(\reg_module/_00600_ ),
    .Q(\reg_module/gprf[600] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20185_  (.CLK(clknet_leaf_9_clk),
    .D(\reg_module/_00601_ ),
    .Q(\reg_module/gprf[601] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20186_  (.CLK(clknet_leaf_199_clk),
    .D(\reg_module/_00602_ ),
    .Q(\reg_module/gprf[602] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20187_  (.CLK(clknet_leaf_203_clk),
    .D(\reg_module/_00603_ ),
    .Q(\reg_module/gprf[603] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20188_  (.CLK(clknet_leaf_209_clk),
    .D(\reg_module/_00604_ ),
    .Q(\reg_module/gprf[604] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20189_  (.CLK(clknet_leaf_209_clk),
    .D(\reg_module/_00605_ ),
    .Q(\reg_module/gprf[605] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20190_  (.CLK(clknet_leaf_213_clk),
    .D(\reg_module/_00606_ ),
    .Q(\reg_module/gprf[606] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20191_  (.CLK(clknet_leaf_213_clk),
    .D(\reg_module/_00607_ ),
    .Q(\reg_module/gprf[607] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20192_  (.CLK(clknet_leaf_178_clk),
    .D(\reg_module/_00608_ ),
    .Q(\reg_module/gprf[608] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20193_  (.CLK(clknet_leaf_178_clk),
    .D(\reg_module/_00609_ ),
    .Q(\reg_module/gprf[609] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20194_  (.CLK(clknet_leaf_167_clk),
    .D(\reg_module/_00610_ ),
    .Q(\reg_module/gprf[610] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20195_  (.CLK(clknet_leaf_164_clk),
    .D(\reg_module/_00611_ ),
    .Q(\reg_module/gprf[611] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20196_  (.CLK(clknet_leaf_163_clk),
    .D(\reg_module/_00612_ ),
    .Q(\reg_module/gprf[612] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20197_  (.CLK(clknet_leaf_163_clk),
    .D(\reg_module/_00613_ ),
    .Q(\reg_module/gprf[613] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20198_  (.CLK(clknet_leaf_150_clk),
    .D(\reg_module/_00614_ ),
    .Q(\reg_module/gprf[614] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20199_  (.CLK(clknet_leaf_151_clk),
    .D(\reg_module/_00615_ ),
    .Q(\reg_module/gprf[615] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20200_  (.CLK(clknet_leaf_146_clk),
    .D(\reg_module/_00616_ ),
    .Q(\reg_module/gprf[616] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20201_  (.CLK(clknet_leaf_140_clk),
    .D(\reg_module/_00617_ ),
    .Q(\reg_module/gprf[617] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20202_  (.CLK(clknet_leaf_140_clk),
    .D(\reg_module/_00618_ ),
    .Q(\reg_module/gprf[618] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20203_  (.CLK(clknet_leaf_140_clk),
    .D(\reg_module/_00619_ ),
    .Q(\reg_module/gprf[619] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20204_  (.CLK(clknet_leaf_108_clk),
    .D(\reg_module/_00620_ ),
    .Q(\reg_module/gprf[620] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20205_  (.CLK(clknet_leaf_106_clk),
    .D(\reg_module/_00621_ ),
    .Q(\reg_module/gprf[621] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20206_  (.CLK(clknet_leaf_107_clk),
    .D(\reg_module/_00622_ ),
    .Q(\reg_module/gprf[622] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20207_  (.CLK(clknet_leaf_107_clk),
    .D(\reg_module/_00623_ ),
    .Q(\reg_module/gprf[623] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20208_  (.CLK(clknet_leaf_107_clk),
    .D(\reg_module/_00624_ ),
    .Q(\reg_module/gprf[624] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20209_  (.CLK(clknet_leaf_102_clk),
    .D(\reg_module/_00625_ ),
    .Q(\reg_module/gprf[625] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20210_  (.CLK(clknet_leaf_76_clk),
    .D(\reg_module/_00626_ ),
    .Q(\reg_module/gprf[626] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20211_  (.CLK(clknet_leaf_76_clk),
    .D(\reg_module/_00627_ ),
    .Q(\reg_module/gprf[627] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20212_  (.CLK(clknet_leaf_77_clk),
    .D(\reg_module/_00628_ ),
    .Q(\reg_module/gprf[628] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20213_  (.CLK(clknet_leaf_70_clk),
    .D(\reg_module/_00629_ ),
    .Q(\reg_module/gprf[629] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20214_  (.CLK(clknet_leaf_70_clk),
    .D(\reg_module/_00630_ ),
    .Q(\reg_module/gprf[630] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20215_  (.CLK(clknet_leaf_70_clk),
    .D(\reg_module/_00631_ ),
    .Q(\reg_module/gprf[631] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20216_  (.CLK(clknet_leaf_10_clk),
    .D(\reg_module/_00632_ ),
    .Q(\reg_module/gprf[632] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20217_  (.CLK(clknet_leaf_10_clk),
    .D(\reg_module/_00633_ ),
    .Q(\reg_module/gprf[633] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20218_  (.CLK(clknet_leaf_200_clk),
    .D(\reg_module/_00634_ ),
    .Q(\reg_module/gprf[634] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20219_  (.CLK(clknet_leaf_201_clk),
    .D(\reg_module/_00635_ ),
    .Q(\reg_module/gprf[635] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20220_  (.CLK(clknet_leaf_209_clk),
    .D(\reg_module/_00636_ ),
    .Q(\reg_module/gprf[636] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20221_  (.CLK(clknet_leaf_202_clk),
    .D(\reg_module/_00637_ ),
    .Q(\reg_module/gprf[637] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20222_  (.CLK(clknet_leaf_213_clk),
    .D(\reg_module/_00638_ ),
    .Q(\reg_module/gprf[638] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20223_  (.CLK(clknet_leaf_212_clk),
    .D(\reg_module/_00639_ ),
    .Q(\reg_module/gprf[639] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20224_  (.CLK(clknet_leaf_176_clk),
    .D(\reg_module/_00640_ ),
    .Q(\reg_module/gprf[640] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20225_  (.CLK(clknet_leaf_171_clk),
    .D(\reg_module/_00641_ ),
    .Q(\reg_module/gprf[641] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20226_  (.CLK(clknet_leaf_171_clk),
    .D(\reg_module/_00642_ ),
    .Q(\reg_module/gprf[642] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20227_  (.CLK(clknet_leaf_161_clk),
    .D(\reg_module/_00643_ ),
    .Q(\reg_module/gprf[643] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20228_  (.CLK(clknet_leaf_170_clk),
    .D(\reg_module/_00644_ ),
    .Q(\reg_module/gprf[644] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20229_  (.CLK(clknet_leaf_170_clk),
    .D(\reg_module/_00645_ ),
    .Q(\reg_module/gprf[645] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20230_  (.CLK(clknet_leaf_166_clk),
    .D(\reg_module/_00646_ ),
    .Q(\reg_module/gprf[646] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20231_  (.CLK(clknet_leaf_186_clk),
    .D(\reg_module/_00647_ ),
    .Q(\reg_module/gprf[647] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20232_  (.CLK(clknet_leaf_133_clk),
    .D(\reg_module/_00648_ ),
    .Q(\reg_module/gprf[648] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20233_  (.CLK(clknet_leaf_130_clk),
    .D(\reg_module/_00649_ ),
    .Q(\reg_module/gprf[649] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20234_  (.CLK(clknet_leaf_137_clk),
    .D(\reg_module/_00650_ ),
    .Q(\reg_module/gprf[650] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20235_  (.CLK(clknet_leaf_127_clk),
    .D(\reg_module/_00651_ ),
    .Q(\reg_module/gprf[651] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20236_  (.CLK(clknet_leaf_128_clk),
    .D(\reg_module/_00652_ ),
    .Q(\reg_module/gprf[652] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20237_  (.CLK(clknet_leaf_138_clk),
    .D(\reg_module/_00653_ ),
    .Q(\reg_module/gprf[653] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20238_  (.CLK(clknet_leaf_127_clk),
    .D(\reg_module/_00654_ ),
    .Q(\reg_module/gprf[654] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20239_  (.CLK(clknet_leaf_128_clk),
    .D(\reg_module/_00655_ ),
    .Q(\reg_module/gprf[655] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20240_  (.CLK(clknet_leaf_126_clk),
    .D(\reg_module/_00656_ ),
    .Q(\reg_module/gprf[656] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20241_  (.CLK(clknet_leaf_126_clk),
    .D(\reg_module/_00657_ ),
    .Q(\reg_module/gprf[657] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20242_  (.CLK(clknet_leaf_126_clk),
    .D(\reg_module/_00658_ ),
    .Q(\reg_module/gprf[658] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20243_  (.CLK(clknet_leaf_124_clk),
    .D(\reg_module/_00659_ ),
    .Q(\reg_module/gprf[659] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20244_  (.CLK(clknet_leaf_123_clk),
    .D(\reg_module/_00660_ ),
    .Q(\reg_module/gprf[660] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20245_  (.CLK(clknet_leaf_123_clk),
    .D(\reg_module/_00661_ ),
    .Q(\reg_module/gprf[661] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20246_  (.CLK(clknet_leaf_195_clk),
    .D(\reg_module/_00662_ ),
    .Q(\reg_module/gprf[662] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20247_  (.CLK(clknet_leaf_192_clk),
    .D(\reg_module/_00663_ ),
    .Q(\reg_module/gprf[663] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20248_  (.CLK(clknet_leaf_9_clk),
    .D(\reg_module/_00664_ ),
    .Q(\reg_module/gprf[664] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20249_  (.CLK(clknet_leaf_9_clk),
    .D(\reg_module/_00665_ ),
    .Q(\reg_module/gprf[665] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20250_  (.CLK(clknet_leaf_9_clk),
    .D(\reg_module/_00666_ ),
    .Q(\reg_module/gprf[666] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20251_  (.CLK(clknet_leaf_199_clk),
    .D(\reg_module/_00667_ ),
    .Q(\reg_module/gprf[667] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20252_  (.CLK(clknet_leaf_209_clk),
    .D(\reg_module/_00668_ ),
    .Q(\reg_module/gprf[668] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20253_  (.CLK(clknet_leaf_209_clk),
    .D(\reg_module/_00669_ ),
    .Q(\reg_module/gprf[669] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20254_  (.CLK(clknet_leaf_216_clk),
    .D(\reg_module/_00670_ ),
    .Q(\reg_module/gprf[670] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20255_  (.CLK(clknet_leaf_216_clk),
    .D(\reg_module/_00671_ ),
    .Q(\reg_module/gprf[671] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20256_  (.CLK(clknet_leaf_176_clk),
    .D(\reg_module/_00672_ ),
    .Q(\reg_module/gprf[672] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20257_  (.CLK(clknet_leaf_174_clk),
    .D(\reg_module/_00673_ ),
    .Q(\reg_module/gprf[673] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20258_  (.CLK(clknet_leaf_173_clk),
    .D(\reg_module/_00674_ ),
    .Q(\reg_module/gprf[674] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20259_  (.CLK(clknet_leaf_169_clk),
    .D(\reg_module/_00675_ ),
    .Q(\reg_module/gprf[675] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20260_  (.CLK(clknet_leaf_169_clk),
    .D(\reg_module/_00676_ ),
    .Q(\reg_module/gprf[676] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20261_  (.CLK(clknet_leaf_169_clk),
    .D(\reg_module/_00677_ ),
    .Q(\reg_module/gprf[677] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20262_  (.CLK(clknet_leaf_186_clk),
    .D(\reg_module/_00678_ ),
    .Q(\reg_module/gprf[678] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20263_  (.CLK(clknet_leaf_186_clk),
    .D(\reg_module/_00679_ ),
    .Q(\reg_module/gprf[679] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20264_  (.CLK(clknet_leaf_186_clk),
    .D(\reg_module/_00680_ ),
    .Q(\reg_module/gprf[680] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20265_  (.CLK(clknet_leaf_134_clk),
    .D(\reg_module/_00681_ ),
    .Q(\reg_module/gprf[681] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20266_  (.CLK(clknet_leaf_130_clk),
    .D(\reg_module/_00682_ ),
    .Q(\reg_module/gprf[682] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20267_  (.CLK(clknet_leaf_131_clk),
    .D(\reg_module/_00683_ ),
    .Q(\reg_module/gprf[683] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20268_  (.CLK(clknet_leaf_127_clk),
    .D(\reg_module/_00684_ ),
    .Q(\reg_module/gprf[684] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20269_  (.CLK(clknet_leaf_127_clk),
    .D(\reg_module/_00685_ ),
    .Q(\reg_module/gprf[685] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20270_  (.CLK(clknet_leaf_117_clk),
    .D(\reg_module/_00686_ ),
    .Q(\reg_module/gprf[686] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20271_  (.CLK(clknet_leaf_118_clk),
    .D(\reg_module/_00687_ ),
    .Q(\reg_module/gprf[687] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20272_  (.CLK(clknet_leaf_126_clk),
    .D(\reg_module/_00688_ ),
    .Q(\reg_module/gprf[688] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20273_  (.CLK(clknet_leaf_126_clk),
    .D(\reg_module/_00689_ ),
    .Q(\reg_module/gprf[689] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20274_  (.CLK(clknet_leaf_126_clk),
    .D(\reg_module/_00690_ ),
    .Q(\reg_module/gprf[690] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20275_  (.CLK(clknet_leaf_123_clk),
    .D(\reg_module/_00691_ ),
    .Q(\reg_module/gprf[691] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20276_  (.CLK(clknet_leaf_123_clk),
    .D(\reg_module/_00692_ ),
    .Q(\reg_module/gprf[692] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20277_  (.CLK(clknet_leaf_123_clk),
    .D(\reg_module/_00693_ ),
    .Q(\reg_module/gprf[693] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20278_  (.CLK(clknet_leaf_196_clk),
    .D(\reg_module/_00694_ ),
    .Q(\reg_module/gprf[694] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20279_  (.CLK(clknet_leaf_11_clk),
    .D(\reg_module/_00695_ ),
    .Q(\reg_module/gprf[695] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20280_  (.CLK(clknet_leaf_7_clk),
    .D(\reg_module/_00696_ ),
    .Q(\reg_module/gprf[696] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20281_  (.CLK(clknet_leaf_7_clk),
    .D(\reg_module/_00697_ ),
    .Q(\reg_module/gprf[697] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20282_  (.CLK(clknet_leaf_8_clk),
    .D(\reg_module/_00698_ ),
    .Q(\reg_module/gprf[698] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20283_  (.CLK(clknet_leaf_203_clk),
    .D(\reg_module/_00699_ ),
    .Q(\reg_module/gprf[699] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20284_  (.CLK(clknet_leaf_204_clk),
    .D(\reg_module/_00700_ ),
    .Q(\reg_module/gprf[700] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20285_  (.CLK(clknet_leaf_207_clk),
    .D(\reg_module/_00701_ ),
    .Q(\reg_module/gprf[701] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20286_  (.CLK(clknet_leaf_217_clk),
    .D(\reg_module/_00702_ ),
    .Q(\reg_module/gprf[702] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20287_  (.CLK(clknet_leaf_214_clk),
    .D(\reg_module/_00703_ ),
    .Q(\reg_module/gprf[703] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20288_  (.CLK(clknet_leaf_176_clk),
    .D(\reg_module/_00704_ ),
    .Q(\reg_module/gprf[704] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20289_  (.CLK(clknet_leaf_177_clk),
    .D(\reg_module/_00705_ ),
    .Q(\reg_module/gprf[705] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20290_  (.CLK(clknet_leaf_169_clk),
    .D(\reg_module/_00706_ ),
    .Q(\reg_module/gprf[706] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20291_  (.CLK(clknet_leaf_162_clk),
    .D(\reg_module/_00707_ ),
    .Q(\reg_module/gprf[707] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20292_  (.CLK(clknet_leaf_162_clk),
    .D(\reg_module/_00708_ ),
    .Q(\reg_module/gprf[708] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20293_  (.CLK(clknet_leaf_162_clk),
    .D(\reg_module/_00709_ ),
    .Q(\reg_module/gprf[709] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20294_  (.CLK(clknet_leaf_153_clk),
    .D(\reg_module/_00710_ ),
    .Q(\reg_module/gprf[710] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20295_  (.CLK(clknet_leaf_153_clk),
    .D(\reg_module/_00711_ ),
    .Q(\reg_module/gprf[711] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20296_  (.CLK(clknet_leaf_135_clk),
    .D(\reg_module/_00712_ ),
    .Q(\reg_module/gprf[712] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20297_  (.CLK(clknet_leaf_136_clk),
    .D(\reg_module/_00713_ ),
    .Q(\reg_module/gprf[713] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20298_  (.CLK(clknet_leaf_137_clk),
    .D(\reg_module/_00714_ ),
    .Q(\reg_module/gprf[714] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20299_  (.CLK(clknet_leaf_136_clk),
    .D(\reg_module/_00715_ ),
    .Q(\reg_module/gprf[715] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20300_  (.CLK(clknet_leaf_109_clk),
    .D(\reg_module/_00716_ ),
    .Q(\reg_module/gprf[716] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20301_  (.CLK(clknet_leaf_108_clk),
    .D(\reg_module/_00717_ ),
    .Q(\reg_module/gprf[717] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20302_  (.CLK(clknet_leaf_108_clk),
    .D(\reg_module/_00718_ ),
    .Q(\reg_module/gprf[718] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20303_  (.CLK(clknet_leaf_109_clk),
    .D(\reg_module/_00719_ ),
    .Q(\reg_module/gprf[719] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20304_  (.CLK(clknet_leaf_109_clk),
    .D(\reg_module/_00720_ ),
    .Q(\reg_module/gprf[720] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20305_  (.CLK(clknet_leaf_109_clk),
    .D(\reg_module/_00721_ ),
    .Q(\reg_module/gprf[721] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20306_  (.CLK(clknet_leaf_122_clk),
    .D(\reg_module/_00722_ ),
    .Q(\reg_module/gprf[722] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20307_  (.CLK(clknet_leaf_122_clk),
    .D(\reg_module/_00723_ ),
    .Q(\reg_module/gprf[723] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20308_  (.CLK(clknet_leaf_122_clk),
    .D(\reg_module/_00724_ ),
    .Q(\reg_module/gprf[724] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20309_  (.CLK(clknet_leaf_123_clk),
    .D(\reg_module/_00725_ ),
    .Q(\reg_module/gprf[725] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20310_  (.CLK(clknet_leaf_196_clk),
    .D(\reg_module/_00726_ ),
    .Q(\reg_module/gprf[726] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20311_  (.CLK(clknet_leaf_73_clk),
    .D(\reg_module/_00727_ ),
    .Q(\reg_module/gprf[727] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20312_  (.CLK(clknet_leaf_7_clk),
    .D(\reg_module/_00728_ ),
    .Q(\reg_module/gprf[728] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20313_  (.CLK(clknet_leaf_14_clk),
    .D(\reg_module/_00729_ ),
    .Q(\reg_module/gprf[729] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20314_  (.CLK(clknet_leaf_8_clk),
    .D(\reg_module/_00730_ ),
    .Q(\reg_module/gprf[730] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20315_  (.CLK(clknet_leaf_4_clk),
    .D(\reg_module/_00731_ ),
    .Q(\reg_module/gprf[731] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20316_  (.CLK(clknet_leaf_206_clk),
    .D(\reg_module/_00732_ ),
    .Q(\reg_module/gprf[732] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20317_  (.CLK(clknet_leaf_207_clk),
    .D(\reg_module/_00733_ ),
    .Q(\reg_module/gprf[733] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20318_  (.CLK(clknet_leaf_217_clk),
    .D(\reg_module/_00734_ ),
    .Q(\reg_module/gprf[734] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20319_  (.CLK(clknet_leaf_213_clk),
    .D(\reg_module/_00735_ ),
    .Q(\reg_module/gprf[735] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20320_  (.CLK(clknet_leaf_176_clk),
    .D(\reg_module/_00736_ ),
    .Q(\reg_module/gprf[736] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20321_  (.CLK(clknet_leaf_177_clk),
    .D(\reg_module/_00737_ ),
    .Q(\reg_module/gprf[737] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20322_  (.CLK(clknet_leaf_169_clk),
    .D(\reg_module/_00738_ ),
    .Q(\reg_module/gprf[738] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20323_  (.CLK(clknet_leaf_169_clk),
    .D(\reg_module/_00739_ ),
    .Q(\reg_module/gprf[739] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20324_  (.CLK(clknet_leaf_169_clk),
    .D(\reg_module/_00740_ ),
    .Q(\reg_module/gprf[740] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20325_  (.CLK(clknet_leaf_169_clk),
    .D(\reg_module/_00741_ ),
    .Q(\reg_module/gprf[741] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20326_  (.CLK(clknet_leaf_166_clk),
    .D(\reg_module/_00742_ ),
    .Q(\reg_module/gprf[742] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20327_  (.CLK(clknet_leaf_134_clk),
    .D(\reg_module/_00743_ ),
    .Q(\reg_module/gprf[743] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20328_  (.CLK(clknet_leaf_133_clk),
    .D(\reg_module/_00744_ ),
    .Q(\reg_module/gprf[744] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20329_  (.CLK(clknet_leaf_129_clk),
    .D(\reg_module/_00745_ ),
    .Q(\reg_module/gprf[745] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20330_  (.CLK(clknet_leaf_129_clk),
    .D(\reg_module/_00746_ ),
    .Q(\reg_module/gprf[746] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20331_  (.CLK(clknet_leaf_128_clk),
    .D(\reg_module/_00747_ ),
    .Q(\reg_module/gprf[747] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20332_  (.CLK(clknet_leaf_138_clk),
    .D(\reg_module/_00748_ ),
    .Q(\reg_module/gprf[748] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20333_  (.CLK(clknet_leaf_117_clk),
    .D(\reg_module/_00749_ ),
    .Q(\reg_module/gprf[749] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20334_  (.CLK(clknet_leaf_127_clk),
    .D(\reg_module/_00750_ ),
    .Q(\reg_module/gprf[750] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20335_  (.CLK(clknet_leaf_117_clk),
    .D(\reg_module/_00751_ ),
    .Q(\reg_module/gprf[751] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20336_  (.CLK(clknet_leaf_138_clk),
    .D(\reg_module/_00752_ ),
    .Q(\reg_module/gprf[752] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20337_  (.CLK(clknet_leaf_118_clk),
    .D(\reg_module/_00753_ ),
    .Q(\reg_module/gprf[753] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20338_  (.CLK(clknet_leaf_122_clk),
    .D(\reg_module/_00754_ ),
    .Q(\reg_module/gprf[754] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20339_  (.CLK(clknet_leaf_122_clk),
    .D(\reg_module/_00755_ ),
    .Q(\reg_module/gprf[755] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20340_  (.CLK(clknet_leaf_123_clk),
    .D(\reg_module/_00756_ ),
    .Q(\reg_module/gprf[756] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20341_  (.CLK(clknet_leaf_11_clk),
    .D(\reg_module/_00757_ ),
    .Q(\reg_module/gprf[757] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20342_  (.CLK(clknet_leaf_196_clk),
    .D(\reg_module/_00758_ ),
    .Q(\reg_module/gprf[758] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20343_  (.CLK(clknet_leaf_12_clk),
    .D(\reg_module/_00759_ ),
    .Q(\reg_module/gprf[759] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20344_  (.CLK(clknet_leaf_10_clk),
    .D(\reg_module/_00760_ ),
    .Q(\reg_module/gprf[760] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20345_  (.CLK(clknet_leaf_12_clk),
    .D(\reg_module/_00761_ ),
    .Q(\reg_module/gprf[761] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20346_  (.CLK(clknet_leaf_12_clk),
    .D(\reg_module/_00762_ ),
    .Q(\reg_module/gprf[762] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20347_  (.CLK(clknet_leaf_203_clk),
    .D(\reg_module/_00763_ ),
    .Q(\reg_module/gprf[763] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20348_  (.CLK(clknet_leaf_209_clk),
    .D(\reg_module/_00764_ ),
    .Q(\reg_module/gprf[764] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20349_  (.CLK(clknet_leaf_202_clk),
    .D(\reg_module/_00765_ ),
    .Q(\reg_module/gprf[765] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20350_  (.CLK(clknet_leaf_213_clk),
    .D(\reg_module/_00766_ ),
    .Q(\reg_module/gprf[766] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20351_  (.CLK(clknet_leaf_191_clk),
    .D(\reg_module/_00767_ ),
    .Q(\reg_module/gprf[767] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20352_  (.CLK(clknet_leaf_189_clk),
    .D(\reg_module/_00768_ ),
    .Q(\reg_module/gprf[768] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20353_  (.CLK(clknet_leaf_184_clk),
    .D(\reg_module/_00769_ ),
    .Q(\reg_module/gprf[769] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20354_  (.CLK(clknet_leaf_184_clk),
    .D(\reg_module/_00770_ ),
    .Q(\reg_module/gprf[770] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20355_  (.CLK(clknet_leaf_186_clk),
    .D(\reg_module/_00771_ ),
    .Q(\reg_module/gprf[771] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20356_  (.CLK(clknet_leaf_166_clk),
    .D(\reg_module/_00772_ ),
    .Q(\reg_module/gprf[772] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20357_  (.CLK(clknet_leaf_153_clk),
    .D(\reg_module/_00773_ ),
    .Q(\reg_module/gprf[773] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20358_  (.CLK(clknet_leaf_153_clk),
    .D(\reg_module/_00774_ ),
    .Q(\reg_module/gprf[774] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20359_  (.CLK(clknet_leaf_154_clk),
    .D(\reg_module/_00775_ ),
    .Q(\reg_module/gprf[775] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20360_  (.CLK(clknet_leaf_136_clk),
    .D(\reg_module/_00776_ ),
    .Q(\reg_module/gprf[776] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20361_  (.CLK(clknet_leaf_136_clk),
    .D(\reg_module/_00777_ ),
    .Q(\reg_module/gprf[777] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20362_  (.CLK(clknet_leaf_138_clk),
    .D(\reg_module/_00778_ ),
    .Q(\reg_module/gprf[778] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20363_  (.CLK(clknet_leaf_136_clk),
    .D(\reg_module/_00779_ ),
    .Q(\reg_module/gprf[779] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20364_  (.CLK(clknet_leaf_112_clk),
    .D(\reg_module/_00780_ ),
    .Q(\reg_module/gprf[780] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20365_  (.CLK(clknet_leaf_110_clk),
    .D(\reg_module/_00781_ ),
    .Q(\reg_module/gprf[781] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20366_  (.CLK(clknet_leaf_112_clk),
    .D(\reg_module/_00782_ ),
    .Q(\reg_module/gprf[782] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20367_  (.CLK(clknet_leaf_112_clk),
    .D(\reg_module/_00783_ ),
    .Q(\reg_module/gprf[783] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20368_  (.CLK(clknet_leaf_112_clk),
    .D(\reg_module/_00784_ ),
    .Q(\reg_module/gprf[784] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20369_  (.CLK(clknet_leaf_112_clk),
    .D(\reg_module/_00785_ ),
    .Q(\reg_module/gprf[785] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20370_  (.CLK(clknet_leaf_121_clk),
    .D(\reg_module/_00786_ ),
    .Q(\reg_module/gprf[786] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20371_  (.CLK(clknet_leaf_114_clk),
    .D(\reg_module/_00787_ ),
    .Q(\reg_module/gprf[787] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20372_  (.CLK(clknet_leaf_70_clk),
    .D(\reg_module/_00788_ ),
    .Q(\reg_module/gprf[788] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20373_  (.CLK(clknet_leaf_70_clk),
    .D(\reg_module/_00789_ ),
    .Q(\reg_module/gprf[789] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20374_  (.CLK(clknet_leaf_70_clk),
    .D(\reg_module/_00790_ ),
    .Q(\reg_module/gprf[790] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20375_  (.CLK(clknet_leaf_74_clk),
    .D(\reg_module/_00791_ ),
    .Q(\reg_module/gprf[791] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20376_  (.CLK(clknet_leaf_194_clk),
    .D(\reg_module/_00792_ ),
    .Q(\reg_module/gprf[792] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20377_  (.CLK(clknet_leaf_194_clk),
    .D(\reg_module/_00793_ ),
    .Q(\reg_module/gprf[793] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20378_  (.CLK(clknet_leaf_194_clk),
    .D(\reg_module/_00794_ ),
    .Q(\reg_module/gprf[794] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20379_  (.CLK(clknet_leaf_191_clk),
    .D(\reg_module/_00795_ ),
    .Q(\reg_module/gprf[795] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20380_  (.CLK(clknet_leaf_190_clk),
    .D(\reg_module/_00796_ ),
    .Q(\reg_module/gprf[796] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20381_  (.CLK(clknet_leaf_190_clk),
    .D(\reg_module/_00797_ ),
    .Q(\reg_module/gprf[797] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20382_  (.CLK(clknet_leaf_181_clk),
    .D(\reg_module/_00798_ ),
    .Q(\reg_module/gprf[798] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20383_  (.CLK(clknet_leaf_180_clk),
    .D(\reg_module/_00799_ ),
    .Q(\reg_module/gprf[799] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20384_  (.CLK(clknet_leaf_189_clk),
    .D(\reg_module/_00800_ ),
    .Q(\reg_module/gprf[800] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20385_  (.CLK(clknet_leaf_189_clk),
    .D(\reg_module/_00801_ ),
    .Q(\reg_module/gprf[801] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20386_  (.CLK(clknet_leaf_188_clk),
    .D(\reg_module/_00802_ ),
    .Q(\reg_module/gprf[802] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20387_  (.CLK(clknet_leaf_189_clk),
    .D(\reg_module/_00803_ ),
    .Q(\reg_module/gprf[803] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20388_  (.CLK(clknet_leaf_153_clk),
    .D(\reg_module/_00804_ ),
    .Q(\reg_module/gprf[804] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20389_  (.CLK(clknet_leaf_153_clk),
    .D(\reg_module/_00805_ ),
    .Q(\reg_module/gprf[805] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20390_  (.CLK(clknet_leaf_135_clk),
    .D(\reg_module/_00806_ ),
    .Q(\reg_module/gprf[806] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20391_  (.CLK(clknet_leaf_135_clk),
    .D(\reg_module/_00807_ ),
    .Q(\reg_module/gprf[807] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20392_  (.CLK(clknet_leaf_135_clk),
    .D(\reg_module/_00808_ ),
    .Q(\reg_module/gprf[808] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20393_  (.CLK(clknet_leaf_135_clk),
    .D(\reg_module/_00809_ ),
    .Q(\reg_module/gprf[809] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20394_  (.CLK(clknet_leaf_139_clk),
    .D(\reg_module/_00810_ ),
    .Q(\reg_module/gprf[810] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20395_  (.CLK(clknet_leaf_139_clk),
    .D(\reg_module/_00811_ ),
    .Q(\reg_module/gprf[811] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20396_  (.CLK(clknet_leaf_95_clk),
    .D(\reg_module/_00812_ ),
    .Q(\reg_module/gprf[812] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20397_  (.CLK(clknet_leaf_95_clk),
    .D(\reg_module/_00813_ ),
    .Q(\reg_module/gprf[813] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20398_  (.CLK(clknet_leaf_95_clk),
    .D(\reg_module/_00814_ ),
    .Q(\reg_module/gprf[814] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20399_  (.CLK(clknet_leaf_95_clk),
    .D(\reg_module/_00815_ ),
    .Q(\reg_module/gprf[815] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20400_  (.CLK(clknet_leaf_95_clk),
    .D(\reg_module/_00816_ ),
    .Q(\reg_module/gprf[816] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20401_  (.CLK(clknet_leaf_95_clk),
    .D(\reg_module/_00817_ ),
    .Q(\reg_module/gprf[817] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20402_  (.CLK(clknet_leaf_79_clk),
    .D(\reg_module/_00818_ ),
    .Q(\reg_module/gprf[818] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20403_  (.CLK(clknet_leaf_79_clk),
    .D(\reg_module/_00819_ ),
    .Q(\reg_module/gprf[819] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20404_  (.CLK(clknet_leaf_69_clk),
    .D(\reg_module/_00820_ ),
    .Q(\reg_module/gprf[820] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20405_  (.CLK(clknet_leaf_69_clk),
    .D(\reg_module/_00821_ ),
    .Q(\reg_module/gprf[821] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20406_  (.CLK(clknet_leaf_68_clk),
    .D(\reg_module/_00822_ ),
    .Q(\reg_module/gprf[822] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20407_  (.CLK(clknet_leaf_68_clk),
    .D(\reg_module/_00823_ ),
    .Q(\reg_module/gprf[823] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20408_  (.CLK(clknet_leaf_197_clk),
    .D(\reg_module/_00824_ ),
    .Q(\reg_module/gprf[824] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20409_  (.CLK(clknet_leaf_194_clk),
    .D(\reg_module/_00825_ ),
    .Q(\reg_module/gprf[825] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20410_  (.CLK(clknet_leaf_192_clk),
    .D(\reg_module/_00826_ ),
    .Q(\reg_module/gprf[826] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20411_  (.CLK(clknet_leaf_191_clk),
    .D(\reg_module/_00827_ ),
    .Q(\reg_module/gprf[827] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20412_  (.CLK(clknet_leaf_190_clk),
    .D(\reg_module/_00828_ ),
    .Q(\reg_module/gprf[828] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20413_  (.CLK(clknet_leaf_190_clk),
    .D(\reg_module/_00829_ ),
    .Q(\reg_module/gprf[829] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20414_  (.CLK(clknet_leaf_210_clk),
    .D(\reg_module/_00830_ ),
    .Q(\reg_module/gprf[830] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20415_  (.CLK(clknet_leaf_181_clk),
    .D(\reg_module/_00831_ ),
    .Q(\reg_module/gprf[831] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20416_  (.CLK(clknet_leaf_181_clk),
    .D(\reg_module/_00832_ ),
    .Q(\reg_module/gprf[832] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20417_  (.CLK(clknet_leaf_181_clk),
    .D(\reg_module/_00833_ ),
    .Q(\reg_module/gprf[833] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20418_  (.CLK(clknet_leaf_185_clk),
    .D(\reg_module/_00834_ ),
    .Q(\reg_module/gprf[834] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20419_  (.CLK(clknet_leaf_166_clk),
    .D(\reg_module/_00835_ ),
    .Q(\reg_module/gprf[835] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20420_  (.CLK(clknet_leaf_153_clk),
    .D(\reg_module/_00836_ ),
    .Q(\reg_module/gprf[836] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20421_  (.CLK(clknet_leaf_154_clk),
    .D(\reg_module/_00837_ ),
    .Q(\reg_module/gprf[837] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20422_  (.CLK(clknet_leaf_152_clk),
    .D(\reg_module/_00838_ ),
    .Q(\reg_module/gprf[838] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20423_  (.CLK(clknet_leaf_152_clk),
    .D(\reg_module/_00839_ ),
    .Q(\reg_module/gprf[839] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20424_  (.CLK(clknet_leaf_136_clk),
    .D(\reg_module/_00840_ ),
    .Q(\reg_module/gprf[840] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20425_  (.CLK(clknet_leaf_140_clk),
    .D(\reg_module/_00841_ ),
    .Q(\reg_module/gprf[841] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20426_  (.CLK(clknet_leaf_139_clk),
    .D(\reg_module/_00842_ ),
    .Q(\reg_module/gprf[842] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20427_  (.CLK(clknet_leaf_139_clk),
    .D(\reg_module/_00843_ ),
    .Q(\reg_module/gprf[843] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20428_  (.CLK(clknet_leaf_108_clk),
    .D(\reg_module/_00844_ ),
    .Q(\reg_module/gprf[844] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20429_  (.CLK(clknet_leaf_108_clk),
    .D(\reg_module/_00845_ ),
    .Q(\reg_module/gprf[845] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20430_  (.CLK(clknet_leaf_111_clk),
    .D(\reg_module/_00846_ ),
    .Q(\reg_module/gprf[846] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20431_  (.CLK(clknet_leaf_111_clk),
    .D(\reg_module/_00847_ ),
    .Q(\reg_module/gprf[847] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20432_  (.CLK(clknet_leaf_110_clk),
    .D(\reg_module/_00848_ ),
    .Q(\reg_module/gprf[848] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20433_  (.CLK(clknet_leaf_110_clk),
    .D(\reg_module/_00849_ ),
    .Q(\reg_module/gprf[849] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20434_  (.CLK(clknet_leaf_115_clk),
    .D(\reg_module/_00850_ ),
    .Q(\reg_module/gprf[850] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20435_  (.CLK(clknet_leaf_75_clk),
    .D(\reg_module/_00851_ ),
    .Q(\reg_module/gprf[851] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20436_  (.CLK(clknet_leaf_72_clk),
    .D(\reg_module/_00852_ ),
    .Q(\reg_module/gprf[852] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20437_  (.CLK(clknet_leaf_72_clk),
    .D(\reg_module/_00853_ ),
    .Q(\reg_module/gprf[853] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20438_  (.CLK(clknet_leaf_72_clk),
    .D(\reg_module/_00854_ ),
    .Q(\reg_module/gprf[854] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20439_  (.CLK(clknet_leaf_73_clk),
    .D(\reg_module/_00855_ ),
    .Q(\reg_module/gprf[855] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20440_  (.CLK(clknet_leaf_196_clk),
    .D(\reg_module/_00856_ ),
    .Q(\reg_module/gprf[856] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20441_  (.CLK(clknet_leaf_195_clk),
    .D(\reg_module/_00857_ ),
    .Q(\reg_module/gprf[857] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20442_  (.CLK(clknet_leaf_201_clk),
    .D(\reg_module/_00858_ ),
    .Q(\reg_module/gprf[858] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20443_  (.CLK(clknet_leaf_201_clk),
    .D(\reg_module/_00859_ ),
    .Q(\reg_module/gprf[859] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20444_  (.CLK(clknet_leaf_181_clk),
    .D(\reg_module/_00860_ ),
    .Q(\reg_module/gprf[860] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20445_  (.CLK(clknet_leaf_210_clk),
    .D(\reg_module/_00861_ ),
    .Q(\reg_module/gprf[861] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20446_  (.CLK(clknet_leaf_210_clk),
    .D(\reg_module/_00862_ ),
    .Q(\reg_module/gprf[862] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20447_  (.CLK(clknet_leaf_210_clk),
    .D(\reg_module/_00863_ ),
    .Q(\reg_module/gprf[863] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20448_  (.CLK(clknet_leaf_182_clk),
    .D(\reg_module/_00864_ ),
    .Q(\reg_module/gprf[864] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20449_  (.CLK(clknet_leaf_182_clk),
    .D(\reg_module/_00865_ ),
    .Q(\reg_module/gprf[865] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20450_  (.CLK(clknet_leaf_185_clk),
    .D(\reg_module/_00866_ ),
    .Q(\reg_module/gprf[866] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20451_  (.CLK(clknet_leaf_165_clk),
    .D(\reg_module/_00867_ ),
    .Q(\reg_module/gprf[867] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20452_  (.CLK(clknet_leaf_154_clk),
    .D(\reg_module/_00868_ ),
    .Q(\reg_module/gprf[868] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20453_  (.CLK(clknet_leaf_165_clk),
    .D(\reg_module/_00869_ ),
    .Q(\reg_module/gprf[869] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20454_  (.CLK(clknet_leaf_136_clk),
    .D(\reg_module/_00870_ ),
    .Q(\reg_module/gprf[870] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20455_  (.CLK(clknet_leaf_136_clk),
    .D(\reg_module/_00871_ ),
    .Q(\reg_module/gprf[871] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20456_  (.CLK(clknet_leaf_140_clk),
    .D(\reg_module/_00872_ ),
    .Q(\reg_module/gprf[872] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20457_  (.CLK(clknet_leaf_140_clk),
    .D(\reg_module/_00873_ ),
    .Q(\reg_module/gprf[873] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20458_  (.CLK(clknet_leaf_140_clk),
    .D(\reg_module/_00874_ ),
    .Q(\reg_module/gprf[874] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20459_  (.CLK(clknet_leaf_141_clk),
    .D(\reg_module/_00875_ ),
    .Q(\reg_module/gprf[875] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20460_  (.CLK(clknet_leaf_108_clk),
    .D(\reg_module/_00876_ ),
    .Q(\reg_module/gprf[876] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20461_  (.CLK(clknet_leaf_107_clk),
    .D(\reg_module/_00877_ ),
    .Q(\reg_module/gprf[877] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20462_  (.CLK(clknet_leaf_107_clk),
    .D(\reg_module/_00878_ ),
    .Q(\reg_module/gprf[878] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20463_  (.CLK(clknet_leaf_111_clk),
    .D(\reg_module/_00879_ ),
    .Q(\reg_module/gprf[879] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20464_  (.CLK(clknet_leaf_111_clk),
    .D(\reg_module/_00880_ ),
    .Q(\reg_module/gprf[880] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20465_  (.CLK(clknet_leaf_107_clk),
    .D(\reg_module/_00881_ ),
    .Q(\reg_module/gprf[881] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20466_  (.CLK(clknet_leaf_76_clk),
    .D(\reg_module/_00882_ ),
    .Q(\reg_module/gprf[882] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20467_  (.CLK(clknet_leaf_77_clk),
    .D(\reg_module/_00883_ ),
    .Q(\reg_module/gprf[883] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20468_  (.CLK(clknet_leaf_77_clk),
    .D(\reg_module/_00884_ ),
    .Q(\reg_module/gprf[884] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20469_  (.CLK(clknet_leaf_70_clk),
    .D(\reg_module/_00885_ ),
    .Q(\reg_module/gprf[885] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20470_  (.CLK(clknet_leaf_70_clk),
    .D(\reg_module/_00886_ ),
    .Q(\reg_module/gprf[886] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20471_  (.CLK(clknet_leaf_70_clk),
    .D(\reg_module/_00887_ ),
    .Q(\reg_module/gprf[887] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20472_  (.CLK(clknet_leaf_197_clk),
    .D(\reg_module/_00888_ ),
    .Q(\reg_module/gprf[888] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20473_  (.CLK(clknet_leaf_197_clk),
    .D(\reg_module/_00889_ ),
    .Q(\reg_module/gprf[889] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20474_  (.CLK(clknet_leaf_197_clk),
    .D(\reg_module/_00890_ ),
    .Q(\reg_module/gprf[890] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20475_  (.CLK(clknet_leaf_191_clk),
    .D(\reg_module/_00891_ ),
    .Q(\reg_module/gprf[891] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20476_  (.CLK(clknet_leaf_190_clk),
    .D(\reg_module/_00892_ ),
    .Q(\reg_module/gprf[892] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20477_  (.CLK(clknet_leaf_201_clk),
    .D(\reg_module/_00893_ ),
    .Q(\reg_module/gprf[893] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20478_  (.CLK(clknet_leaf_210_clk),
    .D(\reg_module/_00894_ ),
    .Q(\reg_module/gprf[894] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20479_  (.CLK(clknet_leaf_211_clk),
    .D(\reg_module/_00895_ ),
    .Q(\reg_module/gprf[895] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20480_  (.CLK(clknet_leaf_172_clk),
    .D(\reg_module/_00896_ ),
    .Q(\reg_module/gprf[896] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20481_  (.CLK(clknet_leaf_175_clk),
    .D(\reg_module/_00897_ ),
    .Q(\reg_module/gprf[897] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20482_  (.CLK(clknet_leaf_172_clk),
    .D(\reg_module/_00898_ ),
    .Q(\reg_module/gprf[898] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20483_  (.CLK(clknet_leaf_171_clk),
    .D(\reg_module/_00899_ ),
    .Q(\reg_module/gprf[899] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20484_  (.CLK(clknet_leaf_170_clk),
    .D(\reg_module/_00900_ ),
    .Q(\reg_module/gprf[900] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20485_  (.CLK(clknet_leaf_161_clk),
    .D(\reg_module/_00901_ ),
    .Q(\reg_module/gprf[901] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20486_  (.CLK(clknet_leaf_134_clk),
    .D(\reg_module/_00902_ ),
    .Q(\reg_module/gprf[902] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20487_  (.CLK(clknet_leaf_134_clk),
    .D(\reg_module/_00903_ ),
    .Q(\reg_module/gprf[903] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20488_  (.CLK(clknet_leaf_135_clk),
    .D(\reg_module/_00904_ ),
    .Q(\reg_module/gprf[904] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20489_  (.CLK(clknet_leaf_130_clk),
    .D(\reg_module/_00905_ ),
    .Q(\reg_module/gprf[905] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20490_  (.CLK(clknet_leaf_129_clk),
    .D(\reg_module/_00906_ ),
    .Q(\reg_module/gprf[906] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20491_  (.CLK(clknet_leaf_129_clk),
    .D(\reg_module/_00907_ ),
    .Q(\reg_module/gprf[907] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20492_  (.CLK(clknet_leaf_114_clk),
    .D(\reg_module/_00908_ ),
    .Q(\reg_module/gprf[908] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20493_  (.CLK(clknet_leaf_114_clk),
    .D(\reg_module/_00909_ ),
    .Q(\reg_module/gprf[909] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20494_  (.CLK(clknet_leaf_114_clk),
    .D(\reg_module/_00910_ ),
    .Q(\reg_module/gprf[910] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20495_  (.CLK(clknet_leaf_114_clk),
    .D(\reg_module/_00911_ ),
    .Q(\reg_module/gprf[911] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20496_  (.CLK(clknet_leaf_114_clk),
    .D(\reg_module/_00912_ ),
    .Q(\reg_module/gprf[912] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20497_  (.CLK(clknet_leaf_114_clk),
    .D(\reg_module/_00913_ ),
    .Q(\reg_module/gprf[913] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20498_  (.CLK(clknet_leaf_74_clk),
    .D(\reg_module/_00914_ ),
    .Q(\reg_module/gprf[914] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20499_  (.CLK(clknet_leaf_73_clk),
    .D(\reg_module/_00915_ ),
    .Q(\reg_module/gprf[915] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20500_  (.CLK(clknet_leaf_74_clk),
    .D(\reg_module/_00916_ ),
    .Q(\reg_module/gprf[916] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20501_  (.CLK(clknet_leaf_73_clk),
    .D(\reg_module/_00917_ ),
    .Q(\reg_module/gprf[917] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20502_  (.CLK(clknet_leaf_13_clk),
    .D(\reg_module/_00918_ ),
    .Q(\reg_module/gprf[918] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20503_  (.CLK(clknet_leaf_12_clk),
    .D(\reg_module/_00919_ ),
    .Q(\reg_module/gprf[919] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20504_  (.CLK(clknet_leaf_9_clk),
    .D(\reg_module/_00920_ ),
    .Q(\reg_module/gprf[920] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20505_  (.CLK(clknet_leaf_9_clk),
    .D(\reg_module/_00921_ ),
    .Q(\reg_module/gprf[921] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20506_  (.CLK(clknet_leaf_198_clk),
    .D(\reg_module/_00922_ ),
    .Q(\reg_module/gprf[922] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20507_  (.CLK(clknet_leaf_203_clk),
    .D(\reg_module/_00923_ ),
    .Q(\reg_module/gprf[923] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20508_  (.CLK(clknet_leaf_202_clk),
    .D(\reg_module/_00924_ ),
    .Q(\reg_module/gprf[924] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20509_  (.CLK(clknet_leaf_202_clk),
    .D(\reg_module/_00925_ ),
    .Q(\reg_module/gprf[925] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20510_  (.CLK(clknet_leaf_216_clk),
    .D(\reg_module/_00926_ ),
    .Q(\reg_module/gprf[926] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20511_  (.CLK(clknet_leaf_216_clk),
    .D(\reg_module/_00927_ ),
    .Q(\reg_module/gprf[927] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20512_  (.CLK(clknet_leaf_179_clk),
    .D(\reg_module/_00928_ ),
    .Q(\reg_module/gprf[928] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20513_  (.CLK(clknet_leaf_177_clk),
    .D(\reg_module/_00929_ ),
    .Q(\reg_module/gprf[929] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20514_  (.CLK(clknet_leaf_183_clk),
    .D(\reg_module/_00930_ ),
    .Q(\reg_module/gprf[930] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20515_  (.CLK(clknet_leaf_168_clk),
    .D(\reg_module/_00931_ ),
    .Q(\reg_module/gprf[931] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20516_  (.CLK(clknet_leaf_168_clk),
    .D(\reg_module/_00932_ ),
    .Q(\reg_module/gprf[932] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20517_  (.CLK(clknet_leaf_167_clk),
    .D(\reg_module/_00933_ ),
    .Q(\reg_module/gprf[933] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20518_  (.CLK(clknet_leaf_187_clk),
    .D(\reg_module/_00934_ ),
    .Q(\reg_module/gprf[934] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20519_  (.CLK(clknet_leaf_188_clk),
    .D(\reg_module/_00935_ ),
    .Q(\reg_module/gprf[935] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20520_  (.CLK(clknet_leaf_188_clk),
    .D(\reg_module/_00936_ ),
    .Q(\reg_module/gprf[936] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20521_  (.CLK(clknet_leaf_125_clk),
    .D(\reg_module/_00937_ ),
    .Q(\reg_module/gprf[937] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20522_  (.CLK(clknet_leaf_125_clk),
    .D(\reg_module/_00938_ ),
    .Q(\reg_module/gprf[938] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20523_  (.CLK(clknet_leaf_125_clk),
    .D(\reg_module/_00939_ ),
    .Q(\reg_module/gprf[939] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20524_  (.CLK(clknet_leaf_118_clk),
    .D(\reg_module/_00940_ ),
    .Q(\reg_module/gprf[940] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20525_  (.CLK(clknet_leaf_118_clk),
    .D(\reg_module/_00941_ ),
    .Q(\reg_module/gprf[941] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20526_  (.CLK(clknet_leaf_119_clk),
    .D(\reg_module/_00942_ ),
    .Q(\reg_module/gprf[942] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20527_  (.CLK(clknet_leaf_117_clk),
    .D(\reg_module/_00943_ ),
    .Q(\reg_module/gprf[943] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20528_  (.CLK(clknet_leaf_119_clk),
    .D(\reg_module/_00944_ ),
    .Q(\reg_module/gprf[944] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20529_  (.CLK(clknet_leaf_119_clk),
    .D(\reg_module/_00945_ ),
    .Q(\reg_module/gprf[945] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20530_  (.CLK(clknet_leaf_122_clk),
    .D(\reg_module/_00946_ ),
    .Q(\reg_module/gprf[946] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20531_  (.CLK(clknet_leaf_73_clk),
    .D(\reg_module/_00947_ ),
    .Q(\reg_module/gprf[947] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20532_  (.CLK(clknet_leaf_73_clk),
    .D(\reg_module/_00948_ ),
    .Q(\reg_module/gprf[948] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20533_  (.CLK(clknet_leaf_73_clk),
    .D(\reg_module/_00949_ ),
    .Q(\reg_module/gprf[949] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20534_  (.CLK(clknet_leaf_14_clk),
    .D(\reg_module/_00950_ ),
    .Q(\reg_module/gprf[950] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20535_  (.CLK(clknet_leaf_14_clk),
    .D(\reg_module/_00951_ ),
    .Q(\reg_module/gprf[951] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20536_  (.CLK(clknet_leaf_7_clk),
    .D(\reg_module/_00952_ ),
    .Q(\reg_module/gprf[952] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20537_  (.CLK(clknet_leaf_8_clk),
    .D(\reg_module/_00953_ ),
    .Q(\reg_module/gprf[953] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20538_  (.CLK(clknet_leaf_4_clk),
    .D(\reg_module/_00954_ ),
    .Q(\reg_module/gprf[954] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20539_  (.CLK(clknet_leaf_4_clk),
    .D(\reg_module/_00955_ ),
    .Q(\reg_module/gprf[955] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20540_  (.CLK(clknet_leaf_204_clk),
    .D(\reg_module/_00956_ ),
    .Q(\reg_module/gprf[956] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20541_  (.CLK(clknet_leaf_204_clk),
    .D(\reg_module/_00957_ ),
    .Q(\reg_module/gprf[957] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20542_  (.CLK(clknet_leaf_213_clk),
    .D(\reg_module/_00958_ ),
    .Q(\reg_module/gprf[958] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20543_  (.CLK(clknet_leaf_212_clk),
    .D(\reg_module/_00959_ ),
    .Q(\reg_module/gprf[959] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20544_  (.CLK(clknet_leaf_179_clk),
    .D(\reg_module/_00960_ ),
    .Q(\reg_module/gprf[960] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20545_  (.CLK(clknet_leaf_179_clk),
    .D(\reg_module/_00961_ ),
    .Q(\reg_module/gprf[961] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20546_  (.CLK(clknet_leaf_183_clk),
    .D(\reg_module/_00962_ ),
    .Q(\reg_module/gprf[962] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20547_  (.CLK(clknet_leaf_183_clk),
    .D(\reg_module/_00963_ ),
    .Q(\reg_module/gprf[963] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20548_  (.CLK(clknet_leaf_167_clk),
    .D(\reg_module/_00964_ ),
    .Q(\reg_module/gprf[964] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20549_  (.CLK(clknet_leaf_167_clk),
    .D(\reg_module/_00965_ ),
    .Q(\reg_module/gprf[965] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20550_  (.CLK(clknet_leaf_186_clk),
    .D(\reg_module/_00966_ ),
    .Q(\reg_module/gprf[966] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20551_  (.CLK(clknet_leaf_132_clk),
    .D(\reg_module/_00967_ ),
    .Q(\reg_module/gprf[967] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20552_  (.CLK(clknet_leaf_133_clk),
    .D(\reg_module/_00968_ ),
    .Q(\reg_module/gprf[968] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20553_  (.CLK(clknet_leaf_133_clk),
    .D(\reg_module/_00969_ ),
    .Q(\reg_module/gprf[969] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20554_  (.CLK(clknet_leaf_129_clk),
    .D(\reg_module/_00970_ ),
    .Q(\reg_module/gprf[970] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20555_  (.CLK(clknet_leaf_128_clk),
    .D(\reg_module/_00971_ ),
    .Q(\reg_module/gprf[971] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20556_  (.CLK(clknet_leaf_117_clk),
    .D(\reg_module/_00972_ ),
    .Q(\reg_module/gprf[972] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20557_  (.CLK(clknet_leaf_116_clk),
    .D(\reg_module/_00973_ ),
    .Q(\reg_module/gprf[973] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20558_  (.CLK(clknet_leaf_116_clk),
    .D(\reg_module/_00974_ ),
    .Q(\reg_module/gprf[974] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20559_  (.CLK(clknet_leaf_116_clk),
    .D(\reg_module/_00975_ ),
    .Q(\reg_module/gprf[975] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20560_  (.CLK(clknet_leaf_116_clk),
    .D(\reg_module/_00976_ ),
    .Q(\reg_module/gprf[976] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20561_  (.CLK(clknet_leaf_116_clk),
    .D(\reg_module/_00977_ ),
    .Q(\reg_module/gprf[977] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20562_  (.CLK(clknet_leaf_121_clk),
    .D(\reg_module/_00978_ ),
    .Q(\reg_module/gprf[978] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20563_  (.CLK(clknet_leaf_121_clk),
    .D(\reg_module/_00979_ ),
    .Q(\reg_module/gprf[979] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20564_  (.CLK(clknet_leaf_12_clk),
    .D(\reg_module/_00980_ ),
    .Q(\reg_module/gprf[980] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20565_  (.CLK(clknet_leaf_73_clk),
    .D(\reg_module/_00981_ ),
    .Q(\reg_module/gprf[981] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20566_  (.CLK(clknet_leaf_12_clk),
    .D(\reg_module/_00982_ ),
    .Q(\reg_module/gprf[982] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20567_  (.CLK(clknet_leaf_12_clk),
    .D(\reg_module/_00983_ ),
    .Q(\reg_module/gprf[983] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20568_  (.CLK(clknet_leaf_14_clk),
    .D(\reg_module/_00984_ ),
    .Q(\reg_module/gprf[984] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20569_  (.CLK(clknet_leaf_7_clk),
    .D(\reg_module/_00985_ ),
    .Q(\reg_module/gprf[985] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20570_  (.CLK(clknet_leaf_8_clk),
    .D(\reg_module/_00986_ ),
    .Q(\reg_module/gprf[986] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20571_  (.CLK(clknet_leaf_204_clk),
    .D(\reg_module/_00987_ ),
    .Q(\reg_module/gprf[987] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20572_  (.CLK(clknet_leaf_207_clk),
    .D(\reg_module/_00988_ ),
    .Q(\reg_module/gprf[988] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20573_  (.CLK(clknet_leaf_209_clk),
    .D(\reg_module/_00989_ ),
    .Q(\reg_module/gprf[989] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20574_  (.CLK(clknet_leaf_217_clk),
    .D(\reg_module/_00990_ ),
    .Q(\reg_module/gprf[990] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20575_  (.CLK(clknet_leaf_215_clk),
    .D(\reg_module/_00991_ ),
    .Q(\reg_module/gprf[991] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20576_  (.CLK(clknet_leaf_175_clk),
    .D(\reg_module/_00992_ ),
    .Q(\reg_module/gprf[992] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20577_  (.CLK(clknet_leaf_179_clk),
    .D(\reg_module/_00993_ ),
    .Q(\reg_module/gprf[993] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20578_  (.CLK(clknet_leaf_168_clk),
    .D(\reg_module/_00994_ ),
    .Q(\reg_module/gprf[994] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20579_  (.CLK(clknet_leaf_169_clk),
    .D(\reg_module/_00995_ ),
    .Q(\reg_module/gprf[995] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20580_  (.CLK(clknet_leaf_167_clk),
    .D(\reg_module/_00996_ ),
    .Q(\reg_module/gprf[996] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20581_  (.CLK(clknet_leaf_164_clk),
    .D(\reg_module/_00997_ ),
    .Q(\reg_module/gprf[997] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20582_  (.CLK(clknet_leaf_134_clk),
    .D(\reg_module/_00998_ ),
    .Q(\reg_module/gprf[998] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20583_  (.CLK(clknet_leaf_134_clk),
    .D(\reg_module/_00999_ ),
    .Q(\reg_module/gprf[999] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20584_  (.CLK(clknet_leaf_133_clk),
    .D(\reg_module/_01000_ ),
    .Q(\reg_module/gprf[1000] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20585_  (.CLK(clknet_leaf_130_clk),
    .D(\reg_module/_01001_ ),
    .Q(\reg_module/gprf[1001] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20586_  (.CLK(clknet_leaf_127_clk),
    .D(\reg_module/_01002_ ),
    .Q(\reg_module/gprf[1002] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20587_  (.CLK(clknet_leaf_128_clk),
    .D(\reg_module/_01003_ ),
    .Q(\reg_module/gprf[1003] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20588_  (.CLK(clknet_leaf_127_clk),
    .D(\reg_module/_01004_ ),
    .Q(\reg_module/gprf[1004] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20589_  (.CLK(clknet_leaf_110_clk),
    .D(\reg_module/_01005_ ),
    .Q(\reg_module/gprf[1005] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20590_  (.CLK(clknet_leaf_116_clk),
    .D(\reg_module/_01006_ ),
    .Q(\reg_module/gprf[1006] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20591_  (.CLK(clknet_leaf_110_clk),
    .D(\reg_module/_01007_ ),
    .Q(\reg_module/gprf[1007] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20592_  (.CLK(clknet_leaf_117_clk),
    .D(\reg_module/_01008_ ),
    .Q(\reg_module/gprf[1008] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20593_  (.CLK(clknet_leaf_113_clk),
    .D(\reg_module/_01009_ ),
    .Q(\reg_module/gprf[1009] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20594_  (.CLK(clknet_leaf_121_clk),
    .D(\reg_module/_01010_ ),
    .Q(\reg_module/gprf[1010] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20595_  (.CLK(clknet_leaf_122_clk),
    .D(\reg_module/_01011_ ),
    .Q(\reg_module/gprf[1011] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20596_  (.CLK(clknet_leaf_71_clk),
    .D(\reg_module/_01012_ ),
    .Q(\reg_module/gprf[1012] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20597_  (.CLK(clknet_leaf_73_clk),
    .D(\reg_module/_01013_ ),
    .Q(\reg_module/gprf[1013] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20598_  (.CLK(clknet_leaf_14_clk),
    .D(\reg_module/_01014_ ),
    .Q(\reg_module/gprf[1014] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20599_  (.CLK(clknet_leaf_12_clk),
    .D(\reg_module/_01015_ ),
    .Q(\reg_module/gprf[1015] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20600_  (.CLK(clknet_leaf_7_clk),
    .D(\reg_module/_01016_ ),
    .Q(\reg_module/gprf[1016] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20601_  (.CLK(clknet_leaf_8_clk),
    .D(\reg_module/_01017_ ),
    .Q(\reg_module/gprf[1017] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20602_  (.CLK(clknet_leaf_198_clk),
    .D(\reg_module/_01018_ ),
    .Q(\reg_module/gprf[1018] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20603_  (.CLK(clknet_leaf_202_clk),
    .D(\reg_module/_01019_ ),
    .Q(\reg_module/gprf[1019] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20604_  (.CLK(clknet_leaf_207_clk),
    .D(\reg_module/_01020_ ),
    .Q(\reg_module/gprf[1020] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20605_  (.CLK(clknet_leaf_210_clk),
    .D(\reg_module/_01021_ ),
    .Q(\reg_module/gprf[1021] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20606_  (.CLK(clknet_leaf_217_clk),
    .D(\reg_module/_01022_ ),
    .Q(\reg_module/gprf[1022] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20607_  (.CLK(clknet_leaf_216_clk),
    .D(\reg_module/_01023_ ),
    .Q(\reg_module/gprf[1023] ));
 sky130_fd_sc_hd__dfxtp_2 \reg_module/_20608_  (.CLK(clknet_leaf_20_clk),
    .D(\reg_module/_01024_ ),
    .Q(\reg_module/rRs1[0] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20609_  (.CLK(clknet_leaf_20_clk),
    .D(\reg_module/_01025_ ),
    .Q(\reg_module/rRs1[1] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20610_  (.CLK(clknet_leaf_20_clk),
    .D(\reg_module/_01026_ ),
    .Q(\reg_module/rRs1[2] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20611_  (.CLK(clknet_leaf_19_clk),
    .D(\reg_module/_01027_ ),
    .Q(\reg_module/rRs1[3] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20612_  (.CLK(clknet_leaf_63_clk),
    .D(\reg_module/_01028_ ),
    .Q(\reg_module/rRs1[4] ));
 sky130_fd_sc_hd__dfxtp_2 \reg_module/_20613_  (.CLK(clknet_leaf_20_clk),
    .D(\reg_module/_01029_ ),
    .Q(\reg_module/rRs2[0] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20614_  (.CLK(clknet_leaf_64_clk),
    .D(\reg_module/_01030_ ),
    .Q(\reg_module/rRs2[1] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20615_  (.CLK(clknet_leaf_19_clk),
    .D(\reg_module/_01031_ ),
    .Q(\reg_module/rRs2[2] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20616_  (.CLK(clknet_leaf_19_clk),
    .D(\reg_module/_01032_ ),
    .Q(\reg_module/rRs2[3] ));
 sky130_fd_sc_hd__dfxtp_1 \reg_module/_20617_  (.CLK(clknet_leaf_19_clk),
    .D(\reg_module/_01033_ ),
    .Q(\reg_module/rRs2[4] ));
 sky130_fd_sc_hd__nor2b_2 \rpc/_238_  (.A(net263),
    .B_N(net1073),
    .Y(\rpc/_032_ ));
 sky130_fd_sc_hd__clkbuf_2 \rpc/_239_  (.A(\rpc/_032_ ),
    .X(\rpc/_033_ ));
 sky130_fd_sc_hd__clkbuf_2 \rpc/_240_  (.A(\rpc/_032_ ),
    .X(\rpc/_034_ ));
 sky130_fd_sc_hd__o21ai_1 \rpc/_241_  (.A1(net378),
    .A2(net960),
    .B1(\rpc/_034_ ),
    .Y(\rpc/_035_ ));
 sky130_fd_sc_hd__a21o_1 \rpc/_242_  (.A1(net960),
    .A2(\wPcNextCond[2] ),
    .B1(\rpc/_035_ ),
    .X(\rpc/_036_ ));
 sky130_fd_sc_hd__o211a_1 \rpc/_243_  (.A1(net378),
    .A2(\rpc/_033_ ),
    .B1(net1027),
    .C1(\rpc/_036_ ),
    .X(\rpc/_000_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_244_  (.A(\rpc/_035_ ),
    .Y(\rpc/_037_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_245_  (.A(net377),
    .B(net379),
    .Y(\rpc/_038_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_246_  (.A(net959),
    .Y(\rpc/_039_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_247_  (.A(\rpc/_032_ ),
    .Y(\rpc/_040_ ));
 sky130_fd_sc_hd__clkbuf_2 \rpc/_248_  (.A(\rpc/_040_ ),
    .X(\rpc/_041_ ));
 sky130_fd_sc_hd__a21o_1 \rpc/_249_  (.A1(\rpc/_038_ ),
    .A2(\rpc/_039_ ),
    .B1(\rpc/_041_ ),
    .X(\rpc/_042_ ));
 sky130_fd_sc_hd__a21o_1 \rpc/_250_  (.A1(net960),
    .A2(\wPcNextCond[3] ),
    .B1(\rpc/_042_ ),
    .X(\rpc/_043_ ));
 sky130_fd_sc_hd__o211a_1 \rpc/_251_  (.A1(net1331),
    .A2(\rpc/_037_ ),
    .B1(net1027),
    .C1(\rpc/_043_ ),
    .X(\rpc/_001_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_252_  (.A(net376),
    .Y(\rpc/_044_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_253_  (.A(\rpc/_044_ ),
    .B(\rpc/_038_ ),
    .Y(\rpc/_045_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_254_  (.A(net959),
    .B(\rpc/_040_ ),
    .Y(\rpc/_046_ ));
 sky130_fd_sc_hd__clkbuf_2 \rpc/_255_  (.A(\rpc/_046_ ),
    .X(\rpc/_047_ ));
 sky130_fd_sc_hd__nand2_2 \rpc/_256_  (.A(\rpc/_032_ ),
    .B(net960),
    .Y(\rpc/_048_ ));
 sky130_fd_sc_hd__o21ai_1 \rpc/_257_  (.A1(\wPcNextCond[4] ),
    .A2(\rpc/_048_ ),
    .B1(net1027),
    .Y(\rpc/_049_ ));
 sky130_fd_sc_hd__a221oi_1 \rpc/_258_  (.A1(\rpc/_045_ ),
    .A2(\rpc/_047_ ),
    .B1(\rpc/_042_ ),
    .B2(\rpc/_044_ ),
    .C1(\rpc/_049_ ),
    .Y(\rpc/_002_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_259_  (.A(\rpc/_048_ ),
    .Y(\rpc/_050_ ));
 sky130_fd_sc_hd__clkbuf_2 \rpc/_260_  (.A(\rpc/_050_ ),
    .X(\rpc/_051_ ));
 sky130_fd_sc_hd__a22o_1 \rpc/_261_  (.A1(net375),
    .A2(\rpc/_041_ ),
    .B1(\rpc/_051_ ),
    .B2(\wPcNextCond[5] ),
    .X(\rpc/_052_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_262_  (.A(net375),
    .B(net161),
    .Y(\rpc/_053_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_263_  (.A(\rpc/_038_ ),
    .B(\rpc/_053_ ),
    .Y(\rpc/_054_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_264_  (.A(\rpc/_046_ ),
    .Y(\rpc/_055_ ));
 sky130_fd_sc_hd__buf_6 \rpc/_265_  (.A(\rpc/_055_ ),
    .X(\rpc/_056_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_266_  (.A(\rpc/_054_ ),
    .B(\rpc/_056_ ),
    .Y(\rpc/_057_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_267_  (.A1(net375),
    .A2(\rpc/_045_ ),
    .B1(\rpc/_057_ ),
    .X(\rpc/_058_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_268_  (.A1(\rpc/_052_ ),
    .A2(\rpc/_058_ ),
    .B1(net1027),
    .X(\rpc/_003_ ));
 sky130_fd_sc_hd__clkbuf_2 \rpc/_269_  (.A(\rpc/_048_ ),
    .X(\rpc/_059_ ));
 sky130_fd_sc_hd__buf_2 \rpc/_270_  (.A(\rpc/_059_ ),
    .X(\rpc/_060_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_271_  (.A(\rpc/_054_ ),
    .B(\rpc/_034_ ),
    .Y(\rpc/_061_ ));
 sky130_fd_sc_hd__xor2_1 \rpc/_272_  (.A(net373),
    .B(\rpc/_061_ ),
    .X(\rpc/_062_ ));
 sky130_fd_sc_hd__clkbuf_2 \rpc/_273_  (.A(\rpc/_048_ ),
    .X(\rpc/_063_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_274_  (.A(\rpc/_062_ ),
    .B(\rpc/_063_ ),
    .Y(\rpc/_064_ ));
 sky130_fd_sc_hd__o211a_1 \rpc/_275_  (.A1(\wPcNextCond[6] ),
    .A2(\rpc/_060_ ),
    .B1(net1029),
    .C1(\rpc/_064_ ),
    .X(\rpc/_004_ ));
 sky130_fd_sc_hd__and2_1 \rpc/_276_  (.A(\rpc/_054_ ),
    .B(net373),
    .X(\rpc/_065_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_277_  (.A(\rpc/_065_ ),
    .B(\rpc/_034_ ),
    .Y(\rpc/_066_ ));
 sky130_fd_sc_hd__xor2_1 \rpc/_278_  (.A(net372),
    .B(\rpc/_066_ ),
    .X(\rpc/_067_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_279_  (.A(\rpc/_067_ ),
    .B(\rpc/_063_ ),
    .Y(\rpc/_068_ ));
 sky130_fd_sc_hd__o211a_1 \rpc/_280_  (.A1(\wPcNextCond[7] ),
    .A2(\rpc/_060_ ),
    .B1(net1029),
    .C1(\rpc/_068_ ),
    .X(\rpc/_005_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_281_  (.A(net165),
    .Y(\rpc/_069_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_282_  (.A(\rpc/_065_ ),
    .B(net372),
    .Y(\rpc/_070_ ));
 sky130_fd_sc_hd__or2_1 \rpc/_283_  (.A(\rpc/_069_ ),
    .B(\rpc/_070_ ),
    .X(\rpc/_071_ ));
 sky130_fd_sc_hd__a21o_1 \rpc/_284_  (.A1(\rpc/_071_ ),
    .A2(\rpc/_039_ ),
    .B1(\rpc/_041_ ),
    .X(\rpc/_072_ ));
 sky130_fd_sc_hd__clkbuf_2 \rpc/_285_  (.A(\rpc/_040_ ),
    .X(\rpc/_073_ ));
 sky130_fd_sc_hd__o21ai_1 \rpc/_286_  (.A1(\rpc/_073_ ),
    .A2(\rpc/_070_ ),
    .B1(\rpc/_069_ ),
    .Y(\rpc/_074_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_287_  (.A(\rpc/_072_ ),
    .B(\rpc/_074_ ),
    .Y(\rpc/_075_ ));
 sky130_fd_sc_hd__clkbuf_2 \rpc/_288_  (.A(\rpc/_050_ ),
    .X(\rpc/_076_ ));
 sky130_fd_sc_hd__clkbuf_2 \rpc/_289_  (.A(\rpc/_076_ ),
    .X(\rpc/_077_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_290_  (.A(\rpc/_077_ ),
    .B(\wPcNextCond[8] ),
    .Y(\rpc/_078_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_291_  (.A(net1028),
    .Y(\rpc/_079_ ));
 sky130_fd_sc_hd__clkbuf_2 \rpc/_292_  (.A(\rpc/_079_ ),
    .X(\rpc/_080_ ));
 sky130_fd_sc_hd__a21oi_1 \rpc/_293_  (.A1(\rpc/_075_ ),
    .A2(\rpc/_078_ ),
    .B1(\rpc/_080_ ),
    .Y(\rpc/_006_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_294_  (.A(\rpc/_072_ ),
    .B(net370),
    .Y(\rpc/_081_ ));
 sky130_fd_sc_hd__or3_1 \rpc/_295_  (.A(net166),
    .B(net959),
    .C(\rpc/_040_ ),
    .X(\rpc/_082_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_296_  (.A(\rpc/_076_ ),
    .B(\wPcNextCond[9] ),
    .Y(\rpc/_083_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_297_  (.A1(\rpc/_082_ ),
    .A2(\rpc/_071_ ),
    .B1(\rpc/_083_ ),
    .X(\rpc/_084_ ));
 sky130_fd_sc_hd__a21oi_1 \rpc/_298_  (.A1(\rpc/_081_ ),
    .A2(\rpc/_084_ ),
    .B1(\rpc/_080_ ),
    .Y(\rpc/_007_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_299_  (.A(net164),
    .B(net374),
    .Y(\rpc/_085_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_300_  (.A(net166),
    .B(net165),
    .Y(\rpc/_086_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_301_  (.A(\rpc/_085_ ),
    .B(\rpc/_086_ ),
    .Y(\rpc/_087_ ));
 sky130_fd_sc_hd__nand2_2 \rpc/_302_  (.A(\rpc/_054_ ),
    .B(\rpc/_087_ ),
    .Y(\rpc/_088_ ));
 sky130_fd_sc_hd__or3_1 \rpc/_303_  (.A(net369),
    .B(\rpc/_040_ ),
    .C(\rpc/_088_ ),
    .X(\rpc/_089_ ));
 sky130_fd_sc_hd__o21ai_1 \rpc/_304_  (.A1(\rpc/_073_ ),
    .A2(\rpc/_088_ ),
    .B1(net369),
    .Y(\rpc/_090_ ));
 sky130_fd_sc_hd__o21ai_1 \rpc/_305_  (.A1(\wPcNextCond[10] ),
    .A2(\rpc/_059_ ),
    .B1(net1027),
    .Y(\rpc/_091_ ));
 sky130_fd_sc_hd__a31o_1 \rpc/_306_  (.A1(\rpc/_089_ ),
    .A2(\rpc/_063_ ),
    .A3(\rpc/_090_ ),
    .B1(\rpc/_091_ ),
    .X(\rpc/_092_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_307_  (.A(\rpc/_092_ ),
    .Y(\rpc/_008_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_308_  (.A(net369),
    .Y(\rpc/_093_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_309_  (.A(\rpc/_093_ ),
    .B(\rpc/_088_ ),
    .Y(\rpc/_094_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_310_  (.A(\rpc/_094_ ),
    .B(\rpc/_034_ ),
    .Y(\rpc/_095_ ));
 sky130_fd_sc_hd__o21ai_1 \rpc/_311_  (.A1(net366),
    .A2(\rpc/_095_ ),
    .B1(\rpc/_059_ ),
    .Y(\rpc/_096_ ));
 sky130_fd_sc_hd__a21o_1 \rpc/_312_  (.A1(net366),
    .A2(\rpc/_095_ ),
    .B1(\rpc/_096_ ),
    .X(\rpc/_097_ ));
 sky130_fd_sc_hd__o211ai_1 \rpc/_313_  (.A1(\wPcNextCond[11] ),
    .A2(\rpc/_060_ ),
    .B1(net1028),
    .C1(\rpc/_097_ ),
    .Y(\rpc/_098_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_314_  (.A(\rpc/_098_ ),
    .Y(\rpc/_009_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_315_  (.A(\rpc/_094_ ),
    .B(net366),
    .Y(\rpc/_099_ ));
 sky130_fd_sc_hd__nor3_1 \rpc/_316_  (.A(net364),
    .B(\rpc/_073_ ),
    .C(\rpc/_099_ ),
    .Y(\rpc/_100_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_317_  (.A1(\rpc/_041_ ),
    .A2(\rpc/_099_ ),
    .B1(net364),
    .X(\rpc/_101_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_318_  (.A1(\wPcNextCond[12] ),
    .A2(\rpc/_059_ ),
    .B1(net1028),
    .X(\rpc/_102_ ));
 sky130_fd_sc_hd__o31ai_1 \rpc/_319_  (.A1(\rpc/_077_ ),
    .A2(\rpc/_100_ ),
    .A3(\rpc/_101_ ),
    .B1(\rpc/_102_ ),
    .Y(\rpc/_103_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_320_  (.A(\rpc/_103_ ),
    .Y(\rpc/_010_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_321_  (.A(net366),
    .B(net368),
    .Y(\rpc/_104_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_322_  (.A(net362),
    .B(net363),
    .Y(\rpc/_105_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_323_  (.A(\rpc/_104_ ),
    .B(\rpc/_105_ ),
    .Y(\rpc/_106_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_324_  (.A(\rpc/_106_ ),
    .Y(\rpc/_107_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_325_  (.A(\rpc/_107_ ),
    .B(\rpc/_088_ ),
    .Y(\rpc/_108_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_326_  (.A(\rpc/_108_ ),
    .Y(\rpc/_109_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_327_  (.A(\rpc/_109_ ),
    .B(\rpc/_047_ ),
    .Y(\rpc/_110_ ));
 sky130_fd_sc_hd__clkbuf_2 \rpc/_328_  (.A(\rpc/_032_ ),
    .X(\rpc/_111_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_329_  (.A(\rpc/_110_ ),
    .B(\rpc/_111_ ),
    .Y(\rpc/_112_ ));
 sky130_fd_sc_hd__and2_1 \rpc/_330_  (.A(\rpc/_112_ ),
    .B(net362),
    .X(\rpc/_113_ ));
 sky130_fd_sc_hd__or2b_1 \rpc/_331_  (.A(\rpc/_099_ ),
    .B_N(net363),
    .X(\rpc/_114_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_332_  (.A(\rpc/_051_ ),
    .B(\wPcNextCond[13] ),
    .Y(\rpc/_115_ ));
 sky130_fd_sc_hd__o21ai_1 \rpc/_333_  (.A1(\rpc/_110_ ),
    .A2(\rpc/_114_ ),
    .B1(\rpc/_115_ ),
    .Y(\rpc/_116_ ));
 sky130_fd_sc_hd__o21ai_1 \rpc/_334_  (.A1(\rpc/_113_ ),
    .A2(\rpc/_116_ ),
    .B1(net1020),
    .Y(\rpc/_117_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_335_  (.A(\rpc/_117_ ),
    .Y(\rpc/_011_ ));
 sky130_fd_sc_hd__and2_1 \rpc/_336_  (.A(\rpc/_112_ ),
    .B(net360),
    .X(\rpc/_118_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_337_  (.A(net360),
    .Y(\rpc/_119_ ));
 sky130_fd_sc_hd__a32o_1 \rpc/_338_  (.A1(\rpc/_108_ ),
    .A2(\rpc/_119_ ),
    .A3(\rpc/_047_ ),
    .B1(\wPcNextCond[14] ),
    .B2(\rpc/_051_ ),
    .X(\rpc/_120_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_339_  (.A1(\rpc/_118_ ),
    .A2(\rpc/_120_ ),
    .B1(net1020),
    .X(\rpc/_012_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_340_  (.A(\rpc/_119_ ),
    .B(\rpc/_109_ ),
    .Y(\rpc/_121_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_341_  (.A(\rpc/_121_ ),
    .B(\rpc/_111_ ),
    .Y(\rpc/_122_ ));
 sky130_fd_sc_hd__xor2_1 \rpc/_342_  (.A(net357),
    .B(\rpc/_122_ ),
    .X(\rpc/_123_ ));
 sky130_fd_sc_hd__o21ai_1 \rpc/_343_  (.A1(\wPcNextCond[15] ),
    .A2(\rpc/_063_ ),
    .B1(net1020),
    .Y(\rpc/_124_ ));
 sky130_fd_sc_hd__a21oi_1 \rpc/_344_  (.A1(\rpc/_123_ ),
    .A2(\rpc/_060_ ),
    .B1(\rpc/_124_ ),
    .Y(\rpc/_013_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_345_  (.A(net357),
    .B(net360),
    .Y(\rpc/_125_ ));
 sky130_fd_sc_hd__o21ai_1 \rpc/_346_  (.A1(\rpc/_125_ ),
    .A2(\rpc/_109_ ),
    .B1(net354),
    .Y(\rpc/_126_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_347_  (.A(\rpc/_125_ ),
    .Y(\rpc/_127_ ));
 sky130_fd_sc_hd__nand3b_1 \rpc/_348_  (.A_N(net354),
    .B(\rpc/_108_ ),
    .C(\rpc/_127_ ),
    .Y(\rpc/_128_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_349_  (.A(\rpc/_126_ ),
    .B(\rpc/_128_ ),
    .Y(\rpc/_129_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_350_  (.A1(\rpc/_039_ ),
    .A2(\wPcNextCond[16] ),
    .B1(\rpc/_033_ ),
    .X(\rpc/_130_ ));
 sky130_fd_sc_hd__o21ai_1 \rpc/_351_  (.A1(net959),
    .A2(\rpc/_129_ ),
    .B1(\rpc/_130_ ),
    .Y(\rpc/_131_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_352_  (.A(\rpc/_073_ ),
    .B(net354),
    .Y(\rpc/_132_ ));
 sky130_fd_sc_hd__a21oi_1 \rpc/_353_  (.A1(\rpc/_131_ ),
    .A2(\rpc/_132_ ),
    .B1(\rpc/_080_ ),
    .Y(\rpc/_014_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_354_  (.A(net352),
    .B(net354),
    .Y(\rpc/_133_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_355_  (.A(\rpc/_125_ ),
    .B(\rpc/_133_ ),
    .Y(\rpc/_134_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_356_  (.A(\rpc/_106_ ),
    .B(\rpc/_134_ ),
    .Y(\rpc/_135_ ));
 sky130_fd_sc_hd__nor2_2 \rpc/_357_  (.A(\rpc/_088_ ),
    .B(\rpc/_135_ ),
    .Y(\rpc/_136_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_358_  (.A(\rpc/_055_ ),
    .B(\rpc/_136_ ),
    .Y(\rpc/_137_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_359_  (.A(\rpc/_137_ ),
    .B(net355),
    .Y(\rpc/_138_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_360_  (.A(\rpc/_121_ ),
    .B(net357),
    .Y(\rpc/_139_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_361_  (.A(\rpc/_076_ ),
    .B(\wPcNextCond[17] ),
    .Y(\rpc/_140_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_362_  (.A1(\rpc/_138_ ),
    .A2(\rpc/_139_ ),
    .B1(\rpc/_140_ ),
    .X(\rpc/_141_ ));
 sky130_fd_sc_hd__or2_1 \rpc/_363_  (.A(\rpc/_040_ ),
    .B(\rpc/_137_ ),
    .X(\rpc/_142_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_364_  (.A(\rpc/_142_ ),
    .B(net353),
    .Y(\rpc/_143_ ));
 sky130_fd_sc_hd__a21o_1 \rpc/_365_  (.A1(\rpc/_141_ ),
    .A2(\rpc/_143_ ),
    .B1(\rpc/_079_ ),
    .X(\rpc/_144_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_366_  (.A(\rpc/_144_ ),
    .Y(\rpc/_015_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_367_  (.A(net350),
    .B(\rpc/_056_ ),
    .Y(\rpc/_145_ ));
 sky130_fd_sc_hd__buf_6 \rpc/_368_  (.A(\rpc/_136_ ),
    .X(\rpc/_146_ ));
 sky130_fd_sc_hd__a22o_1 \rpc/_369_  (.A1(\wPcNextCond[18] ),
    .A2(\rpc/_076_ ),
    .B1(\rpc/_145_ ),
    .B2(\rpc/_146_ ),
    .X(\rpc/_147_ ));
 sky130_fd_sc_hd__and2_1 \rpc/_370_  (.A(\rpc/_142_ ),
    .B(net351),
    .X(\rpc/_148_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_371_  (.A1(\rpc/_147_ ),
    .A2(\rpc/_148_ ),
    .B1(net1028),
    .X(\rpc/_016_ ));
 sky130_fd_sc_hd__nand3_1 \rpc/_372_  (.A(\rpc/_146_ ),
    .B(net351),
    .C(\rpc/_034_ ),
    .Y(\rpc/_149_ ));
 sky130_fd_sc_hd__xor2_1 \rpc/_373_  (.A(net348),
    .B(\rpc/_149_ ),
    .X(\rpc/_150_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_374_  (.A(\rpc/_150_ ),
    .B(\rpc/_063_ ),
    .Y(\rpc/_151_ ));
 sky130_fd_sc_hd__o211a_1 \rpc/_375_  (.A1(\wPcNextCond[19] ),
    .A2(\rpc/_060_ ),
    .B1(net1020),
    .C1(\rpc/_151_ ),
    .X(\rpc/_017_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_376_  (.A(net348),
    .B(net350),
    .Y(\rpc/_152_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_377_  (.A(\rpc/_152_ ),
    .Y(\rpc/_153_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_378_  (.A(\rpc/_136_ ),
    .B(\rpc/_153_ ),
    .Y(\rpc/_154_ ));
 sky130_fd_sc_hd__or2_1 \rpc/_379_  (.A(net346),
    .B(\rpc/_154_ ),
    .X(\rpc/_155_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_380_  (.A(\rpc/_154_ ),
    .B(net346),
    .Y(\rpc/_156_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_381_  (.A(\rpc/_155_ ),
    .B(\rpc/_156_ ),
    .Y(\rpc/_157_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_382_  (.A1(\rpc/_039_ ),
    .A2(\wPcNextCond[20] ),
    .B1(\rpc/_033_ ),
    .X(\rpc/_158_ ));
 sky130_fd_sc_hd__o21ai_1 \rpc/_383_  (.A1(net959),
    .A2(\rpc/_157_ ),
    .B1(\rpc/_158_ ),
    .Y(\rpc/_159_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_384_  (.A(\rpc/_073_ ),
    .B(net346),
    .Y(\rpc/_160_ ));
 sky130_fd_sc_hd__a21oi_1 \rpc/_385_  (.A1(\rpc/_159_ ),
    .A2(\rpc/_160_ ),
    .B1(\rpc/_080_ ),
    .Y(\rpc/_018_ ));
 sky130_fd_sc_hd__nand3_1 \rpc/_386_  (.A(\rpc/_153_ ),
    .B(net345),
    .C(net346),
    .Y(\rpc/_161_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_387_  (.A(\rpc/_161_ ),
    .Y(\rpc/_162_ ));
 sky130_fd_sc_hd__a21o_1 \rpc/_388_  (.A1(\rpc/_146_ ),
    .A2(\rpc/_162_ ),
    .B1(\rpc/_056_ ),
    .X(\rpc/_163_ ));
 sky130_fd_sc_hd__nand2b_1 \rpc/_389_  (.A_N(\rpc/_154_ ),
    .B(net347),
    .Y(\rpc/_164_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_390_  (.A(\rpc/_076_ ),
    .B(\wPcNextCond[21] ),
    .Y(\rpc/_165_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_391_  (.A1(\rpc/_163_ ),
    .A2(\rpc/_164_ ),
    .B1(\rpc/_165_ ),
    .X(\rpc/_166_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_392_  (.A(\rpc/_163_ ),
    .B(\rpc/_111_ ),
    .Y(\rpc/_167_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_393_  (.A(\rpc/_167_ ),
    .B(net345),
    .Y(\rpc/_168_ ));
 sky130_fd_sc_hd__a21oi_1 \rpc/_394_  (.A1(\rpc/_166_ ),
    .A2(\rpc/_168_ ),
    .B1(\rpc/_080_ ),
    .Y(\rpc/_019_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_395_  (.A(net343),
    .B(\rpc/_056_ ),
    .Y(\rpc/_169_ ));
 sky130_fd_sc_hd__and3_1 \rpc/_396_  (.A(\rpc/_034_ ),
    .B(net959),
    .C(\wPcNextCond[22] ),
    .X(\rpc/_170_ ));
 sky130_fd_sc_hd__a31o_1 \rpc/_397_  (.A1(\rpc/_169_ ),
    .A2(\rpc/_146_ ),
    .A3(\rpc/_162_ ),
    .B1(\rpc/_170_ ),
    .X(\rpc/_171_ ));
 sky130_fd_sc_hd__and2_1 \rpc/_398_  (.A(\rpc/_167_ ),
    .B(net343),
    .X(\rpc/_172_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_399_  (.A1(\rpc/_171_ ),
    .A2(\rpc/_172_ ),
    .B1(net1020),
    .X(\rpc/_020_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_400_  (.A(net342),
    .Y(\rpc/_173_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_401_  (.A(\rpc/_173_ ),
    .B(\rpc/_033_ ),
    .Y(\rpc/_174_ ));
 sky130_fd_sc_hd__nand3_1 \rpc/_402_  (.A(\rpc/_146_ ),
    .B(net343),
    .C(\rpc/_162_ ),
    .Y(\rpc/_175_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_403_  (.A(\rpc/_175_ ),
    .B(\rpc/_173_ ),
    .Y(\rpc/_176_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_404_  (.A(\rpc/_173_ ),
    .B(\rpc/_175_ ),
    .Y(\rpc/_177_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_405_  (.A(\rpc/_177_ ),
    .B(\rpc/_033_ ),
    .Y(\rpc/_178_ ));
 sky130_fd_sc_hd__o211ai_1 \rpc/_406_  (.A1(\rpc/_047_ ),
    .A2(\rpc/_174_ ),
    .B1(\rpc/_176_ ),
    .C1(\rpc/_178_ ),
    .Y(\rpc/_179_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_407_  (.A(\rpc/_077_ ),
    .B(\wPcNextCond[23] ),
    .Y(\rpc/_180_ ));
 sky130_fd_sc_hd__a21oi_1 \rpc/_408_  (.A1(\rpc/_179_ ),
    .A2(\rpc/_180_ ),
    .B1(\rpc/_080_ ),
    .Y(\rpc/_021_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_409_  (.A(net340),
    .B(\rpc/_178_ ),
    .Y(\rpc/_181_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_410_  (.A(\rpc/_178_ ),
    .B(net340),
    .Y(\rpc/_182_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_411_  (.A(\rpc/_182_ ),
    .B(\rpc/_063_ ),
    .Y(\rpc/_183_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_412_  (.A1(\wPcNextCond[24] ),
    .A2(\rpc/_059_ ),
    .B1(net1020),
    .X(\rpc/_184_ ));
 sky130_fd_sc_hd__o21ai_1 \rpc/_413_  (.A1(\rpc/_181_ ),
    .A2(\rpc/_183_ ),
    .B1(\rpc/_184_ ),
    .Y(\rpc/_185_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_414_  (.A(\rpc/_185_ ),
    .Y(\rpc/_022_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_415_  (.A(net342),
    .B(net343),
    .Y(\rpc/_186_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_416_  (.A(\rpc/_186_ ),
    .Y(\rpc/_187_ ));
 sky130_fd_sc_hd__nand3_1 \rpc/_417_  (.A(\rpc/_187_ ),
    .B(net339),
    .C(net340),
    .Y(\rpc/_188_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_418_  (.A(\rpc/_188_ ),
    .B(\rpc/_161_ ),
    .Y(\rpc/_189_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_419_  (.A(\rpc/_136_ ),
    .B(\rpc/_189_ ),
    .Y(\rpc/_190_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_420_  (.A(\rpc/_190_ ),
    .B(\rpc/_047_ ),
    .Y(\rpc/_191_ ));
 sky130_fd_sc_hd__nand3b_1 \rpc/_421_  (.A_N(\rpc/_191_ ),
    .B(\rpc/_177_ ),
    .C(net340),
    .Y(\rpc/_192_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_422_  (.A(\rpc/_191_ ),
    .B(\rpc/_111_ ),
    .Y(\rpc/_193_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_423_  (.A(\rpc/_193_ ),
    .B(net339),
    .Y(\rpc/_194_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_424_  (.A(\rpc/_077_ ),
    .B(\wPcNextCond[25] ),
    .Y(\rpc/_195_ ));
 sky130_fd_sc_hd__nand3_1 \rpc/_425_  (.A(\rpc/_192_ ),
    .B(\rpc/_194_ ),
    .C(\rpc/_195_ ),
    .Y(\rpc/_196_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_426_  (.A(\rpc/_196_ ),
    .B(net1021),
    .Y(\rpc/_197_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_427_  (.A(\rpc/_197_ ),
    .Y(\rpc/_023_ ));
 sky130_fd_sc_hd__and2_1 \rpc/_428_  (.A(\rpc/_193_ ),
    .B(net336),
    .X(\rpc/_198_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_429_  (.A(\rpc/_190_ ),
    .Y(\rpc/_199_ ));
 sky130_fd_sc_hd__nor2_1 \rpc/_430_  (.A(net336),
    .B(\rpc/_056_ ),
    .Y(\rpc/_200_ ));
 sky130_fd_sc_hd__a22o_1 \rpc/_431_  (.A1(\wPcNextCond[26] ),
    .A2(\rpc/_051_ ),
    .B1(\rpc/_199_ ),
    .B2(\rpc/_200_ ),
    .X(\rpc/_201_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_432_  (.A1(\rpc/_198_ ),
    .A2(\rpc/_201_ ),
    .B1(net1021),
    .X(\rpc/_024_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_433_  (.A(net335),
    .B(net337),
    .Y(\rpc/_202_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_434_  (.A(\rpc/_202_ ),
    .Y(\rpc/_203_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_435_  (.A(\rpc/_199_ ),
    .B(\rpc/_203_ ),
    .Y(\rpc/_204_ ));
 sky130_fd_sc_hd__or2_1 \rpc/_436_  (.A(\rpc/_041_ ),
    .B(\rpc/_204_ ),
    .X(\rpc/_205_ ));
 sky130_fd_sc_hd__a31o_1 \rpc/_437_  (.A1(\rpc/_146_ ),
    .A2(\rpc/_189_ ),
    .A3(net336),
    .B1(net335),
    .X(\rpc/_206_ ));
 sky130_fd_sc_hd__a21o_1 \rpc/_438_  (.A1(net335),
    .A2(\rpc/_041_ ),
    .B1(\rpc/_047_ ),
    .X(\rpc/_207_ ));
 sky130_fd_sc_hd__nand3_1 \rpc/_439_  (.A(\rpc/_205_ ),
    .B(\rpc/_206_ ),
    .C(\rpc/_207_ ),
    .Y(\rpc/_208_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_440_  (.A(\rpc/_051_ ),
    .B(\wPcNextCond[27] ),
    .Y(\rpc/_209_ ));
 sky130_fd_sc_hd__a21oi_1 \rpc/_441_  (.A1(\rpc/_208_ ),
    .A2(\rpc/_209_ ),
    .B1(\rpc/_079_ ),
    .Y(\rpc/_025_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_442_  (.A(\rpc/_205_ ),
    .B(net333),
    .Y(\rpc/_210_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_443_  (.A(net333),
    .Y(\rpc/_211_ ));
 sky130_fd_sc_hd__nand3b_1 \rpc/_444_  (.A_N(\rpc/_204_ ),
    .B(\rpc/_211_ ),
    .C(\rpc/_033_ ),
    .Y(\rpc/_212_ ));
 sky130_fd_sc_hd__nand3_1 \rpc/_445_  (.A(\rpc/_210_ ),
    .B(\rpc/_060_ ),
    .C(\rpc/_212_ ),
    .Y(\rpc/_213_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_446_  (.A1(\wPcNextCond[28] ),
    .A2(\rpc/_059_ ),
    .B1(net1028),
    .X(\rpc/_214_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_447_  (.A(\rpc/_213_ ),
    .B(\rpc/_214_ ),
    .Y(\rpc/_215_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_448_  (.A(\rpc/_215_ ),
    .Y(\rpc/_026_ ));
 sky130_fd_sc_hd__and3_1 \rpc/_449_  (.A(\rpc/_203_ ),
    .B(net332),
    .C(net333),
    .X(\rpc/_216_ ));
 sky130_fd_sc_hd__nand3_2 \rpc/_450_  (.A(\rpc/_136_ ),
    .B(\rpc/_189_ ),
    .C(\rpc/_216_ ),
    .Y(\rpc/_217_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_451_  (.A(\rpc/_217_ ),
    .B(\rpc/_046_ ),
    .Y(\rpc/_218_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_452_  (.A(\rpc/_218_ ),
    .Y(\rpc/_219_ ));
 sky130_fd_sc_hd__nand3b_1 \rpc/_453_  (.A_N(\rpc/_204_ ),
    .B(net333),
    .C(\rpc/_219_ ),
    .Y(\rpc/_220_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_454_  (.A(\rpc/_218_ ),
    .B(\rpc/_111_ ),
    .Y(\rpc/_221_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_455_  (.A(\rpc/_221_ ),
    .B(net332),
    .Y(\rpc/_222_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_456_  (.A(\rpc/_051_ ),
    .B(\wPcNextCond[29] ),
    .Y(\rpc/_223_ ));
 sky130_fd_sc_hd__a31oi_1 \rpc/_457_  (.A1(\rpc/_220_ ),
    .A2(\rpc/_222_ ),
    .A3(\rpc/_223_ ),
    .B1(\rpc/_079_ ),
    .Y(\rpc/_027_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_458_  (.A(\rpc/_076_ ),
    .B(\wPcNextCond[30] ),
    .Y(\rpc/_224_ ));
 sky130_fd_sc_hd__o31a_1 \rpc/_459_  (.A1(net330),
    .A2(\rpc/_056_ ),
    .A3(\rpc/_217_ ),
    .B1(\rpc/_224_ ),
    .X(\rpc/_225_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_460_  (.A(\rpc/_221_ ),
    .B(net330),
    .Y(\rpc/_226_ ));
 sky130_fd_sc_hd__a21oi_1 \rpc/_461_  (.A1(\rpc/_225_ ),
    .A2(\rpc/_226_ ),
    .B1(\rpc/_079_ ),
    .Y(\rpc/_028_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_462_  (.A(net330),
    .Y(\rpc/_227_ ));
 sky130_fd_sc_hd__o21ai_1 \rpc/_463_  (.A1(\rpc/_227_ ),
    .A2(\rpc/_217_ ),
    .B1(net329),
    .Y(\rpc/_228_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_464_  (.A(\rpc/_217_ ),
    .Y(\rpc/_229_ ));
 sky130_fd_sc_hd__inv_2 \rpc/_465_  (.A(net329),
    .Y(\rpc/_230_ ));
 sky130_fd_sc_hd__nand3_1 \rpc/_466_  (.A(\rpc/_229_ ),
    .B(\rpc/_230_ ),
    .C(net330),
    .Y(\rpc/_231_ ));
 sky130_fd_sc_hd__nand3_1 \rpc/_467_  (.A(\rpc/_228_ ),
    .B(\rpc/_231_ ),
    .C(\rpc/_039_ ),
    .Y(\rpc/_232_ ));
 sky130_fd_sc_hd__o21a_1 \rpc/_468_  (.A1(\rpc/_039_ ),
    .A2(\wPcNextCond[31] ),
    .B1(\rpc/_111_ ),
    .X(\rpc/_233_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_469_  (.A(\rpc/_232_ ),
    .B(\rpc/_233_ ),
    .Y(\rpc/_234_ ));
 sky130_fd_sc_hd__nand2_1 \rpc/_470_  (.A(\rpc/_073_ ),
    .B(net329),
    .Y(\rpc/_235_ ));
 sky130_fd_sc_hd__a21oi_1 \rpc/_471_  (.A1(\rpc/_234_ ),
    .A2(\rpc/_235_ ),
    .B1(\rpc/_079_ ),
    .Y(\rpc/_029_ ));
 sky130_fd_sc_hd__or2_1 \rpc/_472_  (.A(\wPcNextCond[0] ),
    .B(\rpc/_048_ ),
    .X(\rpc/_236_ ));
 sky130_fd_sc_hd__o211a_1 \rpc/_473_  (.A1(net135),
    .A2(\rpc/_077_ ),
    .B1(net1029),
    .C1(\rpc/_236_ ),
    .X(\rpc/_030_ ));
 sky130_fd_sc_hd__or2_1 \rpc/_474_  (.A(\wPcNextCond[1] ),
    .B(\rpc/_048_ ),
    .X(\rpc/_237_ ));
 sky130_fd_sc_hd__o211a_1 \rpc/_475_  (.A1(net146),
    .A2(\rpc/_077_ ),
    .B1(net1030),
    .C1(\rpc/_237_ ),
    .X(\rpc/_031_ ));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_476_  (.CLK(clknet_leaf_50_clk),
    .D(\rpc/_000_ ),
    .Q(net157));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_477_  (.CLK(clknet_leaf_50_clk),
    .D(\rpc/_001_ ),
    .Q(net160));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_478_  (.CLK(clknet_leaf_53_clk),
    .D(\rpc/_002_ ),
    .Q(net161));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_479_  (.CLK(clknet_leaf_50_clk),
    .D(\rpc/_003_ ),
    .Q(net162));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_480_  (.CLK(clknet_leaf_52_clk),
    .D(\rpc/_004_ ),
    .Q(net163));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_481_  (.CLK(clknet_leaf_52_clk),
    .D(\rpc/_005_ ),
    .Q(net164));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_482_  (.CLK(clknet_leaf_50_clk),
    .D(\rpc/_006_ ),
    .Q(net165));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_483_  (.CLK(clknet_leaf_50_clk),
    .D(\rpc/_007_ ),
    .Q(net166));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_484_  (.CLK(clknet_leaf_51_clk),
    .D(\rpc/_008_ ),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_485_  (.CLK(clknet_leaf_39_clk),
    .D(\rpc/_009_ ),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_486_  (.CLK(clknet_leaf_48_clk),
    .D(\rpc/_010_ ),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_487_  (.CLK(clknet_leaf_39_clk),
    .D(\rpc/_011_ ),
    .Q(net139));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_488_  (.CLK(clknet_leaf_40_clk),
    .D(\rpc/_012_ ),
    .Q(net140));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_489_  (.CLK(clknet_leaf_39_clk),
    .D(\rpc/_013_ ),
    .Q(net141));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_490_  (.CLK(clknet_leaf_38_clk),
    .D(\rpc/_014_ ),
    .Q(net142));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_491_  (.CLK(clknet_leaf_49_clk),
    .D(\rpc/_015_ ),
    .Q(net143));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_492_  (.CLK(clknet_leaf_49_clk),
    .D(\rpc/_016_ ),
    .Q(net144));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_493_  (.CLK(clknet_leaf_39_clk),
    .D(\rpc/_017_ ),
    .Q(net145));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_494_  (.CLK(clknet_leaf_38_clk),
    .D(\rpc/_018_ ),
    .Q(net147));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_495_  (.CLK(clknet_leaf_38_clk),
    .D(\rpc/_019_ ),
    .Q(net148));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_496_  (.CLK(clknet_leaf_38_clk),
    .D(\rpc/_020_ ),
    .Q(net149));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_497_  (.CLK(clknet_leaf_38_clk),
    .D(\rpc/_021_ ),
    .Q(net150));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_498_  (.CLK(clknet_leaf_39_clk),
    .D(\rpc/_022_ ),
    .Q(net151));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_499_  (.CLK(clknet_leaf_38_clk),
    .D(\rpc/_023_ ),
    .Q(net152));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_500_  (.CLK(clknet_leaf_38_clk),
    .D(\rpc/_024_ ),
    .Q(net153));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_501_  (.CLK(clknet_leaf_49_clk),
    .D(\rpc/_025_ ),
    .Q(net154));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_502_  (.CLK(clknet_leaf_50_clk),
    .D(\rpc/_026_ ),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_503_  (.CLK(clknet_leaf_49_clk),
    .D(\rpc/_027_ ),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_504_  (.CLK(clknet_leaf_49_clk),
    .D(\rpc/_028_ ),
    .Q(net158));
 sky130_fd_sc_hd__dfxtp_1 \rpc/_505_  (.CLK(clknet_leaf_49_clk),
    .D(\rpc/_029_ ),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_2 \rpc/_506_  (.CLK(clknet_leaf_53_clk),
    .D(\rpc/_030_ ),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_2 \rpc/_507_  (.CLK(clknet_leaf_52_clk),
    .D(\rpc/_031_ ),
    .Q(net146));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Right_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Right_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Right_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Right_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Right_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Right_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Right_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Right_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Right_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Right_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Right_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Right_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Right_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Right_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Right_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Right_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Right_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Right_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Right_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Right_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Right_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Right_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Right_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Right_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Right_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Right_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Right_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Right_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Right_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Right_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Right_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Right_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Right_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Right_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Right_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Right_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Right_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Right_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Right_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Right_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Right_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Right_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Right_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Right_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Right_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Right_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Right_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Right_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Right_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Right_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Right_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Right_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Right_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Right_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Right_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Right_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Right_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Right_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Right_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Right_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Right_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Right_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Right_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Right_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Right_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Right_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Right_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Right_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Right_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Right_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Right_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Right_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Right_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Right_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Right_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Right_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Right_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Right_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Right_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Right_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Right_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Right_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Right_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Right_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Right_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Right_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Right_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Right_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Right_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Right_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Right_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Right_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Right_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Right_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Right_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Right_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Right_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Right_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Right_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Right_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_223 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_224 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_225 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_226 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_227 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_228 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_229 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_230 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_231 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_232 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_233 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_234 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_235 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_236 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_237 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_238 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_239 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_240 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_241 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_242 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_243 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_244 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_245 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_246 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_247 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_248 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_249 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_250 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_251 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_252 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_253 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_254 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_255 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_256 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_257 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_258 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_259 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_260 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_261 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_262 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_263 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_264 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_265 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_266 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_267 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_268 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_269 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_270 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_271 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_272 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_273 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_274 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_275 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_276 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_277 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_278 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_279 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_280 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_281 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_282 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_283 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_284 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_285 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_286 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_287 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_288 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_289 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_290 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_291 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_292 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_293 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_294 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_295 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_296 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_297 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_298 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_299 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_300 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_301 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_302 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_303 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_304 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_305 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_306 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_307 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_308 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_309 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_310 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_311 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_312 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_313 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_314 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_315 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_316 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_317 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_318 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_319 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_320 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_321 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_322 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_323 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_112_Left_324 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_113_Left_325 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_114_Left_326 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_115_Left_327 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_116_Left_328 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_117_Left_329 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_118_Left_330 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_119_Left_331 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_120_Left_332 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_121_Left_333 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_122_Left_334 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_123_Left_335 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_124_Left_336 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_125_Left_337 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_126_Left_338 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_127_Left_339 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_128_Left_340 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_129_Left_341 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_130_Left_342 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_131_Left_343 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_132_Left_344 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_133_Left_345 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_134_Left_346 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_135_Left_347 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_136_Left_348 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_137_Left_349 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_138_Left_350 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_139_Left_351 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_140_Left_352 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_141_Left_353 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_142_Left_354 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_143_Left_355 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_144_Left_356 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_145_Left_357 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_146_Left_358 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_147_Left_359 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_148_Left_360 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_149_Left_361 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_150_Left_362 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_151_Left_363 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_152_Left_364 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_153_Left_365 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_154_Left_366 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_155_Left_367 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_156_Left_368 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_157_Left_369 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_158_Left_370 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_159_Left_371 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_160_Left_372 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_161_Left_373 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_162_Left_374 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_163_Left_375 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_164_Left_376 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_165_Left_377 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_166_Left_378 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_167_Left_379 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_168_Left_380 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_169_Left_381 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_170_Left_382 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_171_Left_383 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_172_Left_384 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_173_Left_385 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_174_Left_386 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_175_Left_387 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_176_Left_388 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_177_Left_389 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_178_Left_390 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_179_Left_391 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_180_Left_392 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_181_Left_393 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_182_Left_394 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_183_Left_395 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_184_Left_396 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_185_Left_397 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_186_Left_398 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_187_Left_399 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_188_Left_400 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_189_Left_401 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_190_Left_402 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_191_Left_403 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_192_Left_404 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_193_Left_405 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_194_Left_406 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_195_Left_407 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_196_Left_408 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_197_Left_409 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_198_Left_410 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_199_Left_411 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_200_Left_412 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_201_Left_413 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_202_Left_414 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_203_Left_415 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_204_Left_416 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_205_Left_417 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_206_Left_418 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_207_Left_419 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_208_Left_420 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_209_Left_421 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_210_Left_422 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_211_Left_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_112_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_113_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_114_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_115_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_116_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_117_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_118_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_119_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_120_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_121_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_122_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_123_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_124_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_125_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_126_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_127_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_128_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_129_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_130_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_131_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_132_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_133_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_134_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_135_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_136_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_137_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_138_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_139_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_140_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_141_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_142_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_143_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_144_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_145_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_146_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_147_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_148_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_149_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_150_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_151_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_152_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_153_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_154_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_155_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_156_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_157_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_158_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_159_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_160_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_161_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_162_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_163_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_164_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_165_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_166_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_167_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_168_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_169_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_170_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_171_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_172_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_173_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_174_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_175_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_176_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_177_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_178_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_179_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_180_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_181_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_182_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_183_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_184_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_185_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_186_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_187_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_188_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_189_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_190_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_191_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_192_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_193_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_194_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_195_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_196_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_197_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_198_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_199_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_200_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_201_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_202_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_203_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_204_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_205_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_206_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_207_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_208_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_209_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_210_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_211_5131 ();
 sky130_fd_sc_hd__buf_1 input1 (.A(clkEn),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(dataBusIn[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input3 (.A(dataBusIn[10]),
    .X(net3));
 sky130_fd_sc_hd__buf_1 input4 (.A(dataBusIn[11]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(dataBusIn[12]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(dataBusIn[13]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input7 (.A(dataBusIn[14]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(dataBusIn[15]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(dataBusIn[16]),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(dataBusIn[17]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(dataBusIn[18]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(dataBusIn[19]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(dataBusIn[1]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(dataBusIn[20]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(dataBusIn[21]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(dataBusIn[22]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(dataBusIn[23]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(dataBusIn[24]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(dataBusIn[25]),
    .X(net19));
 sky130_fd_sc_hd__dlymetal6s2s_1 input20 (.A(dataBusIn[26]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(dataBusIn[27]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(dataBusIn[28]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(dataBusIn[29]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(dataBusIn[2]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(dataBusIn[30]),
    .X(net25));
 sky130_fd_sc_hd__buf_1 input26 (.A(dataBusIn[31]),
    .X(net26));
 sky130_fd_sc_hd__buf_1 input27 (.A(dataBusIn[3]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(dataBusIn[4]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(dataBusIn[5]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input30 (.A(dataBusIn[6]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(dataBusIn[7]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(dataBusIn[8]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(dataBusIn[9]),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 input34 (.A(inst_in[0]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(inst_in[10]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(inst_in[11]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(inst_in[12]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(inst_in[13]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(inst_in[14]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(inst_in[15]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(inst_in[16]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(inst_in[17]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(inst_in[18]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(inst_in[19]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(inst_in[1]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(inst_in[20]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(inst_in[21]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(inst_in[22]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(inst_in[23]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input50 (.A(inst_in[24]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(inst_in[25]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(inst_in[26]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(inst_in[27]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(inst_in[28]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(inst_in[29]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(inst_in[2]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(inst_in[30]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(inst_in[31]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(inst_in[3]),
    .X(net59));
 sky130_fd_sc_hd__dlymetal6s2s_1 input60 (.A(inst_in[4]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(inst_in[5]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(inst_in[6]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(inst_in[7]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(inst_in[8]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(inst_in[9]),
    .X(net65));
 sky130_fd_sc_hd__buf_1 input66 (.A(rstB),
    .X(net66));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(RamMode[0]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(RamMode[1]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(RamMode[2]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(RamMode[3]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(addr[0]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(addr[10]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(addr[11]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(addr[12]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(addr[13]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(addr[14]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(addr[15]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(addr[16]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(addr[17]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(addr[18]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(addr[19]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(addr[1]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(addr[20]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(addr[21]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(addr[22]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(addr[23]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(addr[24]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(addr[25]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(addr[26]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(addr[27]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(addr[28]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(addr[29]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(addr[2]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(addr[30]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(addr[31]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(addr[3]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(addr[4]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(addr[5]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(addr[6]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(addr[7]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(addr[8]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(addr[9]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(dataBusOut[0]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(dataBusOut[10]));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(dataBusOut[11]));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(dataBusOut[12]));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(dataBusOut[13]));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(dataBusOut[14]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(dataBusOut[15]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(dataBusOut[16]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(dataBusOut[17]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(dataBusOut[18]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(dataBusOut[19]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(dataBusOut[1]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(dataBusOut[20]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(dataBusOut[21]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(dataBusOut[22]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(dataBusOut[23]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(dataBusOut[24]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(dataBusOut[25]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(dataBusOut[26]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(dataBusOut[27]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(dataBusOut[28]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(dataBusOut[29]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(dataBusOut[2]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(dataBusOut[30]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(dataBusOut[31]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(dataBusOut[3]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(dataBusOut[4]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(dataBusOut[5]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(dataBusOut[6]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(dataBusOut[7]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(dataBusOut[8]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(dataBusOut[9]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(pc[0]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net368),
    .X(pc[10]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net366),
    .X(pc[11]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net363),
    .X(pc[12]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net362),
    .X(pc[13]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net360),
    .X(pc[14]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net357),
    .X(pc[15]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net354),
    .X(pc[16]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net352),
    .X(pc[17]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net350),
    .X(pc[18]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net348),
    .X(pc[19]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(pc[1]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net346),
    .X(pc[20]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net345),
    .X(pc[21]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net343),
    .X(pc[22]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net342),
    .X(pc[23]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net340),
    .X(pc[24]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net339),
    .X(pc[25]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net336),
    .X(pc[26]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net335),
    .X(pc[27]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net334),
    .X(pc[28]));
 sky130_fd_sc_hd__buf_2 output156 (.A(net332),
    .X(pc[29]));
 sky130_fd_sc_hd__buf_2 output157 (.A(net378),
    .X(pc[2]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net330),
    .X(pc[30]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net329),
    .X(pc[31]));
 sky130_fd_sc_hd__buf_2 output160 (.A(net377),
    .X(pc[3]));
 sky130_fd_sc_hd__buf_2 output161 (.A(net376),
    .X(pc[4]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net375),
    .X(pc[5]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net373),
    .X(pc[6]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net372),
    .X(pc[7]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net371),
    .X(pc[8]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net370),
    .X(pc[9]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(rdEn));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(wrEn));
 sky130_fd_sc_hd__buf_2 fanout169 (.A(net170),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 fanout170 (.A(net174),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_2 fanout171 (.A(net172),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 fanout172 (.A(net174),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_2 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout174 (.A(\wAluB[4] ),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_2 fanout175 (.A(net178),
    .X(net175));
 sky130_fd_sc_hd__buf_1 fanout176 (.A(net178),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_2 fanout177 (.A(net178),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 fanout178 (.A(net182),
    .X(net178));
 sky130_fd_sc_hd__buf_2 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 fanout180 (.A(net182),
    .X(net180));
 sky130_fd_sc_hd__buf_1 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__buf_1 fanout182 (.A(\wAluB[2] ),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 fanout183 (.A(net186),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_2 fanout184 (.A(net185),
    .X(net184));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__buf_1 fanout186 (.A(net189),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_2 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_2 fanout188 (.A(net189),
    .X(net188));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout189 (.A(\wAluB[2] ),
    .X(net189));
 sky130_fd_sc_hd__buf_2 fanout190 (.A(\wAluA[7] ),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 fanout191 (.A(\wAluA[1] ),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_2 fanout192 (.A(\wAluA[31] ),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_2 fanout193 (.A(\wAluA[22] ),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 fanout194 (.A(\wAluA[8] ),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_2 fanout195 (.A(net200),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__buf_2 fanout197 (.A(net200),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 fanout199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__buf_1 fanout200 (.A(net207),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_2 fanout201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_2 fanout202 (.A(net207),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 fanout203 (.A(net206),
    .X(net203));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout204 (.A(net206),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_2 fanout205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_1 fanout207 (.A(\wAluB[3] ),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_2 fanout208 (.A(net209),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 fanout209 (.A(net213),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout213 (.A(net221),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 fanout214 (.A(net216),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_2 fanout215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 fanout216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__buf_1 fanout217 (.A(net221),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_2 fanout218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 fanout219 (.A(net220),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__buf_1 fanout221 (.A(\wAluB[1] ),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_2 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__buf_2 fanout224 (.A(net235),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 fanout225 (.A(net228),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_2 fanout226 (.A(net227),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_2 fanout228 (.A(net235),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_2 fanout229 (.A(net232),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_2 fanout230 (.A(net232),
    .X(net230));
 sky130_fd_sc_hd__buf_1 fanout231 (.A(net232),
    .X(net231));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 fanout234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_2 fanout235 (.A(\wAluB[0] ),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 fanout236 (.A(\wAluA[28] ),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_2 fanout237 (.A(\wAluA[11] ),
    .X(net237));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout238 (.A(net240),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_2 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__buf_1 fanout240 (.A(net242),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 fanout242 (.A(net250),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 fanout243 (.A(net245),
    .X(net243));
 sky130_fd_sc_hd__buf_1 fanout244 (.A(net245),
    .X(net244));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout245 (.A(net250),
    .X(net245));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout246 (.A(net249),
    .X(net246));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout247 (.A(net249),
    .X(net247));
 sky130_fd_sc_hd__buf_1 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 fanout249 (.A(net250),
    .X(net249));
 sky130_fd_sc_hd__buf_1 fanout250 (.A(net259),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_2 fanout251 (.A(net253),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_2 fanout252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 fanout253 (.A(net257),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_2 fanout254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_2 fanout255 (.A(net256),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_2 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_2 fanout257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__buf_2 fanout258 (.A(net259),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 fanout259 (.A(net279),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_2 fanout260 (.A(net262),
    .X(net260));
 sky130_fd_sc_hd__buf_1 fanout261 (.A(net262),
    .X(net261));
 sky130_fd_sc_hd__buf_1 fanout262 (.A(net264),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__buf_1 fanout264 (.A(net270),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_2 fanout265 (.A(net268),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_2 fanout266 (.A(net267),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_2 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 fanout268 (.A(net270),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_2 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__buf_1 fanout270 (.A(net279),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_2 fanout271 (.A(net273),
    .X(net271));
 sky130_fd_sc_hd__buf_1 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__buf_1 fanout273 (.A(net278),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_2 fanout274 (.A(net278),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_2 fanout275 (.A(net276),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_2 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_2 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__buf_1 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_2 fanout279 (.A(wStall),
    .X(net279));
 sky130_fd_sc_hd__buf_1 wire280 (.A(\reg_module/_09687_ ),
    .X(net280));
 sky130_fd_sc_hd__buf_1 wire281 (.A(\reg_module/_08606_ ),
    .X(net281));
 sky130_fd_sc_hd__buf_1 wire282 (.A(\reg_module/_08603_ ),
    .X(net282));
 sky130_fd_sc_hd__buf_1 wire283 (.A(\reg_module/_08547_ ),
    .X(net283));
 sky130_fd_sc_hd__buf_1 wire284 (.A(\reg_module/_08542_ ),
    .X(net284));
 sky130_fd_sc_hd__buf_1 wire285 (.A(\reg_module/_08534_ ),
    .X(net285));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap286 (.A(_0208_),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_2 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_4 fanout288 (.A(\wRegWrData[31] ),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_2 fanout289 (.A(\wRegWrData[30] ),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_2 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__buf_2 fanout291 (.A(\wRegWrData[29] ),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_2 fanout292 (.A(\wRegWrData[28] ),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_2 fanout293 (.A(\wRegWrData[27] ),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_2 fanout294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__buf_2 fanout295 (.A(\wRegWrData[26] ),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_2 fanout296 (.A(net297),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 fanout297 (.A(\wRegWrData[25] ),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_2 fanout298 (.A(\wRegWrData[24] ),
    .X(net298));
 sky130_fd_sc_hd__buf_2 fanout299 (.A(\wRegWrData[23] ),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_4 fanout300 (.A(\wRegWrData[22] ),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_4 fanout301 (.A(\wRegWrData[21] ),
    .X(net301));
 sky130_fd_sc_hd__buf_2 fanout302 (.A(\wRegWrData[20] ),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_4 fanout303 (.A(\wRegWrData[19] ),
    .X(net303));
 sky130_fd_sc_hd__buf_2 fanout304 (.A(\wRegWrData[18] ),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_4 fanout305 (.A(\wRegWrData[17] ),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_4 fanout306 (.A(\wRegWrData[15] ),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_2 fanout307 (.A(\wRegWrData[15] ),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_4 fanout308 (.A(\wRegWrData[14] ),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_4 fanout309 (.A(\wRegWrData[13] ),
    .X(net309));
 sky130_fd_sc_hd__buf_2 fanout310 (.A(\wRegWrData[11] ),
    .X(net310));
 sky130_fd_sc_hd__buf_2 fanout311 (.A(\wRegWrData[10] ),
    .X(net311));
 sky130_fd_sc_hd__buf_2 fanout312 (.A(\wRegWrData[9] ),
    .X(net312));
 sky130_fd_sc_hd__buf_2 fanout313 (.A(\wRegWrData[7] ),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_4 fanout314 (.A(\wRegWrData[5] ),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_4 fanout315 (.A(\wRegWrData[3] ),
    .X(net315));
 sky130_fd_sc_hd__buf_2 fanout316 (.A(\wRegWrData[2] ),
    .X(net316));
 sky130_fd_sc_hd__buf_2 fanout317 (.A(\wRegWrData[1] ),
    .X(net317));
 sky130_fd_sc_hd__buf_2 fanout318 (.A(net319),
    .X(net318));
 sky130_fd_sc_hd__buf_2 fanout319 (.A(\wRegWrData[0] ),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_2 fanout320 (.A(net328),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_2 fanout321 (.A(net327),
    .X(net321));
 sky130_fd_sc_hd__buf_1 fanout322 (.A(net327),
    .X(net322));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout323 (.A(net324),
    .X(net323));
 sky130_fd_sc_hd__buf_1 fanout324 (.A(net325),
    .X(net324));
 sky130_fd_sc_hd__buf_1 fanout325 (.A(net326),
    .X(net325));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout326 (.A(net327),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_2 fanout327 (.A(net328),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_2 fanout328 (.A(op_jal),
    .X(net328));
 sky130_fd_sc_hd__clkbuf_2 fanout329 (.A(net159),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_2 fanout330 (.A(net331),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_2 fanout331 (.A(net158),
    .X(net331));
 sky130_fd_sc_hd__buf_2 fanout332 (.A(net156),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_2 fanout333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_1 fanout334 (.A(net155),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_2 fanout335 (.A(net154),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_2 fanout336 (.A(net337),
    .X(net336));
 sky130_fd_sc_hd__buf_1 fanout337 (.A(net338),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_2 fanout338 (.A(net153),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_2 fanout339 (.A(net152),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_2 fanout340 (.A(net341),
    .X(net340));
 sky130_fd_sc_hd__buf_2 fanout341 (.A(net151),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_4 fanout342 (.A(net150),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 fanout343 (.A(net344),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_2 fanout344 (.A(net149),
    .X(net344));
 sky130_fd_sc_hd__buf_2 fanout345 (.A(net148),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_2 fanout346 (.A(net347),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_2 fanout347 (.A(net147),
    .X(net347));
 sky130_fd_sc_hd__buf_2 fanout348 (.A(net349),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_2 fanout349 (.A(net145),
    .X(net349));
 sky130_fd_sc_hd__buf_2 fanout350 (.A(net351),
    .X(net350));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout351 (.A(net144),
    .X(net351));
 sky130_fd_sc_hd__buf_2 fanout352 (.A(net353),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_2 fanout353 (.A(net143),
    .X(net353));
 sky130_fd_sc_hd__buf_2 fanout354 (.A(net356),
    .X(net354));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout355 (.A(net356),
    .X(net355));
 sky130_fd_sc_hd__buf_2 fanout356 (.A(net142),
    .X(net356));
 sky130_fd_sc_hd__buf_2 fanout357 (.A(net359),
    .X(net357));
 sky130_fd_sc_hd__buf_1 fanout358 (.A(net359),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_2 fanout359 (.A(net141),
    .X(net359));
 sky130_fd_sc_hd__buf_2 fanout360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_2 fanout361 (.A(net140),
    .X(net361));
 sky130_fd_sc_hd__buf_2 fanout362 (.A(net139),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_4 fanout363 (.A(net365),
    .X(net363));
 sky130_fd_sc_hd__buf_1 fanout364 (.A(net365),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_2 fanout365 (.A(net138),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_2 fanout366 (.A(net367),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_2 fanout367 (.A(net137),
    .X(net367));
 sky130_fd_sc_hd__buf_2 fanout368 (.A(net369),
    .X(net368));
 sky130_fd_sc_hd__buf_2 fanout369 (.A(net136),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_4 fanout370 (.A(net166),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_4 fanout371 (.A(net165),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_4 fanout372 (.A(net164),
    .X(net372));
 sky130_fd_sc_hd__buf_2 fanout373 (.A(net163),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_2 fanout374 (.A(net163),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_4 fanout375 (.A(net162),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_4 fanout376 (.A(net161),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_4 fanout377 (.A(net160),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_2 fanout378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_2 fanout379 (.A(net157),
    .X(net379));
 sky130_fd_sc_hd__buf_2 fanout380 (.A(net381),
    .X(net380));
 sky130_fd_sc_hd__buf_2 fanout381 (.A(net387),
    .X(net381));
 sky130_fd_sc_hd__buf_2 fanout382 (.A(net387),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_4 fanout383 (.A(net386),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_2 fanout384 (.A(net385),
    .X(net384));
 sky130_fd_sc_hd__buf_2 fanout385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_2 fanout386 (.A(net387),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_4 fanout387 (.A(\reg_module/rRs2[4] ),
    .X(net387));
 sky130_fd_sc_hd__buf_2 fanout388 (.A(net395),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_2 fanout389 (.A(net390),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_4 fanout390 (.A(net395),
    .X(net390));
 sky130_fd_sc_hd__buf_2 fanout391 (.A(net393),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_1 fanout392 (.A(net393),
    .X(net392));
 sky130_fd_sc_hd__buf_2 fanout393 (.A(net394),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_4 fanout394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_4 fanout395 (.A(\reg_module/rRs2[3] ),
    .X(net395));
 sky130_fd_sc_hd__buf_2 fanout396 (.A(net398),
    .X(net396));
 sky130_fd_sc_hd__buf_1 fanout397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_4 fanout398 (.A(net404),
    .X(net398));
 sky130_fd_sc_hd__buf_2 fanout399 (.A(net403),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_2 fanout400 (.A(net403),
    .X(net400));
 sky130_fd_sc_hd__buf_2 fanout401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__buf_2 fanout402 (.A(net403),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_2 fanout403 (.A(net404),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_4 fanout404 (.A(\reg_module/rRs2[3] ),
    .X(net404));
 sky130_fd_sc_hd__buf_2 fanout405 (.A(net412),
    .X(net405));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout406 (.A(net412),
    .X(net406));
 sky130_fd_sc_hd__buf_2 fanout407 (.A(net411),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_2 fanout408 (.A(net411),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_2 fanout409 (.A(net411),
    .X(net409));
 sky130_fd_sc_hd__buf_1 fanout410 (.A(net411),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_2 fanout411 (.A(net412),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_2 fanout412 (.A(net439),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_2 fanout413 (.A(net420),
    .X(net413));
 sky130_fd_sc_hd__buf_1 fanout414 (.A(net420),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_2 fanout415 (.A(net416),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_2 fanout416 (.A(net418),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_2 fanout417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout418 (.A(net419),
    .X(net418));
 sky130_fd_sc_hd__clkbuf_2 fanout419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_2 fanout420 (.A(net439),
    .X(net420));
 sky130_fd_sc_hd__buf_2 fanout421 (.A(net423),
    .X(net421));
 sky130_fd_sc_hd__buf_1 fanout422 (.A(net423),
    .X(net422));
 sky130_fd_sc_hd__buf_2 fanout423 (.A(net427),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_2 fanout424 (.A(net427),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_2 fanout425 (.A(net426),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_4 fanout426 (.A(net427),
    .X(net426));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout427 (.A(net438),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_2 fanout428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__clkbuf_2 fanout429 (.A(net430),
    .X(net429));
 sky130_fd_sc_hd__buf_2 fanout430 (.A(net438),
    .X(net430));
 sky130_fd_sc_hd__buf_2 fanout431 (.A(net437),
    .X(net431));
 sky130_fd_sc_hd__buf_1 fanout432 (.A(net437),
    .X(net432));
 sky130_fd_sc_hd__buf_2 fanout433 (.A(net436),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_2 fanout434 (.A(net436),
    .X(net434));
 sky130_fd_sc_hd__buf_1 fanout435 (.A(net436),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_2 fanout436 (.A(net437),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_2 fanout437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__buf_2 fanout438 (.A(net439),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_4 fanout439 (.A(\reg_module/rRs2[2] ),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_2 fanout440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__buf_1 fanout441 (.A(net445),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_2 fanout442 (.A(net444),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_2 fanout443 (.A(net444),
    .X(net443));
 sky130_fd_sc_hd__buf_2 fanout444 (.A(net445),
    .X(net444));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout445 (.A(net453),
    .X(net445));
 sky130_fd_sc_hd__clkbuf_2 fanout446 (.A(net449),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_2 fanout447 (.A(net449),
    .X(net447));
 sky130_fd_sc_hd__buf_1 fanout448 (.A(net449),
    .X(net448));
 sky130_fd_sc_hd__clkbuf_2 fanout449 (.A(net453),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_2 fanout450 (.A(net452),
    .X(net450));
 sky130_fd_sc_hd__clkbuf_2 fanout451 (.A(net452),
    .X(net451));
 sky130_fd_sc_hd__buf_2 fanout452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_2 fanout453 (.A(net468),
    .X(net453));
 sky130_fd_sc_hd__buf_2 fanout454 (.A(net455),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_2 fanout455 (.A(net457),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_2 fanout456 (.A(net457),
    .X(net456));
 sky130_fd_sc_hd__buf_1 fanout457 (.A(net459),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_2 fanout458 (.A(net459),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_2 fanout459 (.A(net468),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_2 fanout460 (.A(net467),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_2 fanout461 (.A(net467),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_2 fanout462 (.A(net467),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_2 fanout463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_2 fanout464 (.A(net467),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_2 fanout465 (.A(net466),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_2 fanout466 (.A(net467),
    .X(net466));
 sky130_fd_sc_hd__buf_2 fanout467 (.A(net468),
    .X(net467));
 sky130_fd_sc_hd__buf_2 fanout468 (.A(net504),
    .X(net468));
 sky130_fd_sc_hd__buf_2 fanout469 (.A(net473),
    .X(net469));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout470 (.A(net473),
    .X(net470));
 sky130_fd_sc_hd__clkbuf_2 fanout471 (.A(net473),
    .X(net471));
 sky130_fd_sc_hd__buf_1 fanout472 (.A(net473),
    .X(net472));
 sky130_fd_sc_hd__clkbuf_2 fanout473 (.A(net484),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_2 fanout474 (.A(net477),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_2 fanout475 (.A(net477),
    .X(net475));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout476 (.A(net477),
    .X(net476));
 sky130_fd_sc_hd__buf_2 fanout477 (.A(net484),
    .X(net477));
 sky130_fd_sc_hd__buf_2 fanout478 (.A(net479),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_2 fanout479 (.A(net484),
    .X(net479));
 sky130_fd_sc_hd__buf_2 fanout480 (.A(net483),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_2 fanout481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_2 fanout482 (.A(net483),
    .X(net482));
 sky130_fd_sc_hd__clkbuf_2 fanout483 (.A(net484),
    .X(net483));
 sky130_fd_sc_hd__buf_2 fanout484 (.A(net504),
    .X(net484));
 sky130_fd_sc_hd__buf_2 fanout485 (.A(net488),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_2 fanout486 (.A(net488),
    .X(net486));
 sky130_fd_sc_hd__buf_1 fanout487 (.A(net488),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_2 fanout488 (.A(net503),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_2 fanout489 (.A(net490),
    .X(net489));
 sky130_fd_sc_hd__buf_2 fanout490 (.A(net493),
    .X(net490));
 sky130_fd_sc_hd__buf_2 fanout491 (.A(net493),
    .X(net491));
 sky130_fd_sc_hd__buf_1 fanout492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__buf_1 fanout493 (.A(net503),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_2 fanout494 (.A(net497),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_2 fanout495 (.A(net497),
    .X(net495));
 sky130_fd_sc_hd__buf_1 fanout496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_2 fanout497 (.A(net503),
    .X(net497));
 sky130_fd_sc_hd__clkbuf_2 fanout498 (.A(net502),
    .X(net498));
 sky130_fd_sc_hd__buf_1 fanout499 (.A(net502),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_2 fanout500 (.A(net502),
    .X(net500));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout501 (.A(net502),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_2 fanout502 (.A(net503),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_4 fanout503 (.A(net504),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_4 fanout504 (.A(\reg_module/rRs2[1] ),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_2 fanout505 (.A(net506),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_2 fanout506 (.A(net507),
    .X(net506));
 sky130_fd_sc_hd__clkbuf_2 fanout507 (.A(net515),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_2 fanout508 (.A(net509),
    .X(net508));
 sky130_fd_sc_hd__clkbuf_2 fanout509 (.A(net512),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_2 fanout510 (.A(net511),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_2 fanout511 (.A(net512),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_2 fanout512 (.A(net515),
    .X(net512));
 sky130_fd_sc_hd__clkbuf_2 fanout513 (.A(net514),
    .X(net513));
 sky130_fd_sc_hd__buf_1 fanout514 (.A(net515),
    .X(net514));
 sky130_fd_sc_hd__buf_2 fanout515 (.A(net560),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_2 fanout516 (.A(net518),
    .X(net516));
 sky130_fd_sc_hd__buf_1 fanout517 (.A(net518),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_2 fanout518 (.A(net524),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_2 fanout519 (.A(net523),
    .X(net519));
 sky130_fd_sc_hd__buf_1 fanout520 (.A(net521),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_2 fanout521 (.A(net523),
    .X(net521));
 sky130_fd_sc_hd__clkbuf_2 fanout522 (.A(net523),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_2 fanout523 (.A(net524),
    .X(net523));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout524 (.A(net532),
    .X(net524));
 sky130_fd_sc_hd__clkbuf_2 fanout525 (.A(net528),
    .X(net525));
 sky130_fd_sc_hd__buf_1 fanout526 (.A(net528),
    .X(net526));
 sky130_fd_sc_hd__clkbuf_2 fanout527 (.A(net528),
    .X(net527));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout528 (.A(net532),
    .X(net528));
 sky130_fd_sc_hd__clkbuf_2 fanout529 (.A(net531),
    .X(net529));
 sky130_fd_sc_hd__buf_1 fanout530 (.A(net531),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_2 fanout531 (.A(net532),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_2 fanout532 (.A(net560),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_2 fanout533 (.A(net535),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_2 fanout534 (.A(net535),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_2 fanout535 (.A(net538),
    .X(net535));
 sky130_fd_sc_hd__clkbuf_2 fanout536 (.A(net538),
    .X(net536));
 sky130_fd_sc_hd__clkbuf_2 fanout537 (.A(net538),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_2 fanout538 (.A(net542),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_2 fanout539 (.A(net542),
    .X(net539));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout540 (.A(net541),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_2 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_2 fanout542 (.A(net560),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_2 fanout543 (.A(net545),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_2 fanout544 (.A(net545),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_2 fanout545 (.A(net559),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_2 fanout546 (.A(net547),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_2 fanout547 (.A(net550),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_2 fanout548 (.A(net550),
    .X(net548));
 sky130_fd_sc_hd__buf_1 fanout549 (.A(net550),
    .X(net549));
 sky130_fd_sc_hd__buf_1 fanout550 (.A(net559),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_2 fanout551 (.A(net552),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_2 fanout552 (.A(net554),
    .X(net552));
 sky130_fd_sc_hd__buf_1 fanout553 (.A(net554),
    .X(net553));
 sky130_fd_sc_hd__clkbuf_2 fanout554 (.A(net559),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_2 fanout555 (.A(net556),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_2 fanout556 (.A(net558),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_2 fanout557 (.A(net558),
    .X(net557));
 sky130_fd_sc_hd__buf_1 fanout558 (.A(net559),
    .X(net558));
 sky130_fd_sc_hd__buf_2 fanout559 (.A(net560),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_4 fanout560 (.A(\reg_module/rRs2[0] ),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_2 fanout561 (.A(net564),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_2 fanout562 (.A(net564),
    .X(net562));
 sky130_fd_sc_hd__buf_1 fanout563 (.A(net564),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_2 fanout564 (.A(net578),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_2 fanout565 (.A(net569),
    .X(net565));
 sky130_fd_sc_hd__buf_1 fanout566 (.A(net569),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_2 fanout567 (.A(net569),
    .X(net567));
 sky130_fd_sc_hd__buf_1 fanout568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout569 (.A(net578),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_2 fanout570 (.A(net571),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_2 fanout571 (.A(net577),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_2 fanout572 (.A(net576),
    .X(net572));
 sky130_fd_sc_hd__buf_1 fanout573 (.A(net576),
    .X(net573));
 sky130_fd_sc_hd__clkbuf_2 fanout574 (.A(net576),
    .X(net574));
 sky130_fd_sc_hd__buf_1 fanout575 (.A(net576),
    .X(net575));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout576 (.A(net577),
    .X(net576));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout577 (.A(net578),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_2 fanout578 (.A(net631),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_2 fanout579 (.A(net582),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_2 fanout580 (.A(net582),
    .X(net580));
 sky130_fd_sc_hd__buf_1 fanout581 (.A(net582),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_2 fanout582 (.A(net583),
    .X(net582));
 sky130_fd_sc_hd__buf_2 fanout583 (.A(net592),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_2 fanout584 (.A(net586),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_1 fanout585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_2 fanout586 (.A(net591),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_2 fanout587 (.A(net588),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_2 fanout588 (.A(net591),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_2 fanout589 (.A(net590),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_2 fanout590 (.A(net591),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_2 fanout591 (.A(net592),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_2 fanout592 (.A(net631),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_2 fanout593 (.A(net594),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_2 fanout594 (.A(net601),
    .X(net594));
 sky130_fd_sc_hd__buf_1 fanout595 (.A(net601),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_2 fanout596 (.A(net600),
    .X(net596));
 sky130_fd_sc_hd__buf_1 fanout597 (.A(net600),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_2 fanout598 (.A(net599),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_2 fanout599 (.A(net600),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_2 fanout600 (.A(net601),
    .X(net600));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout601 (.A(net611),
    .X(net601));
 sky130_fd_sc_hd__clkbuf_2 fanout602 (.A(net606),
    .X(net602));
 sky130_fd_sc_hd__buf_1 fanout603 (.A(net606),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_2 fanout604 (.A(net606),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_2 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_2 fanout606 (.A(net611),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_2 fanout607 (.A(net610),
    .X(net607));
 sky130_fd_sc_hd__buf_1 fanout608 (.A(net610),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_2 fanout609 (.A(net610),
    .X(net609));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout610 (.A(net611),
    .X(net610));
 sky130_fd_sc_hd__clkbuf_2 fanout611 (.A(net631),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_2 fanout612 (.A(net613),
    .X(net612));
 sky130_fd_sc_hd__buf_1 fanout613 (.A(net614),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_2 fanout614 (.A(net621),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_2 fanout615 (.A(net620),
    .X(net615));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout616 (.A(net620),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_2 fanout617 (.A(net619),
    .X(net617));
 sky130_fd_sc_hd__buf_1 fanout618 (.A(net619),
    .X(net618));
 sky130_fd_sc_hd__clkbuf_2 fanout619 (.A(net620),
    .X(net619));
 sky130_fd_sc_hd__buf_1 fanout620 (.A(net621),
    .X(net620));
 sky130_fd_sc_hd__buf_1 fanout621 (.A(net630),
    .X(net621));
 sky130_fd_sc_hd__clkbuf_2 fanout622 (.A(net623),
    .X(net622));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout623 (.A(net625),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_2 fanout624 (.A(net625),
    .X(net624));
 sky130_fd_sc_hd__buf_1 fanout625 (.A(net630),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_2 fanout626 (.A(net629),
    .X(net626));
 sky130_fd_sc_hd__clkbuf_2 fanout627 (.A(net629),
    .X(net627));
 sky130_fd_sc_hd__clkbuf_2 fanout628 (.A(net629),
    .X(net628));
 sky130_fd_sc_hd__clkbuf_2 fanout629 (.A(net630),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_2 fanout630 (.A(net631),
    .X(net630));
 sky130_fd_sc_hd__clkbuf_4 fanout631 (.A(\reg_module/rRs2[0] ),
    .X(net631));
 sky130_fd_sc_hd__buf_2 fanout632 (.A(net635),
    .X(net632));
 sky130_fd_sc_hd__buf_2 fanout633 (.A(net635),
    .X(net633));
 sky130_fd_sc_hd__buf_1 fanout634 (.A(net635),
    .X(net634));
 sky130_fd_sc_hd__buf_4 fanout635 (.A(net639),
    .X(net635));
 sky130_fd_sc_hd__buf_2 fanout636 (.A(net637),
    .X(net636));
 sky130_fd_sc_hd__buf_2 fanout637 (.A(net639),
    .X(net637));
 sky130_fd_sc_hd__clkbuf_4 fanout638 (.A(net639),
    .X(net638));
 sky130_fd_sc_hd__buf_2 fanout639 (.A(\reg_module/rRs1[4] ),
    .X(net639));
 sky130_fd_sc_hd__buf_2 fanout640 (.A(net641),
    .X(net640));
 sky130_fd_sc_hd__clkbuf_2 fanout641 (.A(net642),
    .X(net641));
 sky130_fd_sc_hd__clkbuf_4 fanout642 (.A(net655),
    .X(net642));
 sky130_fd_sc_hd__clkbuf_2 fanout643 (.A(net645),
    .X(net643));
 sky130_fd_sc_hd__buf_1 fanout644 (.A(net645),
    .X(net644));
 sky130_fd_sc_hd__buf_2 fanout645 (.A(net646),
    .X(net645));
 sky130_fd_sc_hd__clkbuf_4 fanout646 (.A(net655),
    .X(net646));
 sky130_fd_sc_hd__buf_2 fanout647 (.A(net648),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_2 fanout648 (.A(net650),
    .X(net648));
 sky130_fd_sc_hd__buf_2 fanout649 (.A(net650),
    .X(net649));
 sky130_fd_sc_hd__clkbuf_2 fanout650 (.A(net654),
    .X(net650));
 sky130_fd_sc_hd__buf_2 fanout651 (.A(net652),
    .X(net651));
 sky130_fd_sc_hd__clkbuf_4 fanout652 (.A(net654),
    .X(net652));
 sky130_fd_sc_hd__buf_2 fanout653 (.A(net654),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_4 fanout654 (.A(net655),
    .X(net654));
 sky130_fd_sc_hd__clkbuf_4 fanout655 (.A(\reg_module/rRs1[3] ),
    .X(net655));
 sky130_fd_sc_hd__buf_2 fanout656 (.A(net662),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_2 fanout657 (.A(net662),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_2 fanout658 (.A(net659),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_2 fanout659 (.A(net661),
    .X(net659));
 sky130_fd_sc_hd__buf_2 fanout660 (.A(net661),
    .X(net660));
 sky130_fd_sc_hd__buf_2 fanout661 (.A(net662),
    .X(net661));
 sky130_fd_sc_hd__clkbuf_2 fanout662 (.A(net688),
    .X(net662));
 sky130_fd_sc_hd__buf_2 fanout663 (.A(net670),
    .X(net663));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout664 (.A(net670),
    .X(net664));
 sky130_fd_sc_hd__clkbuf_2 fanout665 (.A(net668),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_2 fanout666 (.A(net667),
    .X(net666));
 sky130_fd_sc_hd__clkbuf_2 fanout667 (.A(net668),
    .X(net667));
 sky130_fd_sc_hd__clkbuf_2 fanout668 (.A(net669),
    .X(net668));
 sky130_fd_sc_hd__buf_2 fanout669 (.A(net670),
    .X(net669));
 sky130_fd_sc_hd__clkbuf_2 fanout670 (.A(net688),
    .X(net670));
 sky130_fd_sc_hd__buf_2 fanout671 (.A(net672),
    .X(net671));
 sky130_fd_sc_hd__clkbuf_2 fanout672 (.A(net673),
    .X(net672));
 sky130_fd_sc_hd__clkbuf_2 fanout673 (.A(net677),
    .X(net673));
 sky130_fd_sc_hd__buf_2 fanout674 (.A(net675),
    .X(net674));
 sky130_fd_sc_hd__buf_2 fanout675 (.A(net676),
    .X(net675));
 sky130_fd_sc_hd__buf_2 fanout676 (.A(net677),
    .X(net676));
 sky130_fd_sc_hd__buf_2 fanout677 (.A(net688),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_2 fanout678 (.A(net687),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_2 fanout679 (.A(net686),
    .X(net679));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout680 (.A(net686),
    .X(net680));
 sky130_fd_sc_hd__clkbuf_2 fanout681 (.A(net685),
    .X(net681));
 sky130_fd_sc_hd__buf_1 fanout682 (.A(net685),
    .X(net682));
 sky130_fd_sc_hd__clkbuf_2 fanout683 (.A(net684),
    .X(net683));
 sky130_fd_sc_hd__clkbuf_2 fanout684 (.A(net685),
    .X(net684));
 sky130_fd_sc_hd__buf_1 fanout685 (.A(net686),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_2 fanout686 (.A(net687),
    .X(net686));
 sky130_fd_sc_hd__clkbuf_2 fanout687 (.A(net688),
    .X(net687));
 sky130_fd_sc_hd__buf_4 fanout688 (.A(\reg_module/rRs1[2] ),
    .X(net688));
 sky130_fd_sc_hd__clkbuf_2 fanout689 (.A(net690),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_2 fanout690 (.A(net701),
    .X(net690));
 sky130_fd_sc_hd__buf_2 fanout691 (.A(net693),
    .X(net691));
 sky130_fd_sc_hd__clkbuf_2 fanout692 (.A(net693),
    .X(net692));
 sky130_fd_sc_hd__buf_2 fanout693 (.A(net701),
    .X(net693));
 sky130_fd_sc_hd__clkbuf_2 fanout694 (.A(net697),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_2 fanout695 (.A(net697),
    .X(net695));
 sky130_fd_sc_hd__clkbuf_2 fanout696 (.A(net697),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_2 fanout697 (.A(net701),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_2 fanout698 (.A(net700),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_2 fanout699 (.A(net700),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_2 fanout700 (.A(net701),
    .X(net700));
 sky130_fd_sc_hd__buf_2 fanout701 (.A(net753),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_2 fanout702 (.A(net705),
    .X(net702));
 sky130_fd_sc_hd__buf_1 fanout703 (.A(net705),
    .X(net703));
 sky130_fd_sc_hd__clkbuf_2 fanout704 (.A(net705),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_2 fanout705 (.A(net707),
    .X(net705));
 sky130_fd_sc_hd__buf_2 fanout706 (.A(net707),
    .X(net706));
 sky130_fd_sc_hd__clkbuf_2 fanout707 (.A(net716),
    .X(net707));
 sky130_fd_sc_hd__buf_2 fanout708 (.A(net711),
    .X(net708));
 sky130_fd_sc_hd__clkbuf_2 fanout709 (.A(net711),
    .X(net709));
 sky130_fd_sc_hd__clkbuf_2 fanout710 (.A(net711),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_2 fanout711 (.A(net716),
    .X(net711));
 sky130_fd_sc_hd__clkbuf_2 fanout712 (.A(net715),
    .X(net712));
 sky130_fd_sc_hd__clkbuf_2 fanout713 (.A(net715),
    .X(net713));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout714 (.A(net715),
    .X(net714));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout715 (.A(net716),
    .X(net715));
 sky130_fd_sc_hd__clkbuf_2 fanout716 (.A(net753),
    .X(net716));
 sky130_fd_sc_hd__buf_2 fanout717 (.A(net721),
    .X(net717));
 sky130_fd_sc_hd__buf_1 fanout718 (.A(net721),
    .X(net718));
 sky130_fd_sc_hd__clkbuf_2 fanout719 (.A(net721),
    .X(net719));
 sky130_fd_sc_hd__buf_1 fanout720 (.A(net721),
    .X(net720));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout721 (.A(net734),
    .X(net721));
 sky130_fd_sc_hd__clkbuf_2 fanout722 (.A(net726),
    .X(net722));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout723 (.A(net726),
    .X(net723));
 sky130_fd_sc_hd__clkbuf_2 fanout724 (.A(net725),
    .X(net724));
 sky130_fd_sc_hd__buf_2 fanout725 (.A(net726),
    .X(net725));
 sky130_fd_sc_hd__buf_1 fanout726 (.A(net734),
    .X(net726));
 sky130_fd_sc_hd__clkbuf_2 fanout727 (.A(net728),
    .X(net727));
 sky130_fd_sc_hd__buf_2 fanout728 (.A(net734),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_2 fanout729 (.A(net733),
    .X(net729));
 sky130_fd_sc_hd__buf_1 fanout730 (.A(net733),
    .X(net730));
 sky130_fd_sc_hd__clkbuf_2 fanout731 (.A(net733),
    .X(net731));
 sky130_fd_sc_hd__buf_1 fanout732 (.A(net733),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_2 fanout733 (.A(net734),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_4 fanout734 (.A(net753),
    .X(net734));
 sky130_fd_sc_hd__buf_2 fanout735 (.A(net738),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_2 fanout736 (.A(net738),
    .X(net736));
 sky130_fd_sc_hd__buf_1 fanout737 (.A(net738),
    .X(net737));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout738 (.A(net752),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_2 fanout739 (.A(net741),
    .X(net739));
 sky130_fd_sc_hd__buf_1 fanout740 (.A(net741),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_2 fanout741 (.A(net743),
    .X(net741));
 sky130_fd_sc_hd__buf_2 fanout742 (.A(net743),
    .X(net742));
 sky130_fd_sc_hd__clkbuf_2 fanout743 (.A(net752),
    .X(net743));
 sky130_fd_sc_hd__clkbuf_2 fanout744 (.A(net746),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_2 fanout745 (.A(net746),
    .X(net745));
 sky130_fd_sc_hd__buf_2 fanout746 (.A(net752),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_2 fanout747 (.A(net751),
    .X(net747));
 sky130_fd_sc_hd__buf_1 fanout748 (.A(net751),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_2 fanout749 (.A(net750),
    .X(net749));
 sky130_fd_sc_hd__buf_2 fanout750 (.A(net751),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_2 fanout751 (.A(net752),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_4 fanout752 (.A(net753),
    .X(net752));
 sky130_fd_sc_hd__buf_4 fanout753 (.A(\reg_module/rRs1[1] ),
    .X(net753));
 sky130_fd_sc_hd__clkbuf_2 fanout754 (.A(net764),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_2 fanout755 (.A(net756),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_2 fanout756 (.A(net764),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_2 fanout757 (.A(net761),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_2 fanout758 (.A(net761),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_2 fanout759 (.A(net760),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_2 fanout760 (.A(net761),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_2 fanout761 (.A(net763),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_2 fanout762 (.A(net763),
    .X(net762));
 sky130_fd_sc_hd__clkbuf_2 fanout763 (.A(net764),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_2 fanout764 (.A(net809),
    .X(net764));
 sky130_fd_sc_hd__clkbuf_2 fanout765 (.A(net767),
    .X(net765));
 sky130_fd_sc_hd__buf_1 fanout766 (.A(net767),
    .X(net766));
 sky130_fd_sc_hd__buf_2 fanout767 (.A(net774),
    .X(net767));
 sky130_fd_sc_hd__clkbuf_2 fanout768 (.A(net769),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_2 fanout769 (.A(net773),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_2 fanout770 (.A(net773),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_2 fanout771 (.A(net773),
    .X(net771));
 sky130_fd_sc_hd__buf_1 fanout772 (.A(net773),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_2 fanout773 (.A(net774),
    .X(net773));
 sky130_fd_sc_hd__buf_1 fanout774 (.A(net781),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_2 fanout775 (.A(net778),
    .X(net775));
 sky130_fd_sc_hd__buf_1 fanout776 (.A(net778),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_2 fanout777 (.A(net778),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_2 fanout778 (.A(net781),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_2 fanout779 (.A(net780),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_2 fanout780 (.A(net781),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_2 fanout781 (.A(net809),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_2 fanout782 (.A(net784),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_2 fanout783 (.A(net784),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_2 fanout784 (.A(net787),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_2 fanout785 (.A(net787),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_2 fanout786 (.A(net787),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_2 fanout787 (.A(net808),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_2 fanout788 (.A(net790),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_2 fanout789 (.A(net790),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_2 fanout790 (.A(net808),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_2 fanout791 (.A(net794),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_2 fanout792 (.A(net794),
    .X(net792));
 sky130_fd_sc_hd__buf_1 fanout793 (.A(net794),
    .X(net793));
 sky130_fd_sc_hd__clkbuf_2 fanout794 (.A(net807),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_2 fanout795 (.A(net796),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_2 fanout796 (.A(net799),
    .X(net796));
 sky130_fd_sc_hd__clkbuf_2 fanout797 (.A(net799),
    .X(net797));
 sky130_fd_sc_hd__clkbuf_2 fanout798 (.A(net799),
    .X(net798));
 sky130_fd_sc_hd__buf_1 fanout799 (.A(net807),
    .X(net799));
 sky130_fd_sc_hd__clkbuf_2 fanout800 (.A(net801),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_2 fanout801 (.A(net802),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_2 fanout802 (.A(net807),
    .X(net802));
 sky130_fd_sc_hd__clkbuf_2 fanout803 (.A(net804),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_2 fanout804 (.A(net806),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_2 fanout805 (.A(net806),
    .X(net805));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout806 (.A(net807),
    .X(net806));
 sky130_fd_sc_hd__buf_2 fanout807 (.A(net808),
    .X(net807));
 sky130_fd_sc_hd__buf_2 fanout808 (.A(net809),
    .X(net808));
 sky130_fd_sc_hd__buf_2 fanout809 (.A(\reg_module/rRs1[0] ),
    .X(net809));
 sky130_fd_sc_hd__clkbuf_2 fanout810 (.A(net811),
    .X(net810));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout811 (.A(net814),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_2 fanout812 (.A(net814),
    .X(net812));
 sky130_fd_sc_hd__buf_1 fanout813 (.A(net814),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_1 fanout814 (.A(net829),
    .X(net814));
 sky130_fd_sc_hd__clkbuf_2 fanout815 (.A(net819),
    .X(net815));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout816 (.A(net819),
    .X(net816));
 sky130_fd_sc_hd__clkbuf_2 fanout817 (.A(net819),
    .X(net817));
 sky130_fd_sc_hd__buf_1 fanout818 (.A(net819),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_2 fanout819 (.A(net829),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_2 fanout820 (.A(net821),
    .X(net820));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout821 (.A(net823),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_2 fanout822 (.A(net823),
    .X(net822));
 sky130_fd_sc_hd__buf_1 fanout823 (.A(net829),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_2 fanout824 (.A(net825),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_2 fanout825 (.A(net828),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_2 fanout826 (.A(net828),
    .X(net826));
 sky130_fd_sc_hd__buf_1 fanout827 (.A(net828),
    .X(net827));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout828 (.A(net829),
    .X(net828));
 sky130_fd_sc_hd__buf_2 fanout829 (.A(net881),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_2 fanout830 (.A(net831),
    .X(net830));
 sky130_fd_sc_hd__clkbuf_2 fanout831 (.A(net832),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_2 fanout832 (.A(net844),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_2 fanout833 (.A(net834),
    .X(net833));
 sky130_fd_sc_hd__buf_1 fanout834 (.A(net844),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_2 fanout835 (.A(net836),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_2 fanout836 (.A(net843),
    .X(net836));
 sky130_fd_sc_hd__buf_1 fanout837 (.A(net843),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_2 fanout838 (.A(net839),
    .X(net838));
 sky130_fd_sc_hd__buf_1 fanout839 (.A(net842),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_2 fanout840 (.A(net841),
    .X(net840));
 sky130_fd_sc_hd__clkbuf_2 fanout841 (.A(net842),
    .X(net841));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout842 (.A(net843),
    .X(net842));
 sky130_fd_sc_hd__buf_1 fanout843 (.A(net844),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_2 fanout844 (.A(net881),
    .X(net844));
 sky130_fd_sc_hd__clkbuf_2 fanout845 (.A(net846),
    .X(net845));
 sky130_fd_sc_hd__buf_2 fanout846 (.A(net851),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_2 fanout847 (.A(net850),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_2 fanout848 (.A(net850),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_2 fanout849 (.A(net850),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_2 fanout850 (.A(net851),
    .X(net850));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout851 (.A(net880),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_2 fanout852 (.A(net854),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_2 fanout853 (.A(net854),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_2 fanout854 (.A(net860),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_2 fanout855 (.A(net860),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_2 fanout856 (.A(net859),
    .X(net856));
 sky130_fd_sc_hd__buf_1 fanout857 (.A(net859),
    .X(net857));
 sky130_fd_sc_hd__clkbuf_2 fanout858 (.A(net859),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_2 fanout859 (.A(net860),
    .X(net859));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout860 (.A(net880),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_2 fanout861 (.A(net862),
    .X(net861));
 sky130_fd_sc_hd__buf_1 fanout862 (.A(net864),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_2 fanout863 (.A(net864),
    .X(net863));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout864 (.A(net879),
    .X(net864));
 sky130_fd_sc_hd__clkbuf_2 fanout865 (.A(net869),
    .X(net865));
 sky130_fd_sc_hd__buf_1 fanout866 (.A(net869),
    .X(net866));
 sky130_fd_sc_hd__clkbuf_2 fanout867 (.A(net868),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_2 fanout868 (.A(net869),
    .X(net868));
 sky130_fd_sc_hd__buf_1 fanout869 (.A(net879),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_2 fanout870 (.A(net873),
    .X(net870));
 sky130_fd_sc_hd__buf_1 fanout871 (.A(net873),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_2 fanout872 (.A(net873),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_2 fanout873 (.A(net879),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_2 fanout874 (.A(net878),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_2 fanout875 (.A(net878),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_2 fanout876 (.A(net877),
    .X(net876));
 sky130_fd_sc_hd__buf_1 fanout877 (.A(net878),
    .X(net877));
 sky130_fd_sc_hd__buf_1 fanout878 (.A(net879),
    .X(net878));
 sky130_fd_sc_hd__buf_2 fanout879 (.A(net880),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_2 fanout880 (.A(net881),
    .X(net880));
 sky130_fd_sc_hd__buf_2 fanout881 (.A(\reg_module/rRs1[0] ),
    .X(net881));
 sky130_fd_sc_hd__clkbuf_2 fanout882 (.A(net883),
    .X(net882));
 sky130_fd_sc_hd__clkbuf_2 fanout883 (.A(net887),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_2 fanout884 (.A(net886),
    .X(net884));
 sky130_fd_sc_hd__buf_1 fanout885 (.A(net886),
    .X(net885));
 sky130_fd_sc_hd__clkbuf_4 fanout886 (.A(net887),
    .X(net886));
 sky130_fd_sc_hd__clkbuf_2 fanout887 (.A(\dec/rStall1 ),
    .X(net887));
 sky130_fd_sc_hd__buf_2 fanout888 (.A(net891),
    .X(net888));
 sky130_fd_sc_hd__clkbuf_2 fanout889 (.A(net891),
    .X(net889));
 sky130_fd_sc_hd__buf_1 fanout890 (.A(net891),
    .X(net890));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout891 (.A(\dec/rStall2 ),
    .X(net891));
 sky130_fd_sc_hd__clkbuf_2 fanout892 (.A(net895),
    .X(net892));
 sky130_fd_sc_hd__clkbuf_2 fanout893 (.A(net895),
    .X(net893));
 sky130_fd_sc_hd__clkbuf_2 fanout894 (.A(net895),
    .X(net894));
 sky130_fd_sc_hd__buf_1 fanout895 (.A(\dec/rStall2 ),
    .X(net895));
 sky130_fd_sc_hd__buf_2 fanout896 (.A(net897),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_2 fanout897 (.A(b_type),
    .X(net897));
 sky130_fd_sc_hd__clkbuf_2 fanout898 (.A(net899),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_2 fanout899 (.A(op_jalr),
    .X(net899));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout900 (.A(net901),
    .X(net900));
 sky130_fd_sc_hd__clkbuf_2 fanout901 (.A(net906),
    .X(net901));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout902 (.A(net903),
    .X(net902));
 sky130_fd_sc_hd__buf_1 fanout903 (.A(net904),
    .X(net903));
 sky130_fd_sc_hd__buf_1 fanout904 (.A(net905),
    .X(net904));
 sky130_fd_sc_hd__buf_1 fanout905 (.A(net906),
    .X(net905));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout906 (.A(op_jalr),
    .X(net906));
 sky130_fd_sc_hd__clkbuf_2 fanout907 (.A(net914),
    .X(net907));
 sky130_fd_sc_hd__buf_1 fanout908 (.A(net914),
    .X(net908));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout909 (.A(net910),
    .X(net909));
 sky130_fd_sc_hd__clkbuf_2 fanout910 (.A(net914),
    .X(net910));
 sky130_fd_sc_hd__buf_1 fanout911 (.A(net912),
    .X(net911));
 sky130_fd_sc_hd__buf_1 fanout912 (.A(net913),
    .X(net912));
 sky130_fd_sc_hd__buf_1 fanout913 (.A(net914),
    .X(net913));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout914 (.A(net921),
    .X(net914));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout915 (.A(net917),
    .X(net915));
 sky130_fd_sc_hd__buf_1 fanout916 (.A(net920),
    .X(net916));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout917 (.A(net920),
    .X(net917));
 sky130_fd_sc_hd__buf_1 fanout918 (.A(net919),
    .X(net918));
 sky130_fd_sc_hd__clkbuf_2 fanout919 (.A(net920),
    .X(net919));
 sky130_fd_sc_hd__clkbuf_2 fanout920 (.A(net921),
    .X(net920));
 sky130_fd_sc_hd__buf_2 fanout921 (.A(op_auipc),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_2 fanout922 (.A(net924),
    .X(net922));
 sky130_fd_sc_hd__clkbuf_2 fanout923 (.A(net924),
    .X(net923));
 sky130_fd_sc_hd__clkbuf_2 fanout924 (.A(net928),
    .X(net924));
 sky130_fd_sc_hd__clkbuf_2 fanout925 (.A(net926),
    .X(net925));
 sky130_fd_sc_hd__clkbuf_2 fanout926 (.A(net927),
    .X(net926));
 sky130_fd_sc_hd__clkbuf_2 fanout927 (.A(net928),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_2 fanout928 (.A(op_lui),
    .X(net928));
 sky130_fd_sc_hd__clkbuf_2 fanout929 (.A(net931),
    .X(net929));
 sky130_fd_sc_hd__buf_1 fanout930 (.A(net931),
    .X(net930));
 sky130_fd_sc_hd__buf_1 fanout931 (.A(net938),
    .X(net931));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout932 (.A(net938),
    .X(net932));
 sky130_fd_sc_hd__clkbuf_2 fanout933 (.A(net937),
    .X(net933));
 sky130_fd_sc_hd__buf_1 fanout934 (.A(net937),
    .X(net934));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout935 (.A(net937),
    .X(net935));
 sky130_fd_sc_hd__buf_1 fanout936 (.A(net937),
    .X(net936));
 sky130_fd_sc_hd__buf_1 fanout937 (.A(net938),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_2 fanout938 (.A(\brancher/rAdder_b[13] ),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_2 fanout939 (.A(net941),
    .X(net939));
 sky130_fd_sc_hd__buf_1 fanout940 (.A(net941),
    .X(net940));
 sky130_fd_sc_hd__buf_2 fanout941 (.A(\brancher/rOp_jal ),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_2 fanout942 (.A(net943),
    .X(net942));
 sky130_fd_sc_hd__clkbuf_2 fanout943 (.A(net944),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_2 fanout944 (.A(\brancher/rOp_jal ),
    .X(net944));
 sky130_fd_sc_hd__clkbuf_2 fanout945 (.A(net947),
    .X(net945));
 sky130_fd_sc_hd__buf_1 fanout946 (.A(net947),
    .X(net946));
 sky130_fd_sc_hd__clkbuf_2 fanout947 (.A(\brancher/rOp_jalr ),
    .X(net947));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout948 (.A(net950),
    .X(net948));
 sky130_fd_sc_hd__buf_1 fanout949 (.A(net950),
    .X(net949));
 sky130_fd_sc_hd__buf_1 fanout950 (.A(net953),
    .X(net950));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout951 (.A(net953),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_2 fanout952 (.A(net953),
    .X(net952));
 sky130_fd_sc_hd__buf_1 fanout953 (.A(\brancher/rAdder_jal[21] ),
    .X(net953));
 sky130_fd_sc_hd__clkbuf_2 fanout954 (.A(\brancher/rPc_current_reg3[28] ),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_2 fanout955 (.A(\brancher/rPc_current_reg3[27] ),
    .X(net955));
 sky130_fd_sc_hd__clkbuf_2 fanout956 (.A(\brancher/rPc_current_reg3[26] ),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_2 fanout957 (.A(\brancher/rPc_current_reg3[25] ),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_2 fanout958 (.A(\brancher/rPc_current_reg3[21] ),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_2 fanout959 (.A(net961),
    .X(net959));
 sky130_fd_sc_hd__buf_1 fanout960 (.A(net961),
    .X(net960));
 sky130_fd_sc_hd__clkbuf_2 fanout961 (.A(net2072),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_4 fanout962 (.A(\rReg_d2[4] ),
    .X(net962));
 sky130_fd_sc_hd__buf_2 fanout963 (.A(net965),
    .X(net963));
 sky130_fd_sc_hd__buf_1 fanout964 (.A(net965),
    .X(net964));
 sky130_fd_sc_hd__buf_1 fanout965 (.A(net966),
    .X(net965));
 sky130_fd_sc_hd__buf_1 fanout966 (.A(net967),
    .X(net966));
 sky130_fd_sc_hd__clkbuf_4 fanout967 (.A(net970),
    .X(net967));
 sky130_fd_sc_hd__buf_2 fanout968 (.A(net970),
    .X(net968));
 sky130_fd_sc_hd__buf_1 fanout969 (.A(net970),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_4 fanout970 (.A(\rReg_d2[3] ),
    .X(net970));
 sky130_fd_sc_hd__buf_2 fanout971 (.A(net975),
    .X(net971));
 sky130_fd_sc_hd__buf_1 fanout972 (.A(net975),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_2 fanout973 (.A(net974),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_2 fanout974 (.A(net975),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_4 fanout975 (.A(\rReg_d2[3] ),
    .X(net975));
 sky130_fd_sc_hd__clkbuf_2 fanout976 (.A(net977),
    .X(net976));
 sky130_fd_sc_hd__buf_2 fanout977 (.A(net980),
    .X(net977));
 sky130_fd_sc_hd__buf_2 fanout978 (.A(net979),
    .X(net978));
 sky130_fd_sc_hd__clkbuf_2 fanout979 (.A(net980),
    .X(net979));
 sky130_fd_sc_hd__buf_2 fanout980 (.A(net993),
    .X(net980));
 sky130_fd_sc_hd__clkbuf_2 fanout981 (.A(net984),
    .X(net981));
 sky130_fd_sc_hd__clkbuf_2 fanout982 (.A(net984),
    .X(net982));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout983 (.A(net984),
    .X(net983));
 sky130_fd_sc_hd__buf_2 fanout984 (.A(net993),
    .X(net984));
 sky130_fd_sc_hd__clkbuf_2 fanout985 (.A(net987),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_1 fanout986 (.A(net987),
    .X(net986));
 sky130_fd_sc_hd__clkbuf_4 fanout987 (.A(net993),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_2 fanout988 (.A(net989),
    .X(net988));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout989 (.A(net990),
    .X(net989));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout990 (.A(net992),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_2 fanout991 (.A(net992),
    .X(net991));
 sky130_fd_sc_hd__clkbuf_2 fanout992 (.A(net993),
    .X(net992));
 sky130_fd_sc_hd__buf_4 fanout993 (.A(\rReg_d2[2] ),
    .X(net993));
 sky130_fd_sc_hd__clkbuf_4 fanout994 (.A(\rReg_d2[1] ),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_4 fanout995 (.A(\rReg_d2[0] ),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_2 fanout996 (.A(net998),
    .X(net996));
 sky130_fd_sc_hd__buf_1 fanout997 (.A(net998),
    .X(net997));
 sky130_fd_sc_hd__clkbuf_2 fanout998 (.A(rOp_memLd2),
    .X(net998));
 sky130_fd_sc_hd__buf_2 fanout999 (.A(net1003),
    .X(net999));
 sky130_fd_sc_hd__clkbuf_2 fanout1000 (.A(net1002),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_2 fanout1001 (.A(net1003),
    .X(net1001));
 sky130_fd_sc_hd__buf_1 fanout1002 (.A(net1003),
    .X(net1002));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1003 (.A(rOp_memLd2),
    .X(net1003));
 sky130_fd_sc_hd__clkbuf_2 fanout1004 (.A(net1008),
    .X(net1004));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1005 (.A(net1008),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_2 fanout1006 (.A(net1008),
    .X(net1006));
 sky130_fd_sc_hd__buf_1 fanout1007 (.A(net1008),
    .X(net1007));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1008 (.A(net1009),
    .X(net1008));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1009 (.A(net1031),
    .X(net1009));
 sky130_fd_sc_hd__clkbuf_2 fanout1010 (.A(net1011),
    .X(net1010));
 sky130_fd_sc_hd__clkbuf_2 fanout1011 (.A(net1013),
    .X(net1011));
 sky130_fd_sc_hd__buf_2 fanout1012 (.A(net1013),
    .X(net1012));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1013 (.A(net1014),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_4 fanout1014 (.A(net1031),
    .X(net1014));
 sky130_fd_sc_hd__clkbuf_2 fanout1015 (.A(net1016),
    .X(net1015));
 sky130_fd_sc_hd__clkbuf_2 fanout1016 (.A(net1022),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_2 fanout1017 (.A(net1018),
    .X(net1017));
 sky130_fd_sc_hd__buf_1 fanout1018 (.A(net1019),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_2 fanout1019 (.A(net1022),
    .X(net1019));
 sky130_fd_sc_hd__clkbuf_2 fanout1020 (.A(net1021),
    .X(net1020));
 sky130_fd_sc_hd__clkbuf_1 fanout1021 (.A(net1022),
    .X(net1021));
 sky130_fd_sc_hd__clkbuf_2 fanout1022 (.A(net1031),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_2 fanout1023 (.A(net1025),
    .X(net1023));
 sky130_fd_sc_hd__buf_1 fanout1024 (.A(net1025),
    .X(net1024));
 sky130_fd_sc_hd__clkbuf_2 fanout1025 (.A(net1026),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_4 fanout1026 (.A(net1030),
    .X(net1026));
 sky130_fd_sc_hd__clkbuf_2 fanout1027 (.A(net1028),
    .X(net1027));
 sky130_fd_sc_hd__buf_2 fanout1028 (.A(net1029),
    .X(net1028));
 sky130_fd_sc_hd__buf_2 fanout1029 (.A(net1030),
    .X(net1029));
 sky130_fd_sc_hd__clkbuf_2 fanout1030 (.A(net1031),
    .X(net1030));
 sky130_fd_sc_hd__buf_4 fanout1031 (.A(net1068),
    .X(net1031));
 sky130_fd_sc_hd__clkbuf_2 fanout1032 (.A(net1034),
    .X(net1032));
 sky130_fd_sc_hd__buf_1 fanout1033 (.A(net1034),
    .X(net1033));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1034 (.A(net1046),
    .X(net1034));
 sky130_fd_sc_hd__clkbuf_2 fanout1035 (.A(net1036),
    .X(net1035));
 sky130_fd_sc_hd__clkbuf_2 fanout1036 (.A(net1037),
    .X(net1036));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1037 (.A(net1046),
    .X(net1037));
 sky130_fd_sc_hd__clkbuf_2 fanout1038 (.A(net1041),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_2 fanout1039 (.A(net1041),
    .X(net1039));
 sky130_fd_sc_hd__clkbuf_2 fanout1040 (.A(net1041),
    .X(net1040));
 sky130_fd_sc_hd__clkbuf_2 fanout1041 (.A(net1046),
    .X(net1041));
 sky130_fd_sc_hd__clkbuf_2 fanout1042 (.A(net1045),
    .X(net1042));
 sky130_fd_sc_hd__buf_1 fanout1043 (.A(net1045),
    .X(net1043));
 sky130_fd_sc_hd__clkbuf_2 fanout1044 (.A(net1045),
    .X(net1044));
 sky130_fd_sc_hd__clkbuf_2 fanout1045 (.A(net1046),
    .X(net1045));
 sky130_fd_sc_hd__buf_2 fanout1046 (.A(net1057),
    .X(net1046));
 sky130_fd_sc_hd__buf_2 fanout1047 (.A(net1052),
    .X(net1047));
 sky130_fd_sc_hd__clkbuf_2 fanout1048 (.A(net1050),
    .X(net1048));
 sky130_fd_sc_hd__buf_1 fanout1049 (.A(net1050),
    .X(net1049));
 sky130_fd_sc_hd__buf_1 fanout1050 (.A(net1051),
    .X(net1050));
 sky130_fd_sc_hd__clkbuf_2 fanout1051 (.A(net1052),
    .X(net1051));
 sky130_fd_sc_hd__clkbuf_2 fanout1052 (.A(net1057),
    .X(net1052));
 sky130_fd_sc_hd__clkbuf_2 fanout1053 (.A(net1056),
    .X(net1053));
 sky130_fd_sc_hd__clkbuf_2 fanout1054 (.A(net1056),
    .X(net1054));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1055 (.A(net1056),
    .X(net1055));
 sky130_fd_sc_hd__clkbuf_2 fanout1056 (.A(net1057),
    .X(net1056));
 sky130_fd_sc_hd__buf_2 fanout1057 (.A(net1068),
    .X(net1057));
 sky130_fd_sc_hd__buf_2 fanout1058 (.A(net1062),
    .X(net1058));
 sky130_fd_sc_hd__clkbuf_2 fanout1059 (.A(net1060),
    .X(net1059));
 sky130_fd_sc_hd__buf_1 fanout1060 (.A(net1061),
    .X(net1060));
 sky130_fd_sc_hd__clkbuf_2 fanout1061 (.A(net1062),
    .X(net1061));
 sky130_fd_sc_hd__buf_1 fanout1062 (.A(net1067),
    .X(net1062));
 sky130_fd_sc_hd__clkbuf_2 fanout1063 (.A(net1064),
    .X(net1063));
 sky130_fd_sc_hd__buf_1 fanout1064 (.A(net1065),
    .X(net1064));
 sky130_fd_sc_hd__clkbuf_2 fanout1065 (.A(net1066),
    .X(net1065));
 sky130_fd_sc_hd__buf_2 fanout1066 (.A(net1067),
    .X(net1066));
 sky130_fd_sc_hd__buf_2 fanout1067 (.A(net1068),
    .X(net1067));
 sky130_fd_sc_hd__buf_4 fanout1068 (.A(net66),
    .X(net1068));
 sky130_fd_sc_hd__buf_1 fanout1069 (.A(net1071),
    .X(net1069));
 sky130_fd_sc_hd__buf_1 fanout1070 (.A(net1071),
    .X(net1070));
 sky130_fd_sc_hd__clkbuf_2 fanout1071 (.A(net1072),
    .X(net1071));
 sky130_fd_sc_hd__buf_1 fanout1072 (.A(net1073),
    .X(net1072));
 sky130_fd_sc_hd__buf_2 fanout1073 (.A(net1),
    .X(net1073));
 sky130_fd_sc_hd__conb_1 \brancher/_2171__1074  (.LO(net1074));
 sky130_fd_sc_hd__conb_1 _1877__1077 (.LO(net1077));
 sky130_fd_sc_hd__conb_1 _1885__1079 (.LO(net1079));
 sky130_fd_sc_hd__conb_1 _1892__1081 (.LO(net1081));
 sky130_fd_sc_hd__conb_1 _1897__1083 (.LO(net1083));
 sky130_fd_sc_hd__conb_1 _1902__1085 (.LO(net1085));
 sky130_fd_sc_hd__conb_1 _1906__1087 (.LO(net1087));
 sky130_fd_sc_hd__conb_1 _1911__1089 (.LO(net1089));
 sky130_fd_sc_hd__conb_1 _1917__1091 (.LO(net1091));
 sky130_fd_sc_hd__conb_1 _1922__1093 (.LO(net1093));
 sky130_fd_sc_hd__conb_1 _1926__1095 (.LO(net1095));
 sky130_fd_sc_hd__conb_1 _1931__1097 (.LO(net1097));
 sky130_fd_sc_hd__conb_1 _1935__1099 (.LO(net1099));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_44_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_45_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_46_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_47_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_48_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_49_clk (.A(clknet_4_5__leaf_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_50_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_51_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_52_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_53_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_54_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_55_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_56_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_57_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_58_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_59_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_60_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_61_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_62_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_63_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_64_clk (.A(clknet_4_4__leaf_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_65_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_66_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_67_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_68_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_69_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_70_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_71_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_72_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_73_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_74_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_75_clk (.A(clknet_4_3__leaf_clk),
    .X(clknet_leaf_75_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_76_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_77_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_77_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_78_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_78_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_79_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_79_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_80_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_81_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_82_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_83_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_83_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_84_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_85_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_85_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_86_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_86_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_87_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_87_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_88_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_88_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_89_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_89_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_90_clk (.A(clknet_4_6__leaf_clk),
    .X(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_91_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_91_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_92_clk (.A(clknet_4_7__leaf_clk),
    .X(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_95_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_95_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_96_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_97_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_98_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_98_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_99_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_99_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_100_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_101_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_101_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_102_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_103_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_103_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_104_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_105_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_106_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_107_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_108_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_108_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_109_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_110_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_111_clk (.A(clknet_4_15__leaf_clk),
    .X(clknet_leaf_111_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_112_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_112_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_113_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_114_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_115_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_115_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_116_clk (.A(clknet_4_13__leaf_clk),
    .X(clknet_leaf_116_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_117_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_118_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_119_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_120_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_121_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_122_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_122_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_123_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_123_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_124_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_125_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_126_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_127_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_128_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_129_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_130_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_130_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_131_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_132_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_133_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_134_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_134_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_135_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_135_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_136_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_136_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_137_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_138_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_139_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_140_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_141_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_141_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_142_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_143_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_143_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_144_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_144_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_145_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_146_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_147_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_148_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_149_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_150_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_150_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_151_clk (.A(clknet_4_14__leaf_clk),
    .X(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_152_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_153_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_154_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_155_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_156_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_156_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_157_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_157_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_158_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_158_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_159_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_159_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_160_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_161_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_162_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_162_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_163_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_163_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_164_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_165_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_165_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_166_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_167_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_167_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_168_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_169_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_169_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_170_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_171_clk (.A(clknet_4_10__leaf_clk),
    .X(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_172_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_173_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_174_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_175_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_175_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_176_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_176_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_177_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_178_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_178_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_179_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_179_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_180_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_181_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_182_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_183_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_184_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_185_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_185_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_186_clk (.A(clknet_4_11__leaf_clk),
    .X(clknet_leaf_186_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_187_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_188_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_189_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_189_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_190_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_191_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_192_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_193_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_193_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_194_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_195_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_196_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_197_clk (.A(clknet_4_12__leaf_clk),
    .X(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_198_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_198_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_199_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_200_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_201_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_202_clk (.A(clknet_4_9__leaf_clk),
    .X(clknet_leaf_202_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_203_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_204_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_205_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_206_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_206_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_207_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_207_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_208_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_209_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_209_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_210_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_210_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_211_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_212_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_213_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_214_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_214_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_215_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_215_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_216_clk (.A(clknet_4_8__leaf_clk),
    .X(clknet_leaf_216_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_217_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_217_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_218_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_218_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_219_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_219_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_220_clk (.A(clknet_4_0__leaf_clk),
    .X(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_221_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_222_clk (.A(clknet_4_2__leaf_clk),
    .X(clknet_leaf_222_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_223_clk (.A(clknet_4_1__leaf_clk),
    .X(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_clk (.A(clknet_0_clk),
    .X(clknet_2_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_clk (.A(clknet_0_clk),
    .X(clknet_2_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_clk (.A(clknet_0_clk),
    .X(clknet_2_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_clk (.A(clknet_0_clk),
    .X(clknet_2_3_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3__f_clk (.A(clknet_2_0_0_clk),
    .X(clknet_4_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7__f_clk (.A(clknet_2_1_0_clk),
    .X(clknet_4_7__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_8__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11__f_clk (.A(clknet_2_2_0_clk),
    .X(clknet_4_11__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_12__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15__f_clk (.A(clknet_2_3_0_clk),
    .X(clknet_4_15__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload0 (.A(clknet_4_0__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_4_1__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload2 (.A(clknet_4_2__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload3 (.A(clknet_4_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload4 (.A(clknet_4_5__leaf_clk));
 sky130_fd_sc_hd__inv_12 clkload5 (.A(clknet_4_7__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload6 (.A(clknet_4_9__leaf_clk));
 sky130_fd_sc_hd__inv_12 clkload7 (.A(clknet_4_10__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload8 (.A(clknet_4_11__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload9 (.A(clknet_4_13__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload10 (.A(clknet_4_14__leaf_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload11 (.A(clknet_4_15__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload12 (.A(clknet_leaf_204_clk));
 sky130_fd_sc_hd__clkinv_4 clkload13 (.A(clknet_leaf_205_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload14 (.A(clknet_leaf_206_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload15 (.A(clknet_leaf_207_clk));
 sky130_fd_sc_hd__inv_6 clkload16 (.A(clknet_leaf_208_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload17 (.A(clknet_leaf_213_clk));
 sky130_fd_sc_hd__clkinv_2 clkload18 (.A(clknet_leaf_219_clk));
 sky130_fd_sc_hd__inv_6 clkload19 (.A(clknet_leaf_220_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload20 (.A(clknet_leaf_0_clk));
 sky130_fd_sc_hd__clkinv_2 clkload21 (.A(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload22 (.A(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkinv_4 clkload23 (.A(clknet_leaf_199_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload24 (.A(clknet_leaf_203_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload25 (.A(clknet_leaf_221_clk));
 sky130_fd_sc_hd__clkinv_2 clkload26 (.A(clknet_leaf_223_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload27 (.A(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload28 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload29 (.A(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload30 (.A(clknet_leaf_9_clk));
 sky130_fd_sc_hd__bufinv_16 clkload31 (.A(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload32 (.A(clknet_leaf_15_clk));
 sky130_fd_sc_hd__bufinv_16 clkload33 (.A(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload34 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__inv_6 clkload35 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload36 (.A(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload37 (.A(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkinv_2 clkload38 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload39 (.A(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkinv_4 clkload40 (.A(clknet_leaf_71_clk));
 sky130_fd_sc_hd__inv_6 clkload41 (.A(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload42 (.A(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkinv_4 clkload43 (.A(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkinv_4 clkload44 (.A(clknet_leaf_75_clk));
 sky130_fd_sc_hd__inv_8 clkload45 (.A(clknet_leaf_19_clk));
 sky130_fd_sc_hd__inv_8 clkload46 (.A(clknet_leaf_20_clk));
 sky130_fd_sc_hd__inv_8 clkload47 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__inv_6 clkload48 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__inv_12 clkload49 (.A(clknet_leaf_23_clk));
 sky130_fd_sc_hd__inv_6 clkload50 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload51 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkinv_4 clkload52 (.A(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload53 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkinv_8 clkload54 (.A(clknet_leaf_43_clk));
 sky130_fd_sc_hd__inv_8 clkload55 (.A(clknet_leaf_44_clk));
 sky130_fd_sc_hd__inv_6 clkload56 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkinv_8 clkload57 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__inv_8 clkload58 (.A(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload59 (.A(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkinv_2 clkload60 (.A(clknet_leaf_26_clk));
 sky130_fd_sc_hd__bufinv_16 clkload61 (.A(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkinv_2 clkload62 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkinv_4 clkload63 (.A(clknet_leaf_33_clk));
 sky130_fd_sc_hd__bufinv_16 clkload64 (.A(clknet_leaf_34_clk));
 sky130_fd_sc_hd__inv_8 clkload65 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__inv_8 clkload66 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__inv_6 clkload67 (.A(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload68 (.A(clknet_leaf_38_clk));
 sky130_fd_sc_hd__inv_6 clkload69 (.A(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkinv_4 clkload70 (.A(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkinv_4 clkload71 (.A(clknet_leaf_41_clk));
 sky130_fd_sc_hd__inv_8 clkload72 (.A(clknet_leaf_47_clk));
 sky130_fd_sc_hd__inv_8 clkload73 (.A(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkinv_4 clkload74 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload75 (.A(clknet_leaf_60_clk));
 sky130_fd_sc_hd__inv_6 clkload76 (.A(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkinv_4 clkload77 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkinv_4 clkload78 (.A(clknet_leaf_67_clk));
 sky130_fd_sc_hd__inv_8 clkload79 (.A(clknet_leaf_68_clk));
 sky130_fd_sc_hd__inv_6 clkload80 (.A(clknet_leaf_69_clk));
 sky130_fd_sc_hd__inv_8 clkload81 (.A(clknet_leaf_76_clk));
 sky130_fd_sc_hd__clkinv_8 clkload82 (.A(clknet_leaf_77_clk));
 sky130_fd_sc_hd__inv_6 clkload83 (.A(clknet_leaf_78_clk));
 sky130_fd_sc_hd__inv_8 clkload84 (.A(clknet_leaf_79_clk));
 sky130_fd_sc_hd__inv_8 clkload85 (.A(clknet_leaf_80_clk));
 sky130_fd_sc_hd__clkinv_8 clkload86 (.A(clknet_leaf_85_clk));
 sky130_fd_sc_hd__inv_6 clkload87 (.A(clknet_leaf_86_clk));
 sky130_fd_sc_hd__inv_6 clkload88 (.A(clknet_leaf_87_clk));
 sky130_fd_sc_hd__inv_8 clkload89 (.A(clknet_leaf_88_clk));
 sky130_fd_sc_hd__inv_12 clkload90 (.A(clknet_leaf_89_clk));
 sky130_fd_sc_hd__inv_8 clkload91 (.A(clknet_leaf_90_clk));
 sky130_fd_sc_hd__clkinv_8 clkload92 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__inv_12 clkload93 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__bufinv_16 clkload94 (.A(clknet_leaf_52_clk));
 sky130_fd_sc_hd__inv_8 clkload95 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__inv_12 clkload96 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload97 (.A(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload98 (.A(clknet_leaf_57_clk));
 sky130_fd_sc_hd__inv_6 clkload99 (.A(clknet_leaf_58_clk));
 sky130_fd_sc_hd__inv_12 clkload100 (.A(clknet_leaf_91_clk));
 sky130_fd_sc_hd__inv_12 clkload101 (.A(clknet_leaf_92_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload102 (.A(clknet_leaf_172_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload103 (.A(clknet_leaf_173_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload104 (.A(clknet_leaf_174_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload105 (.A(clknet_leaf_176_clk));
 sky130_fd_sc_hd__bufinv_16 clkload106 (.A(clknet_leaf_177_clk));
 sky130_fd_sc_hd__clkinv_4 clkload107 (.A(clknet_leaf_178_clk));
 sky130_fd_sc_hd__bufinv_16 clkload108 (.A(clknet_leaf_179_clk));
 sky130_fd_sc_hd__bufinv_16 clkload109 (.A(clknet_leaf_180_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload110 (.A(clknet_leaf_181_clk));
 sky130_fd_sc_hd__clkinv_2 clkload111 (.A(clknet_leaf_182_clk));
 sky130_fd_sc_hd__clkinv_4 clkload112 (.A(clknet_leaf_183_clk));
 sky130_fd_sc_hd__clkinv_2 clkload113 (.A(clknet_leaf_210_clk));
 sky130_fd_sc_hd__inv_6 clkload114 (.A(clknet_leaf_211_clk));
 sky130_fd_sc_hd__clkinv_4 clkload115 (.A(clknet_leaf_212_clk));
 sky130_fd_sc_hd__clkinv_4 clkload116 (.A(clknet_leaf_214_clk));
 sky130_fd_sc_hd__bufinv_16 clkload117 (.A(clknet_leaf_215_clk));
 sky130_fd_sc_hd__bufinv_16 clkload118 (.A(clknet_leaf_216_clk));
 sky130_fd_sc_hd__bufinv_16 clkload119 (.A(clknet_leaf_125_clk));
 sky130_fd_sc_hd__clkinv_4 clkload120 (.A(clknet_leaf_131_clk));
 sky130_fd_sc_hd__clkinv_4 clkload121 (.A(clknet_leaf_132_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload122 (.A(clknet_leaf_184_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload123 (.A(clknet_leaf_187_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload124 (.A(clknet_leaf_188_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload125 (.A(clknet_leaf_189_clk));
 sky130_fd_sc_hd__bufinv_16 clkload126 (.A(clknet_leaf_190_clk));
 sky130_fd_sc_hd__clkinv_4 clkload127 (.A(clknet_leaf_191_clk));
 sky130_fd_sc_hd__clkinv_4 clkload128 (.A(clknet_leaf_192_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload129 (.A(clknet_leaf_194_clk));
 sky130_fd_sc_hd__clkinv_4 clkload130 (.A(clknet_leaf_198_clk));
 sky130_fd_sc_hd__bufinv_16 clkload131 (.A(clknet_leaf_200_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload132 (.A(clknet_leaf_201_clk));
 sky130_fd_sc_hd__clkinv_2 clkload133 (.A(clknet_leaf_202_clk));
 sky130_fd_sc_hd__inv_6 clkload134 (.A(clknet_leaf_159_clk));
 sky130_fd_sc_hd__inv_6 clkload135 (.A(clknet_leaf_160_clk));
 sky130_fd_sc_hd__clkinv_2 clkload136 (.A(clknet_leaf_161_clk));
 sky130_fd_sc_hd__clkinv_4 clkload137 (.A(clknet_leaf_162_clk));
 sky130_fd_sc_hd__bufinv_16 clkload138 (.A(clknet_leaf_163_clk));
 sky130_fd_sc_hd__inv_6 clkload139 (.A(clknet_leaf_164_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload140 (.A(clknet_leaf_167_clk));
 sky130_fd_sc_hd__bufinv_16 clkload141 (.A(clknet_leaf_168_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload142 (.A(clknet_leaf_170_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload143 (.A(clknet_leaf_171_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload144 (.A(clknet_leaf_133_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload145 (.A(clknet_leaf_134_clk));
 sky130_fd_sc_hd__inv_8 clkload146 (.A(clknet_leaf_149_clk));
 sky130_fd_sc_hd__clkinv_4 clkload147 (.A(clknet_leaf_152_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload148 (.A(clknet_leaf_153_clk));
 sky130_fd_sc_hd__clkinv_2 clkload149 (.A(clknet_leaf_154_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload150 (.A(clknet_leaf_155_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload151 (.A(clknet_leaf_156_clk));
 sky130_fd_sc_hd__bufinv_16 clkload152 (.A(clknet_leaf_157_clk));
 sky130_fd_sc_hd__inv_8 clkload153 (.A(clknet_leaf_158_clk));
 sky130_fd_sc_hd__inv_8 clkload154 (.A(clknet_leaf_165_clk));
 sky130_fd_sc_hd__inv_6 clkload155 (.A(clknet_leaf_166_clk));
 sky130_fd_sc_hd__clkinv_4 clkload156 (.A(clknet_leaf_185_clk));
 sky130_fd_sc_hd__bufinv_16 clkload157 (.A(clknet_leaf_186_clk));
 sky130_fd_sc_hd__bufinv_16 clkload158 (.A(clknet_leaf_117_clk));
 sky130_fd_sc_hd__clkinv_4 clkload159 (.A(clknet_leaf_118_clk));
 sky130_fd_sc_hd__clkinv_2 clkload160 (.A(clknet_leaf_119_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload161 (.A(clknet_leaf_120_clk));
 sky130_fd_sc_hd__clkinv_4 clkload162 (.A(clknet_leaf_121_clk));
 sky130_fd_sc_hd__clkinv_2 clkload163 (.A(clknet_leaf_122_clk));
 sky130_fd_sc_hd__bufinv_16 clkload164 (.A(clknet_leaf_124_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload165 (.A(clknet_leaf_126_clk));
 sky130_fd_sc_hd__clkinv_2 clkload166 (.A(clknet_leaf_127_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload167 (.A(clknet_leaf_128_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload168 (.A(clknet_leaf_129_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload169 (.A(clknet_leaf_130_clk));
 sky130_fd_sc_hd__bufinv_16 clkload170 (.A(clknet_leaf_195_clk));
 sky130_fd_sc_hd__clkinv_4 clkload171 (.A(clknet_leaf_196_clk));
 sky130_fd_sc_hd__clkinv_4 clkload172 (.A(clknet_leaf_197_clk));
 sky130_fd_sc_hd__clkinv_4 clkload173 (.A(clknet_leaf_81_clk));
 sky130_fd_sc_hd__clkinv_4 clkload174 (.A(clknet_leaf_82_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload175 (.A(clknet_leaf_83_clk));
 sky130_fd_sc_hd__bufinv_16 clkload176 (.A(clknet_leaf_84_clk));
 sky130_fd_sc_hd__clkinv_4 clkload177 (.A(clknet_leaf_110_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload178 (.A(clknet_leaf_112_clk));
 sky130_fd_sc_hd__inv_6 clkload179 (.A(clknet_leaf_113_clk));
 sky130_fd_sc_hd__clkinv_2 clkload180 (.A(clknet_leaf_114_clk));
 sky130_fd_sc_hd__clkinv_2 clkload181 (.A(clknet_leaf_115_clk));
 sky130_fd_sc_hd__bufinv_16 clkload182 (.A(clknet_leaf_116_clk));
 sky130_fd_sc_hd__bufinv_16 clkload183 (.A(clknet_leaf_135_clk));
 sky130_fd_sc_hd__inv_6 clkload184 (.A(clknet_leaf_137_clk));
 sky130_fd_sc_hd__clkinv_4 clkload185 (.A(clknet_leaf_138_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload186 (.A(clknet_leaf_139_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload187 (.A(clknet_leaf_140_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload188 (.A(clknet_leaf_141_clk));
 sky130_fd_sc_hd__inv_6 clkload189 (.A(clknet_leaf_142_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload190 (.A(clknet_leaf_143_clk));
 sky130_fd_sc_hd__bufinv_16 clkload191 (.A(clknet_leaf_144_clk));
 sky130_fd_sc_hd__bufinv_16 clkload192 (.A(clknet_leaf_145_clk));
 sky130_fd_sc_hd__clkinv_4 clkload193 (.A(clknet_leaf_146_clk));
 sky130_fd_sc_hd__clkinv_2 clkload194 (.A(clknet_leaf_147_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload195 (.A(clknet_leaf_148_clk));
 sky130_fd_sc_hd__clkinv_4 clkload196 (.A(clknet_leaf_151_clk));
 sky130_fd_sc_hd__clkinv_4 clkload197 (.A(clknet_leaf_96_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload198 (.A(clknet_leaf_97_clk));
 sky130_fd_sc_hd__clkinv_4 clkload199 (.A(clknet_leaf_99_clk));
 sky130_fd_sc_hd__inv_6 clkload200 (.A(clknet_leaf_100_clk));
 sky130_fd_sc_hd__clkinv_4 clkload201 (.A(clknet_leaf_101_clk));
 sky130_fd_sc_hd__inv_8 clkload202 (.A(clknet_leaf_102_clk));
 sky130_fd_sc_hd__clkinv_4 clkload203 (.A(clknet_leaf_103_clk));
 sky130_fd_sc_hd__inv_6 clkload204 (.A(clknet_leaf_104_clk));
 sky130_fd_sc_hd__clkinv_4 clkload205 (.A(clknet_leaf_105_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload206 (.A(clknet_leaf_106_clk));
 sky130_fd_sc_hd__clkinv_4 clkload207 (.A(clknet_leaf_107_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload208 (.A(clknet_leaf_108_clk));
 sky130_fd_sc_hd__inv_6 clkload209 (.A(clknet_leaf_109_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload210 (.A(clknet_leaf_111_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\rWrData[1] ),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\dec/rInstrustion1[16] ),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\dec/rInstrustion1[19] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\dec/rInstrustion1[14] ),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\dec/rInstrustion1[5] ),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\dec/rInstrustion1[23] ),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\dec/rInstrustion1[8] ),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\dec/rInstrustion1[0] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\dec/rInstrustion1[22] ),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\dec/rInstrustion1[28] ),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\dec/rInstrustion1[11] ),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\dec/rInstrustion1[21] ),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\dec/rInstrustion1[3] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\dec/rInstrustion1[29] ),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(rOp_memLd),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\dec/rInstrustion1[1] ),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\dec/rInstrustion1[2] ),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\dec/rInstrustion1[9] ),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\dec/rInstrustion1[18] ),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\dec/rInstrustion1[20] ),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\dec/rInstrustion1[31] ),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\dec/rInstrustion1[24] ),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\dec/rInstrustion1[26] ),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\dec/rInstrustion1[17] ),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\dec/rInstrustion1[6] ),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\dec/rInstrustion1[10] ),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\dec/rInstrustion1[13] ),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\dec/rInstrustion1[30] ),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\dec/rInstrustion1[4] ),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\dec/rInstrustion1[27] ),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\dec/rInstrustion1[7] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\dec/rInstrustion1[15] ),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\dec/rInstrustion1[25] ),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\rWrData[27] ),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\imm21_j[15] ),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\imm13_b[11] ),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\rWrData[18] ),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\rWrData[16] ),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\imm21_j[11] ),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\imm13_b[4] ),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\rWrData[30] ),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\imm21_j[18] ),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\rWrData[31] ),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\dec/rInstrustion1[12] ),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\imm13_b[2] ),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\rWrData[29] ),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\rWrData[24] ),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\imm13_b[3] ),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\imm21_j[19] ),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\imm21_j[17] ),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\rWrData[14] ),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\imm13_b[1] ),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\imm21_j[2] ),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\imm21_j[16] ),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\rWrData[23] ),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\rWrData[2] ),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\rWrData[19] ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\imm21_j[14] ),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\rWrData[3] ),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\rWrData[25] ),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(i_type),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\rWrData[0] ),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\imm21_j[3] ),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\rWrData[10] ),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\rWrData[8] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\rReg_d[3] ),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\rWrData[13] ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\rReg_d[4] ),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(op_ecb),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\rWrData[4] ),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(u_type),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\imm21_j[4] ),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\Op_code[6] ),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\Op_code[5] ),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\Op_code[4] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\rWrData[5] ),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\rWrData[28] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\rWrData[22] ),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(op_efence),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\rWrData[11] ),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\Op_code[1] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\rWrData[21] ),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\Op_code[3] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\Op_code[0] ),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\Op_code[2] ),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(rRegWrEn),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\rWrData[26] ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\rWrData[12] ),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\rWrData[20] ),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\imm21_j[13] ),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\rWrData[17] ),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\imm21_j[12] ),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\rWrData[6] ),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\reg_module/gprf[993] ),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\reg_module/gprf[1016] ),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\reg_module/gprf[1014] ),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\reg_module/gprf[1018] ),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\reg_module/gprf[1017] ),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\reg_module/gprf[1012] ),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\reg_module/gprf[1020] ),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\reg_module/gprf[1004] ),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(op_memLd),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\reg_module/gprf[998] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(j_type),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\reg_module/gprf[1015] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\reg_module/gprf[1013] ),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\reg_module/gprf[1021] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\reg_module/gprf[1003] ),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\reg_module/gprf[1006] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\reg_module/gprf[1010] ),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\reg_module/gprf[996] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\reg_module/gprf[1008] ),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\reg_module/gprf[1011] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\reg_module/gprf[1000] ),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\rWrData[9] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\reg_module/gprf[999] ),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\reg_module/gprf[1019] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\reg_module/gprf[1001] ),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\reg_module/gprf[997] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\reg_module/gprf[994] ),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\reg_module/gprf[1005] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\reg_module/gprf[1002] ),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\reg_module/gprf[1023] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\reg_module/gprf[1022] ),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\reg_module/gprf[1007] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\rWrData[15] ),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\reg_module/gprf[995] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\reg_module/gprf[353] ),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\reg_module/gprf[979] ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\reg_module/gprf[429] ),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\reg_module/gprf[382] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\reg_module/gprf[442] ),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\reg_module/gprf[633] ),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\reg_module/gprf[694] ),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\reg_module/gprf[291] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\reg_module/gprf[672] ),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\reg_module/gprf[443] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\reg_module/gprf[745] ),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\reg_module/gprf[379] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\reg_module/gprf[305] ),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\reg_module/gprf[615] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\reg_module/gprf[503] ),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\reg_module/gprf[695] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\reg_module/gprf[504] ),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\reg_module/gprf[747] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\reg_module/gprf[426] ),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\reg_module/gprf[708] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\reg_module/gprf[124] ),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\reg_module/gprf[673] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\reg_module/gprf[444] ),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\reg_module/gprf[447] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\reg_module/gprf[617] ),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\reg_module/gprf[449] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\reg_module/gprf[693] ),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\reg_module/gprf[472] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\reg_module/gprf[985] ),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\reg_module/gprf[612] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\reg_module/gprf[188] ),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\reg_module/gprf[689] ),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\reg_module/gprf[377] ),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\reg_module/gprf[296] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\reg_module/gprf[482] ),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\reg_module/gprf[381] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\reg_module/gprf[624] ),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\reg_module/gprf[796] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\reg_module/gprf[280] ),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\reg_module/gprf[88] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\reg_module/gprf[33] ),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\reg_module/gprf[686] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\reg_module/gprf[1009] ),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\reg_module/gprf[753] ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\reg_module/gprf[575] ),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\reg_module/gprf[505] ),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\reg_module/gprf[510] ),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\reg_module/gprf[511] ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\reg_module/gprf[314] ),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\reg_module/gprf[981] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\reg_module/gprf[317] ),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\reg_module/gprf[297] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\reg_module/gprf[431] ),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\reg_module/gprf[691] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\reg_module/gprf[761] ),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\reg_module/gprf[621] ),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\reg_module/gprf[308] ),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\reg_module/gprf[574] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\reg_module/gprf[430] ),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\reg_module/gprf[759] ),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\reg_module/gprf[698] ),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\reg_module/gprf[43] ),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\reg_module/gprf[697] ),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\reg_module/gprf[425] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\reg_module/gprf[618] ),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\reg_module/gprf[298] ),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\reg_module/gprf[638] ),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\reg_module/gprf[692] ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\reg_module/gprf[334] ),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\reg_module/gprf[197] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\reg_module/gprf[187] ),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\reg_module/gprf[676] ),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\reg_module/gprf[632] ),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\reg_module/gprf[795] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\reg_module/gprf[725] ),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\reg_module/gprf[127] ),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\reg_module/gprf[115] ),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\reg_module/gprf[636] ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\reg_module/gprf[770] ),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\reg_module/gprf[212] ),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\reg_module/gprf[345] ),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\reg_module/gprf[730] ),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\reg_module/gprf[569] ),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\reg_module/gprf[185] ),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\reg_module/gprf[739] ),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\reg_module/gprf[111] ),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\reg_module/gprf[78] ),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\reg_module/gprf[375] ),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\reg_module/gprf[73] ),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\reg_module/gprf[755] ),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\reg_module/gprf[988] ),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\reg_module/gprf[34] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\reg_module/gprf[378] ),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\reg_module/gprf[545] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\reg_module/gprf[338] ),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\reg_module/gprf[507] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\reg_module/gprf[162] ),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\reg_module/gprf[278] ),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\reg_module/gprf[502] ),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\reg_module/gprf[493] ),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\reg_module/gprf[309] ),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\reg_module/gprf[380] ),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\reg_module/gprf[348] ),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\reg_module/gprf[623] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(net160),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\reg_module/gprf[161] ),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\reg_module/gprf[365] ),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\reg_module/gprf[751] ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\reg_module/gprf[726] ),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\reg_module/gprf[984] ),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\reg_module/gprf[295] ),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\reg_module/gprf[677] ),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\reg_module/gprf[468] ),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\reg_module/gprf[784] ),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\reg_module/gprf[64] ),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\reg_module/gprf[798] ),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\reg_module/gprf[41] ),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\reg_module/gprf[72] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\reg_module/gprf[428] ),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\reg_module/gprf[799] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\reg_module/gprf[776] ),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\reg_module/gprf[474] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\reg_module/gprf[789] ),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\reg_module/gprf[321] ),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\reg_module/gprf[366] ),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\reg_module/gprf[77] ),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\reg_module/gprf[344] ),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\reg_module/gprf[793] ),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\reg_module/gprf[42] ),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\reg_module/gprf[331] ),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\reg_module/gprf[93] ),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\reg_module/gprf[550] ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\reg_module/gprf[432] ),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\reg_module/gprf[961] ),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\reg_module/gprf[611] ),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\reg_module/gprf[108] ),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\reg_module/gprf[433] ),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\reg_module/gprf[763] ),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\reg_module/gprf[374] ),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\reg_module/gprf[794] ),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\reg_module/gprf[310] ),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\reg_module/gprf[221] ),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\reg_module/gprf[706] ),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\reg_module/gprf[40] ),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\reg_module/gprf[96] ),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\reg_module/gprf[470] ),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\reg_module/gprf[217] ),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\reg_module/gprf[471] ),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\reg_module/gprf[106] ),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\reg_module/gprf[635] ),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\reg_module/gprf[323] ),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\reg_module/gprf[289] ),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\reg_module/gprf[741] ),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\reg_module/gprf[304] ),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\reg_module/gprf[707] ),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\reg_module/gprf[714] ),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\reg_module/gprf[95] ),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\reg_module/gprf[990] ),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\reg_module/gprf[222] ),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\reg_module/gprf[987] ),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\reg_module/gprf[271] ),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\reg_module/gprf[639] ),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\reg_module/gprf[727] ),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\reg_module/gprf[288] ),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\reg_module/gprf[351] ),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\reg_module/gprf[35] ),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\reg_module/gprf[889] ),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\reg_module/gprf[473] ),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\reg_module/gprf[704] ),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\reg_module/gprf[416] ),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\reg_module/gprf[58] ),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\reg_module/gprf[456] ),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\reg_module/gprf[343] ),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\reg_module/gprf[220] ),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\imm21_j[1] ),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\reg_module/gprf[479] ),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\reg_module/gprf[746] ),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\reg_module/gprf[480] ),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\reg_module/gprf[113] ),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\reg_module/gprf[329] ),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\reg_module/gprf[508] ),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\reg_module/gprf[438] ),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\reg_module/gprf[448] ),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\reg_module/gprf[356] ),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\reg_module/gprf[437] ),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\reg_module/gprf[186] ),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\reg_module/gprf[705] ),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\reg_module/gprf[126] ),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\reg_module/gprf[978] ),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\reg_module/gprf[485] ),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\reg_module/gprf[461] ),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\reg_module/gprf[737] ),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\reg_module/gprf[783] ),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\reg_module/gprf[171] ),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\reg_module/gprf[109] ),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\reg_module/gprf[196] ),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\reg_module/gprf[980] ),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\reg_module/gprf[328] ),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\reg_module/gprf[120] ),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\reg_module/gprf[76] ),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\reg_module/gprf[613] ),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\reg_module/gprf[484] ),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\reg_module/gprf[300] ),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\reg_module/gprf[340] ),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\reg_module/gprf[481] ),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\reg_module/gprf[724] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\reg_module/gprf[100] ),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\reg_module/gprf[71] ),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\reg_module/gprf[110] ),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\reg_module/gprf[184] ),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\reg_module/gprf[506] ),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\reg_module/gprf[982] ),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\reg_module/gprf[84] ),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\reg_module/gprf[551] ),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\reg_module/gprf[614] ),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\reg_module/gprf[208] ),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\reg_module/gprf[568] ),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\reg_module/gprf[347] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\reg_module/gprf[591] ),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\reg_module/gprf[594] ),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\reg_module/gprf[359] ),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\reg_module/gprf[777] ),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\reg_module/gprf[89] ),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\reg_module/gprf[320] ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\reg_module/gprf[454] ),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\reg_module/gprf[209] ),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\reg_module/gprf[723] ),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\reg_module/gprf[620] ),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\reg_module/gprf[496] ),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\reg_module/gprf[101] ),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\reg_module/gprf[970] ),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\reg_module/gprf[977] ),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\reg_module/gprf[59] ),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\reg_module/gprf[711] ),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\reg_module/gprf[722] ),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\reg_module/gprf[976] ),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\reg_module/gprf[68] ),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\reg_module/gprf[261] ),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\reg_module/gprf[337] ),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\reg_module/gprf[589] ),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\reg_module/gprf[299] ),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\reg_module/gprf[446] ),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\reg_module/gprf[703] ),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\reg_module/gprf[103] ),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\reg_module/gprf[260] ),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\reg_module/gprf[341] ),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\reg_module/gprf[330] ),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\reg_module/gprf[690] ),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\reg_module/gprf[206] ),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\reg_module/gprf[774] ),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\reg_module/gprf[991] ),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\reg_module/gprf[696] ),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\reg_module/gprf[459] ),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\reg_module/gprf[455] ),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\reg_module/gprf[322] ),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\reg_module/gprf[893] ),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\reg_module/gprf[39] ),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\reg_module/gprf[674] ),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\reg_module/gprf[595] ),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\reg_module/gprf[70] ),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\reg_module/gprf[189] ),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\reg_module/gprf[460] ),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\reg_module/gprf[223] ),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\reg_module/gprf[782] ),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\reg_module/gprf[335] ),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\reg_module/gprf[207] ),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\reg_module/gprf[500] ),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\reg_module/gprf[262] ),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\reg_module/gprf[436] ),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\reg_module/gprf[316] ),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\reg_module/gprf[790] ),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\reg_module/gprf[272] ),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\reg_module/gprf[738] ),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\reg_module/gprf[303] ),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\reg_module/gprf[333] ),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\reg_module/gprf[797] ),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\reg_module/gprf[218] ),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\reg_module/gprf[79] ),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\reg_module/gprf[765] ),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\reg_module/gprf[350] ),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\reg_module/gprf[287] ),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(rHazardStallRs1),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(_0632_),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\reg_module/gprf[285] ),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\reg_module/gprf[609] ),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\reg_module/gprf[92] ),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\reg_module/gprf[509] ),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\reg_module/gprf[358] ),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\reg_module/gprf[792] ),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\reg_module/gprf[572] ),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\reg_module/gprf[423] ),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\reg_module/gprf[342] ),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\reg_module/gprf[688] ),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\reg_module/gprf[501] ),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\reg_module/gprf[57] ),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\reg_module/gprf[489] ),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\reg_module/gprf[865] ),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\reg_module/gprf[346] ),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\reg_module/gprf[975] ),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\reg_module/gprf[324] ),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\reg_module/gprf[326] ),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\reg_module/gprf[181] ),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\reg_module/gprf[292] ),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\reg_module/gprf[830] ),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\reg_module/gprf[894] ),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\reg_module/gprf[364] ),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\reg_module/gprf[105] ),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\reg_module/gprf[268] ),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\reg_module/gprf[785] ),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\reg_module/gprf[114] ),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\reg_module/gprf[373] ),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\reg_module/gprf[710] ),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\reg_module/gprf[119] ),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\reg_module/gprf[458] ),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\reg_module/gprf[182] ),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\reg_module/gprf[966] ),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\reg_module/gprf[166] ),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\reg_module/gprf[478] ),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\reg_module/gprf[466] ),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\reg_module/gprf[102] ),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\reg_module/gprf[891] ),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\reg_module/gprf[453] ),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\reg_module/gprf[332] ),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\reg_module/gprf[270] ),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\reg_module/gprf[339] ),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\reg_module/gprf[325] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\reg_module/gprf[198] ),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\reg_module/gprf[637] ),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\reg_module/gprf[315] ),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\reg_module/gprf[216] ),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(op_intRegImm),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\reg_module/gprf[720] ),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\reg_module/gprf[769] ),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\reg_module/gprf[90] ),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\reg_module/gprf[701] ),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\reg_module/gprf[974] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\reg_module/gprf[192] ),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\reg_module/gprf[439] ),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\reg_module/gprf[36] ),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\reg_module/gprf[441] ),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\reg_module/gprf[742] ),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\reg_module/gprf[492] ),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\reg_module/gprf[49] ),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\reg_module/gprf[548] ),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\reg_module/gprf[892] ),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\reg_module/gprf[69] ),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\reg_module/gprf[211] ),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\reg_module/gprf[554] ),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\reg_module/gprf[74] ),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\reg_module/gprf[972] ),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\reg_module/gprf[200] ),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\reg_module/gprf[258] ),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\reg_module/gprf[678] ),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\reg_module/gprf[743] ),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\reg_module/gprf[125] ),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\reg_module/gprf[679] ),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\reg_module/gprf[773] ),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\reg_module/gprf[83] ),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\reg_module/gprf[702] ),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\reg_module/gprf[464] ),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\reg_module/gprf[716] ),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\reg_module/gprf[445] ),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\reg_module/gprf[549] ),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\reg_module/gprf[190] ),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\reg_module/gprf[962] ),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\reg_module/gprf[191] ),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\reg_module/gprf[465] ),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\reg_module/gprf[592] ),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\reg_module/gprf[631] ),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\reg_module/gprf[75] ),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\reg_module/gprf[486] ),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\reg_module/gprf[372] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\reg_module/gprf[475] ),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\reg_module/gprf[179] ),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\reg_module/gprf[194] ),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\reg_module/gprf[38] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\reg_module/gprf[967] ),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\reg_module/gprf[327] ),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\reg_module/gprf[176] ),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\reg_module/gprf[37] ),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\reg_module/gprf[264] ),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\reg_module/gprf[973] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\reg_module/gprf[169] ),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\reg_module/gprf[193] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\reg_module/gprf[281] ),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\reg_module/gprf[293] ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\reg_module/gprf[420] ),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\reg_module/gprf[579] ),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\reg_module/gprf[457] ),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\reg_module/gprf[583] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\reg_module/gprf[48] ),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\reg_module/gprf[597] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\reg_module/gprf[888] ),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\reg_module/gprf[376] ),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\reg_module/gprf[294] ),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\reg_module/gprf[749] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\reg_module/gprf[214] ),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\reg_module/gprf[864] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\reg_module/gprf[121] ),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\reg_module/gprf[85] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\reg_module/gprf[969] ),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\reg_module/gprf[992] ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\reg_module/gprf[628] ),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\reg_module/gprf[964] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\reg_module/gprf[91] ),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\reg_module/gprf[649] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\reg_module/gprf[66] ),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\reg_module/gprf[733] ),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\reg_module/gprf[488] ),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\reg_module/gprf[573] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\reg_module/gprf[203] ),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\reg_module/gprf[634] ),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\reg_module/gprf[607] ),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\reg_module/gprf[483] ),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\reg_module/gprf[118] ),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\reg_module/gprf[546] ),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\reg_module/gprf[469] ),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\reg_module/gprf[947] ),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\reg_module/gprf[273] ),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\reg_module/gprf[107] ),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(\reg_module/gprf[670] ),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\reg_module/gprf[766] ),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\reg_module/gprf[452] ),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\reg_module/gprf[213] ),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\reg_module/gprf[112] ),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\reg_module/gprf[576] ),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\reg_module/gprf[63] ),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\reg_module/gprf[487] ),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\reg_module/gprf[578] ),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\reg_module/gprf[180] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\reg_module/gprf[422] ),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\reg_module/gprf[417] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\reg_module/gprf[177] ),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\reg_module/gprf[752] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\reg_module/gprf[362] ),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\reg_module/gprf[930] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\reg_module/gprf[491] ),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\reg_module/gprf[463] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\reg_module/gprf[650] ),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\reg_module/gprf[219] ),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\reg_module/gprf[719] ),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\reg_module/gprf[104] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\reg_module/gprf[588] ),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\reg_module/gprf[302] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\reg_module/gprf[307] ),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\reg_module/gprf[183] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\reg_module/gprf[825] ),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\reg_module/gprf[424] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\reg_module/gprf[168] ),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\reg_module/gprf[45] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\reg_module/gprf[853] ),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\reg_module/gprf[666] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\reg_module/gprf[87] ),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\reg_module/gprf[60] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\reg_module/gprf[772] ),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\reg_module/gprf[629] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\reg_module/gprf[357] ),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\reg_module/gprf[544] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\reg_module/gprf[764] ),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\reg_module/gprf[467] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\reg_module/gprf[586] ),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\reg_module/gprf[286] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\reg_module/gprf[654] ),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\reg_module/gprf[599] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\reg_module/gprf[175] ),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\reg_module/gprf[319] ),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\reg_module/gprf[497] ),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\reg_module/gprf[201] ),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(\reg_module/gprf[596] ),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\reg_module/gprf[630] ),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\reg_module/gprf[895] ),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\reg_module/gprf[778] ),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\reg_module/gprf[419] ),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\reg_module/gprf[598] ),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(\reg_module/gprf[835] ),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\reg_module/gprf[499] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\reg_module/gprf[606] ),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\reg_module/gprf[626] ),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\reg_module/gprf[734] ),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\reg_module/gprf[781] ),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\reg_module/gprf[651] ),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\reg_module/gprf[349] ),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\reg_module/gprf[744] ),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\reg_module/gprf[167] ),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\reg_module/gprf[81] ),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\reg_module/gprf[553] ),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(\reg_module/gprf[24] ),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\reg_module/gprf[683] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\reg_module/gprf[352] ),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\reg_module/gprf[750] ),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\reg_module/gprf[667] ),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\reg_module/gprf[660] ),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\reg_module/gprf[757] ),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\reg_module/gprf[163] ),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\reg_module/gprf[644] ),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\rReg_d[2] ),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\reg_module/gprf[6] ),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\reg_module/gprf[580] ),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\reg_module/gprf[462] ),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\reg_module/gprf[28] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\reg_module/gprf[856] ),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\reg_module/gprf[668] ),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\reg_module/gprf[450] ),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\reg_module/gprf[829] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\reg_module/gprf[627] ),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\reg_module/gprf[80] ),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\reg_module/gprf[838] ),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\reg_module/gprf[675] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\reg_module/gprf[46] ),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\reg_module/gprf[361] ),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\reg_module/gprf[210] ),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\reg_module/gprf[842] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\reg_module/gprf[290] ),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\reg_module/gprf[768] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\reg_module/gprf[313] ),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\reg_module/gprf[832] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\reg_module/gprf[542] ),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\reg_module/gprf[363] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\reg_module/gprf[989] ),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\reg_module/gprf[284] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\reg_module/gprf[263] ),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\reg_module/gprf[841] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\reg_module/gprf[585] ),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\reg_module/gprf[533] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\reg_module/gprf[199] ),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\reg_module/gprf[873] ),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\reg_module/gprf[440] ),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\reg_module/gprf[418] ),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\reg_module/gprf[983] ),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\reg_module/gprf[204] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\reg_module/gprf[736] ),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\reg_module/gprf[960] ),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\reg_module/gprf[754] ),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\reg_module/gprf[824] ),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\reg_module/gprf[94] ),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\reg_module/gprf[879] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\reg_module/gprf[839] ),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\reg_module/gprf[699] ),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\reg_module/gprf[949] ),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\reg_module/gprf[56] ),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\reg_module/gprf[664] ),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\reg_module/gprf[29] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\reg_module/gprf[779] ),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\reg_module/gprf[543] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\reg_module/gprf[717] ),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\reg_module/gprf[215] ),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\reg_module/gprf[170] ),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\reg_module/gprf[640] ),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\reg_module/gprf[15] ),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\reg_module/gprf[451] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\reg_module/gprf[659] ),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\reg_module/gprf[311] ),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\reg_module/gprf[852] ),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\reg_module/gprf[622] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\reg_module/gprf[367] ),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\reg_module/gprf[847] ),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\reg_module/gprf[427] ),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\reg_module/gprf[848] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\reg_module/gprf[965] ),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\reg_module/gprf[495] ),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\reg_module/gprf[25] ),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\reg_module/gprf[662] ),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\reg_module/gprf[477] ),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\reg_module/gprf[826] ),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\reg_module/gprf[476] ),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\reg_module/gprf[490] ),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\reg_module/gprf[534] ),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\reg_module/gprf[661] ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\reg_module/gprf[808] ),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\reg_module/gprf[14] ),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\reg_module/gprf[178] ),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\reg_module/gprf[807] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\reg_module/gprf[26] ),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\reg_module/gprf[82] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\reg_module/gprf[748] ),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\reg_module/gprf[713] ),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\reg_module/gprf[946] ),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\reg_module/gprf[669] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(\reg_module/gprf[874] ),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\reg_module/gprf[312] ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\reg_module/gprf[7] ),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\reg_module/gprf[828] ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\reg_module/gprf[863] ),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\reg_module/gprf[13] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\reg_module/gprf[123] ),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\reg_module/gprf[521] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\reg_module/gprf[336] ),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\reg_module/gprf[581] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\reg_module/gprf[383] ),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\reg_module/gprf[494] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(\reg_module/gprf[47] ),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\reg_module/gprf[928] ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\reg_module/gprf[956] ),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\reg_module/gprf[643] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(\reg_module/gprf[800] ),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\reg_module/gprf[257] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\reg_module/gprf[876] ),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\reg_module/gprf[570] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(\reg_module/gprf[160] ),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\reg_module/gprf[760] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\reg_module/gprf[646] ),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\reg_module/gprf[30] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\reg_module/gprf[265] ),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\reg_module/gprf[582] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\reg_module/gprf[8] ),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\reg_module/gprf[687] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\reg_module/gprf[600] ),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\reg_module/gprf[728] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\reg_module/gprf[968] ),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\reg_module/gprf[619] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\reg_module/gprf[729] ),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\reg_module/gprf[647] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\reg_module/gprf[604] ),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\reg_module/gprf[648] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\reg_module/gprf[354] ),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\reg_module/gprf[555] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\reg_module/gprf[844] ),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\reg_module/gprf[886] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\reg_module/gprf[657] ),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\reg_module/gprf[608] ),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\reg_module/gprf[301] ),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\reg_module/gprf[857] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\reg_module/gprf[858] ),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\reg_module/gprf[27] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\reg_module/gprf[860] ),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\reg_module/gprf[23] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\rReg_d[1] ),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\reg_module/gprf[684] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\reg_module/gprf[61] ),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\reg_module/gprf[653] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(\reg_module/gprf[539] ),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\reg_module/gprf[498] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(\reg_module/gprf[20] ),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\reg_module/gprf[567] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\reg_module/gprf[172] ),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\reg_module/gprf[890] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(\reg_module/gprf[205] ),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\reg_module/gprf[122] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(\reg_module/gprf[931] ),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\funct7[3] ),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(\reg_module/gprf[953] ),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\reg_module/gprf[528] ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(\reg_module/gprf[665] ),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\reg_module/gprf[963] ),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(\reg_module/gprf[371] ),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\reg_module/gprf[869] ),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\reg_module/gprf[877] ),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\reg_module/gprf[861] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(\reg_module/gprf[86] ),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\reg_module/gprf[862] ),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(\reg_module/gprf[843] ),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\reg_module/gprf[788] ),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(\reg_module/gprf[658] ),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\reg_module/gprf[655] ),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(\reg_module/gprf[948] ),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\reg_module/gprf[883] ),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\reg_module/gprf[671] ),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\reg_module/gprf[306] ),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\reg_module/gprf[855] ),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\reg_module/gprf[712] ),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\reg_module/gprf[31] ),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\reg_module/gprf[12] ),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\reg_module/gprf[277] ),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\reg_module/gprf[625] ),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\reg_module/gprf[195] ),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\reg_module/gprf[652] ),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(\reg_module/gprf[851] ),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\reg_module/gprf[538] ),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(\reg_module/gprf[283] ),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\reg_module/gprf[571] ),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\reg_module/gprf[700] ),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\reg_module/gprf[810] ),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\reg_module/gprf[740] ),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\reg_module/gprf[360] ),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(\reg_module/gprf[859] ),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\reg_module/gprf[880] ),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\reg_module/gprf[421] ),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\reg_module/gprf[780] ),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(\reg_module/gprf[610] ),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\reg_module/gprf[831] ),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(\reg_module/gprf[518] ),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\reg_module/gprf[849] ),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(\reg_module/gprf[5] ),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\reg_module/gprf[4] ),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(\reg_module/gprf[809] ),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\reg_module/gprf[806] ),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(\reg_module/gprf[971] ),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\reg_module/gprf[805] ),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(\reg_module/gprf[174] ),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\reg_module/gprf[318] ),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(\reg_module/gprf[709] ),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\reg_module/gprf[854] ),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(\reg_module/gprf[67] ),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\reg_module/gprf[718] ),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(\reg_module/gprf[731] ),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\reg_module/gprf[680] ),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(\reg_module/gprf[827] ),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\reg_module/gprf[685] ),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(\reg_module/gprf[986] ),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\reg_module/gprf[16] ),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(\reg_module/gprf[944] ),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\reg_module/gprf[866] ),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(\reg_module/gprf[836] ),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\reg_module/gprf[804] ),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(\reg_module/gprf[850] ),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\reg_module/gprf[602] ),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(\reg_module/gprf[52] ),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\reg_module/gprf[682] ),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(\reg_module/gprf[929] ),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\reg_module/gprf[771] ),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(\reg_module/gprf[276] ),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\reg_module/gprf[868] ),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\reg_module/gprf[601] ),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\reg_module/gprf[282] ),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(\reg_module/gprf[846] ),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\reg_module/gprf[845] ),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(\reg_module/gprf[590] ),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\reg_module/gprf[552] ),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(\reg_module/gprf[955] ),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\reg_module/gprf[9] ),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(\reg_module/gprf[18] ),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\reg_module/gprf[22] ),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\reg_module/gprf[950] ),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\reg_module/gprf[11] ),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\reg_module/gprf[882] ),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\reg_module/gprf[522] ),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(\reg_module/gprf[645] ),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\reg_module/gprf[840] ),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(\reg_module/gprf[202] ),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\reg_module/gprf[559] ),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(\reg_module/gprf[837] ),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\reg_module/gprf[801] ),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(\reg_module/gprf[867] ),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\reg_module/gprf[577] ),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(\reg_module/gprf[10] ),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\reg_module/gprf[44] ),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(\reg_module/gprf[519] ),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\reg_module/gprf[762] ),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(\reg_module/gprf[21] ),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\reg_module/gprf[885] ),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(\reg_module/gprf[656] ),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\reg_module/gprf[735] ),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(\reg_module/gprf[527] ),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\reg_module/gprf[116] ),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(\rReg_d[0] ),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\reg_module/gprf[566] ),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(\reg_module/gprf[173] ),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\reg_module/gprf[775] ),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(\brancher/rPc_current_reg2[22] ),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\reg_module/gprf[878] ),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(\reg_module/gprf[19] ),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\reg_module/gprf[732] ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(\reg_module/gprf[721] ),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\reg_module/gprf[564] ),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(\funct7[0] ),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\reg_module/gprf[540] ),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(\reg_module/gprf[97] ),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\reg_module/gprf[952] ),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(\reg_module/gprf[164] ),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\reg_module/gprf[535] ),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(\brancher/rPc_current_reg2[24] ),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\reg_module/gprf[756] ),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(\reg_module/gprf[811] ),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\reg_module/gprf[515] ),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(\reg_module/gprf[99] ),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\reg_module/gprf[603] ),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(\reg_module/gprf[941] ),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\reg_module/gprf[62] ),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(\reg_module/gprf[875] ),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\reg_module/gprf[517] ),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(\reg_module/gprf[32] ),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\reg_module/gprf[557] ),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(\reg_module/gprf[565] ),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\reg_module/gprf[2] ),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(\reg_module/gprf[536] ),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\reg_module/gprf[642] ),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(\reg_module/gprf[516] ),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\reg_module/gprf[541] ),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(\reg_module/gprf[786] ),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\reg_module/gprf[524] ),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(\reg_module/gprf[563] ),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\reg_module/gprf[884] ),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(\reg_module/gprf[1] ),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\reg_module/gprf[933] ),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(\reg_module/gprf[593] ),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\reg_module/gprf[959] ),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(\reg_module/gprf[3] ),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\reg_module/gprf[562] ),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(\reg_module/gprf[872] ),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\reg_module/gprf[51] ),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(\reg_module/gprf[0] ),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\reg_module/gprf[881] ),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(\reg_module/gprf[833] ),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\reg_module/gprf[54] ),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(\reg_module/gprf[560] ),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\reg_module/gprf[715] ),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(\reg_module/gprf[556] ),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\reg_module/gprf[938] ),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(\reg_module/gprf[932] ),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\reg_module/gprf[802] ),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(\reg_module/gprf[17] ),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\reg_module/gprf[943] ),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(\reg_module/gprf[65] ),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\reg_module/gprf[815] ),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(\reg_module/gprf[117] ),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\reg_module/gprf[942] ),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(\brancher/rPc_current_reg2[30] ),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\reg_module/gprf[681] ),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(\reg_module/gprf[958] ),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\reg_module/gprf[758] ),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(\brancher/rPc_current_reg2[18] ),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\reg_module/gprf[939] ),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(\reg_module/gprf[537] ),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\reg_module/gprf[370] ),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(\reg_module/gprf[547] ),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(op_consShf),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(\brancher/rPc_current_reg2[14] ),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\reg_module/gprf[819] ),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(\reg_module/gprf[165] ),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\reg_module/gprf[814] ),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(\reg_module/gprf[818] ),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\funct7[5] ),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(\reg_module/gprf[921] ),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\brancher/rPc_current_reg2[17] ),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(\reg_module/gprf[937] ),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\reg_module/gprf[957] ),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(\funct7[5] ),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\reg_module/gprf[605] ),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(\brancher/rPc_current_reg2[21] ),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\reg_module/gprf[616] ),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(\reg_module/gprf[834] ),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\brancher/rPc_current_reg2[26] ),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(\brancher/rPc_current_reg2[29] ),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\reg_module/gprf[917] ),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(\reg_module/gprf[525] ),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\reg_module/gprf[904] ),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(\reg_module/gprf[369] ),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\brancher/rPc_current_reg2[19] ),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(\reg_module/gprf[355] ),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(op_intRegReg),
    .X(net2066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(\funct7[4] ),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\reg_module/gprf[918] ),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(\funct7[1] ),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\reg_module/gprf[871] ),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(\reg_module/gprf[920] ),
    .X(net2071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(rJumping1),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(\funct7[4] ),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\reg_module/gprf[951] ),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(\brancher/rPc_current_reg2[31] ),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\reg_module/gprf[817] ),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(\reg_module/gprf[927] ),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\reg_module/gprf[520] ),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(\reg_module/gprf[954] ),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\reg_module/gprf[935] ),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(\brancher/rPc_current_reg2[20] ),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\reg_module/gprf[916] ),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(\brancher/rPc_current_reg2[13] ),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\reg_module/gprf[907] ),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(\reg_module/gprf[915] ),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\brancher/rPc_current_reg2[28] ),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(\brancher/rPc_current_reg2[16] ),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\reg_module/gprf[53] ),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(\reg_module/gprf[434] ),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\reg_module/gprf[923] ),
    .X(net2090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(\reg_module/gprf[822] ),
    .X(net2091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\brancher/rPc_current_reg2[23] ),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(\reg_module/gprf[913] ),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\reg_module/gprf[50] ),
    .X(net2094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(\brancher/rPc_current_reg2[7] ),
    .X(net2095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\reg_module/gprf[821] ),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(\reg_module/gprf[561] ),
    .X(net2097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\imm12_i_s[9] ),
    .X(net2098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(\brancher/rPc_current_reg2[12] ),
    .X(net2099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\reg_module/gprf[816] ),
    .X(net2100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(\reg_module/gprf[905] ),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\brancher/rPc_current_reg2[25] ),
    .X(net2102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(\reg_module/gprf[902] ),
    .X(net2103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\reg_module/gprf[887] ),
    .X(net2104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(\brancher/rPc_current_reg2[27] ),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\imm12_i_s[10] ),
    .X(net2106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(\reg_module/gprf[587] ),
    .X(net2107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\reg_module/gprf[940] ),
    .X(net2108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(\funct7[2] ),
    .X(net2109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\reg_module/gprf[526] ),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(\reg_module/gprf[906] ),
    .X(net2111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\brancher/rPc_current_reg2[8] ),
    .X(net2112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(\brancher/rPc_current_reg2[6] ),
    .X(net2113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\reg_module/gprf[267] ),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(\brancher/rPc_current_reg2[15] ),
    .X(net2115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\reg_module/gprf[903] ),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(\reg_module/gprf[870] ),
    .X(net2117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\brancher/rPc_current_reg2[5] ),
    .X(net2118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(\reg_module/gprf[529] ),
    .X(net2119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\brancher/rPc_current_reg2[11] ),
    .X(net2120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(\brancher/rPc_current_reg2[4] ),
    .X(net2121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\reg_module/gprf[924] ),
    .X(net2122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(\reg_module/gprf[936] ),
    .X(net2123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\reg_module/gprf[531] ),
    .X(net2124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(\reg_module/gprf[919] ),
    .X(net2125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\reg_module/gprf[926] ),
    .X(net2126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(\reg_module/gprf[514] ),
    .X(net2127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\reg_module/gprf[812] ),
    .X(net2128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(\reg_module/gprf[787] ),
    .X(net2129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\reg_module/gprf[55] ),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(\reg_module/gprf[368] ),
    .X(net2131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\brancher/rPc_current_reg2[2] ),
    .X(net2132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(\reg_module/gprf[523] ),
    .X(net2133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\reg_module/gprf[558] ),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(\imm12_i_s[5] ),
    .X(net2135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\reg_module/gprf[922] ),
    .X(net2136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(\reg_module/gprf[925] ),
    .X(net2137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\brancher/rPc_current_reg2[0] ),
    .X(net2138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(\reg_module/gprf[945] ),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\reg_module/gprf[98] ),
    .X(net2140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(\reg_module/gprf[813] ),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\imm12_i_s[7] ),
    .X(net2142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(\reg_module/gprf[532] ),
    .X(net2143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\reg_module/gprf[791] ),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(\reg_module/gprf[914] ),
    .X(net2145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\funct3[1] ),
    .X(net2146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(\brancher/rPc_current_reg2[1] ),
    .X(net2147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\reg_module/gprf[934] ),
    .X(net2148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(\brancher/rPc_current_reg2[3] ),
    .X(net2149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\reg_module/gprf[245] ),
    .X(net2150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(op_lui),
    .X(net2151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\reg_module/gprf[803] ),
    .X(net2152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(\reg_module/gprf[820] ),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\reg_module/gprf[254] ),
    .X(net2154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(\reg_s1[3] ),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\reg_module/gprf[398] ),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(\reg_module/gprf[231] ),
    .X(net2157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(\reg_module/gprf[275] ),
    .X(net2158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(\reg_module/gprf[399] ),
    .X(net2159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\reg_module/gprf[392] ),
    .X(net2160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(\reg_module/gprf[394] ),
    .X(net2161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\reg_module/gprf[243] ),
    .X(net2162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(\reg_module/gprf[912] ),
    .X(net2163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\reg_module/gprf[390] ),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(\imm12_i_s[11] ),
    .X(net2165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\reg_module/gprf[249] ),
    .X(net2166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(\reg_module/gprf[274] ),
    .X(net2167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\reg_module/gprf[393] ),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(\reg_module/gprf[259] ),
    .X(net2169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\reg_module/gprf[225] ),
    .X(net2170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(\reg_module/gprf[251] ),
    .X(net2171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\reg_module/gprf[253] ),
    .X(net2172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(\reg_module/gprf[133] ),
    .X(net2173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\reg_module/gprf[157] ),
    .X(net2174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(\reg_module/gprf[141] ),
    .X(net2175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\reg_module/gprf[391] ),
    .X(net2176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(\reg_module/gprf[405] ),
    .X(net2177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\funct7[6] ),
    .X(net2178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(\funct3[0] ),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\reg_module/gprf[412] ),
    .X(net2180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(op_memSt),
    .X(net2181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\reg_module/gprf[584] ),
    .X(net2182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(\reg_module/gprf[250] ),
    .X(net2183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(\reg_module/gprf[158] ),
    .X(net2184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(\reg_module/gprf[248] ),
    .X(net2185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\reg_module/gprf[404] ),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(\reg_module/gprf[823] ),
    .X(net2187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\reg_module/gprf[256] ),
    .X(net2188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(\reg_module/gprf[132] ),
    .X(net2189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\reg_module/gprf[400] ),
    .X(net2190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(\imm12_i_s[0] ),
    .X(net2191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\reg_module/gprf[224] ),
    .X(net2192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(\reg_module/gprf[641] ),
    .X(net2193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\reg_module/gprf[530] ),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(\reg_module/gprf[910] ),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\reg_module/gprf[247] ),
    .X(net2196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(\reg_module/gprf[407] ),
    .X(net2197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\reg_module/gprf[911] ),
    .X(net2198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(\reg_module/gprf[397] ),
    .X(net2199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\reg_module/gprf[395] ),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(\reg_module/gprf[246] ),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\reg_module/gprf[406] ),
    .X(net2202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(\reg_module/gprf[140] ),
    .X(net2203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\reg_module/gprf[159] ),
    .X(net2204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(\reg_module/gprf[138] ),
    .X(net2205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\reg_module/gprf[155] ),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(\reg_module/gprf[279] ),
    .X(net2207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\reg_module/gprf[909] ),
    .X(net2208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(\reg_module/gprf[150] ),
    .X(net2209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\reg_module/gprf[238] ),
    .X(net2210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(\imm12_i_s[4] ),
    .X(net2211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\reg_module/gprf[414] ),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(\reg_module/gprf[411] ),
    .X(net2213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\reg_module/gprf[135] ),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(\reg_module/gprf[240] ),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\reg_module/gprf[237] ),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(\reg_module/gprf[129] ),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(\reg_module/gprf[226] ),
    .X(net2218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(\reg_module/gprf[233] ),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\reg_module/gprf[232] ),
    .X(net2220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(\imm12_i_s[1] ),
    .X(net2221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\reg_module/gprf[269] ),
    .X(net2222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(\reg_module/gprf[153] ),
    .X(net2223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\reg_module/gprf[241] ),
    .X(net2224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(\reg_module/gprf[255] ),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\imm21_j[13] ),
    .X(net2226));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_0676_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\funct7[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\imm12_i_s[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\wAluA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\wAluA[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\wAluA[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\wAluOut[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\wAluOut[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\wRegWrData[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\wRegWrData[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\wRegWrData[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\wRegWrData[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(\wRegWrData[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(\wRegWrData[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(\wRegWrData[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\wRegWrData[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\wRegWrData[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\wRegWrData[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\wRs1Data[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\wRs1Data[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\wRs1Data[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\wRs1Data[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\wRs1Data[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\wRs1Data[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(\wRs1Data[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\wRs1Data[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\wRs1Data[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\wRs1Data[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\wRs1Data[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\wRs1Data[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\wRs1Data[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\wRs1Data[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\wRs1Data[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\wRs1Data[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(\wRs1Data[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(\wRs1Data[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(\wRs1Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(\wRs1Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(\wRs1Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(\wRs1Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(\wRs1Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(\wRs1Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(\wRs1Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(\wRs1Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(\wRs1Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(\wRs1Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(\wRs1Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(\wRs1Data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(\wRs2Data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(\wRs2Data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(\wRs2Data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(\wRs2Data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(\wRs2Data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(\wRs2Data[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(\wRs2Data[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(\wRs2Data[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(\wRs2Data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(\wRs2Data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(\wRs2Data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(\wRs2Data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(\wRs2Data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(\wRs2Data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(\wRs2Data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(\wRs2Data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(\wRs2Data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(\wRs2Data[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(\wRs2Data[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(\wRs2Data[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(\wRs2Data[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(\wRs2Data[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(\wRs2Data[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(\wRs2Data[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(\wRs2Data[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(\wRs2Data[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(\wRs2Data[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(\wRs2Data[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(\wRs2Data[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(\wRs2Data[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(\wRs2Data[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(\wRs2Data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(\wRs2Data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(\wRs2Data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(\wRs2Data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(\wRs2Data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(\wRs2Data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(\wRs2Data[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(\wRs2Data[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(\wRs2Data[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(\wRs2Data[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(\wRs2Data[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(\wRs2Data[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(\wRs2Data[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(\wRs2Data[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(\wRs2Data[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(\wRs2Data[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(\wRs2Data[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(\wRs2Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(\wRs2Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(\wRs2Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(\wRs2Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(\wRs2Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(\wRs2Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(\wRs2Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(\wRs2Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(\wRs2Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(\wRs2Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(\wRs2Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(\wRs2Data[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(\wRs2Data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(\wRs2Data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(\wRs2Data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(\wRs2Data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(\wRs2Data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(\wRs2Data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(\wRs2Data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(\wRs2Data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(\wRs2Data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(\wRs2Data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(\wRs2Data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(\wRs2Data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(\wRs2Data[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(\wRs2Data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(\alu/_0017_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(\brancher/rPc_current_reg1[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(\brancher/rPc_current_reg1[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(\brancher/rPc_current_reg1[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(\reg_module/_01147_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(\reg_module/_01147_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(\reg_module/_01147_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(\reg_module/_01147_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(\reg_module/_01147_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(\reg_module/_01147_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(\reg_module/_01147_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(\reg_module/_01147_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(\reg_module/_01147_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(\reg_module/_01147_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(\reg_module/_01147_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(\reg_module/_01147_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(\reg_module/_01147_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(\reg_module/_01147_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(\reg_module/_01151_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(\reg_module/_01151_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(\reg_module/_01151_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(\reg_module/_01155_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(\reg_module/_01155_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(\reg_module/_01155_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(\reg_module/_01155_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(\reg_module/_01155_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(\reg_module/_01156_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(\reg_module/_01183_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(\reg_module/_01183_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(\reg_module/_01183_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(\reg_module/_01254_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(\reg_module/_01254_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(\reg_module/_01254_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(\reg_module/_01254_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(\reg_module/_01254_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(\reg_module/_01283_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(\reg_module/_01283_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(\reg_module/_01283_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(\reg_module/_01283_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(\reg_module/_01301_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(\reg_module/_01301_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(\reg_module/_01301_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(\reg_module/_01301_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(\reg_module/_01301_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(\reg_module/_01315_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(\reg_module/_01348_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(\reg_module/_01371_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(\reg_module/_01371_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(\reg_module/_01371_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(\reg_module/_01371_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(\reg_module/_01382_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(\reg_module/_01382_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(\reg_module/_01382_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(\reg_module/_01382_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(\reg_module/_01408_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(\reg_module/_01408_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(\reg_module/_01408_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(\reg_module/_01412_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(\reg_module/_01412_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(\reg_module/_01412_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(\reg_module/_01412_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(\reg_module/_01412_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(\reg_module/_01412_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(\reg_module/_01455_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(\reg_module/_01455_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(\reg_module/_01455_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(\reg_module/_01542_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(\reg_module/_01542_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(\reg_module/_01542_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(\reg_module/_01619_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(\reg_module/_01619_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(\reg_module/_01619_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(\reg_module/_01699_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(\reg_module/_01699_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(\reg_module/_01699_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(\reg_module/_01699_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(\reg_module/_01699_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(\reg_module/_01699_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(\reg_module/_01771_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(\reg_module/_01771_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(\reg_module/_01771_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(\reg_module/_01858_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(\reg_module/_01858_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(\reg_module/_01868_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(\reg_module/_01868_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(\reg_module/_01868_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(\reg_module/_01932_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(\reg_module/_01932_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(\reg_module/_01974_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(\reg_module/_01974_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(\reg_module/_02022_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(\reg_module/_02022_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(\reg_module/_02022_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(\reg_module/_02075_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(\reg_module/_02075_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(\reg_module/_02111_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(\reg_module/_02111_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(\reg_module/_02170_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(\reg_module/_02194_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(\reg_module/_02194_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(\reg_module/_02198_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(\reg_module/_02284_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(\reg_module/_02491_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(\reg_module/_02491_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(\reg_module/_02492_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(\reg_module/_02492_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(\reg_module/_02498_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(\reg_module/_02498_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(\reg_module/_02498_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(\reg_module/_02503_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(\reg_module/_02503_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(\reg_module/_02503_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(\reg_module/_02503_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(\reg_module/_02513_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(\reg_module/_02516_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(\reg_module/_02522_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(\reg_module/_02522_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(\reg_module/_02522_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(\reg_module/_02522_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(\reg_module/_02523_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(\reg_module/_02523_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(\reg_module/_02530_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(\reg_module/_02535_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(\reg_module/_02538_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(\reg_module/_02538_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(\reg_module/_02538_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(\reg_module/_02545_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(\reg_module/_02545_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(\reg_module/_02545_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(\reg_module/_02545_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(\reg_module/_02545_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(\reg_module/_02545_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(\reg_module/_02545_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(\reg_module/_02553_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(\reg_module/_02553_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(\reg_module/_02562_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(\reg_module/_02562_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(\reg_module/_02562_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(\reg_module/_02562_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(\reg_module/_02565_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(\reg_module/_02565_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(\reg_module/_02584_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(\reg_module/_02584_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(\reg_module/_02584_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(\reg_module/_02587_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(\reg_module/_02587_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(\reg_module/_02587_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(\reg_module/_02595_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(\reg_module/_02595_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(\reg_module/_02595_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(\reg_module/_02604_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(\reg_module/_02614_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(\reg_module/_02614_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(\reg_module/_02736_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(\reg_module/_02736_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(\reg_module/_02736_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(\reg_module/_02897_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(\reg_module/_02897_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(\reg_module/_04154_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(\reg_module/_05034_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(\reg_module/_05034_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(\reg_module/_05034_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(\reg_module/_05034_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(\reg_module/_05034_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(\reg_module/_05034_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(\reg_module/_05034_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(\reg_module/_05034_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(\reg_module/_05034_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(\reg_module/_05048_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(\reg_module/_05048_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(\reg_module/_05048_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(\reg_module/_05086_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(\reg_module/_05086_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(\reg_module/_05086_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(\reg_module/_05091_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(\reg_module/_05091_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(\reg_module/_05094_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(\reg_module/_05094_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(\reg_module/_05100_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(\reg_module/_05100_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(\reg_module/_05100_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(\reg_module/_05109_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(\reg_module/_05204_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(\reg_module/_05204_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(\reg_module/_05282_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(\reg_module/_05282_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(\reg_module/_05282_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(\reg_module/_05282_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(\reg_module/_05287_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(\reg_module/_05287_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(\reg_module/_05287_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(\reg_module/_05287_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(\reg_module/_05290_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(\reg_module/_05290_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(\reg_module/_05290_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(\reg_module/_05290_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(\reg_module/_05477_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(\reg_module/_05538_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(\reg_module/_05538_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(\reg_module/_05538_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(\reg_module/_05964_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(\reg_module/_06905_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(\reg_module/_07632_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_328 (.DIODE(\reg_module/_07632_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_329 (.DIODE(\reg_module/_07632_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_330 (.DIODE(\reg_module/_07632_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_331 (.DIODE(\reg_module/_07632_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_332 (.DIODE(\reg_module/_07641_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_333 (.DIODE(\reg_module/_07641_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_334 (.DIODE(\reg_module/_07641_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_335 (.DIODE(\reg_module/_07641_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_336 (.DIODE(\reg_module/_07645_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_337 (.DIODE(\reg_module/_07648_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_338 (.DIODE(\reg_module/_07648_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_339 (.DIODE(\reg_module/_07655_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_340 (.DIODE(\reg_module/_07655_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_341 (.DIODE(\reg_module/_07655_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_342 (.DIODE(\reg_module/_07655_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_343 (.DIODE(\reg_module/_07655_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_344 (.DIODE(\reg_module/_07662_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_345 (.DIODE(\reg_module/_07662_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_346 (.DIODE(\reg_module/_07768_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_347 (.DIODE(\reg_module/_07768_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_348 (.DIODE(\reg_module/_07781_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_349 (.DIODE(\reg_module/_07781_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_350 (.DIODE(\reg_module/_07781_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_351 (.DIODE(\reg_module/_07781_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_352 (.DIODE(\reg_module/_07812_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_353 (.DIODE(\reg_module/_07812_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_354 (.DIODE(\reg_module/_07812_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_355 (.DIODE(\reg_module/_07812_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_356 (.DIODE(\reg_module/_07812_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_357 (.DIODE(\reg_module/_07818_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_358 (.DIODE(\reg_module/_07819_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_359 (.DIODE(\reg_module/_07819_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_360 (.DIODE(\reg_module/_07819_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_361 (.DIODE(\reg_module/_07819_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_362 (.DIODE(\reg_module/_07986_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_363 (.DIODE(\reg_module/_08017_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_364 (.DIODE(\reg_module/_08017_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_365 (.DIODE(\reg_module/_08017_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_366 (.DIODE(\reg_module/_08017_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_367 (.DIODE(\reg_module/_08020_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_368 (.DIODE(\reg_module/_08020_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_369 (.DIODE(\reg_module/_08020_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_370 (.DIODE(\reg_module/_08178_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_371 (.DIODE(\reg_module/_08178_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_372 (.DIODE(\reg_module/_08178_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_373 (.DIODE(\reg_module/_08178_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_374 (.DIODE(\reg_module/_08178_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_375 (.DIODE(\reg_module/_08184_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_376 (.DIODE(\reg_module/_08186_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_377 (.DIODE(\reg_module/_08186_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_378 (.DIODE(\reg_module/_08186_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_379 (.DIODE(\reg_module/_08274_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_380 (.DIODE(\reg_module/_08361_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_381 (.DIODE(\reg_module/_08361_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_382 (.DIODE(\reg_module/_08361_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_383 (.DIODE(\reg_module/_08361_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_384 (.DIODE(\reg_module/_08361_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_385 (.DIODE(\reg_module/_08361_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_386 (.DIODE(\reg_module/_08364_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_387 (.DIODE(\reg_module/_08364_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_388 (.DIODE(\reg_module/_08364_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_389 (.DIODE(\reg_module/_08372_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_390 (.DIODE(\reg_module/_08372_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_391 (.DIODE(\reg_module/_08372_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_392 (.DIODE(\reg_module/_08372_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_393 (.DIODE(\reg_module/_08418_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_394 (.DIODE(\reg_module/_08422_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_395 (.DIODE(\reg_module/_08523_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_396 (.DIODE(\reg_module/_08523_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_397 (.DIODE(\reg_module/_08523_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_398 (.DIODE(\reg_module/_08523_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_399 (.DIODE(\reg_module/_08523_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_400 (.DIODE(\reg_module/_08523_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_401 (.DIODE(\reg_module/_08526_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_402 (.DIODE(\reg_module/_08526_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_403 (.DIODE(\reg_module/_08544_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_404 (.DIODE(\reg_module/_08544_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_405 (.DIODE(\reg_module/_08649_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_406 (.DIODE(\reg_module/_08649_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_407 (.DIODE(\reg_module/_08649_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_408 (.DIODE(\reg_module/_08649_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_409 (.DIODE(\reg_module/_08649_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_410 (.DIODE(\reg_module/_08653_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_411 (.DIODE(\reg_module/_08653_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_412 (.DIODE(\reg_module/_08653_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_413 (.DIODE(\reg_module/_08663_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_414 (.DIODE(\reg_module/_08663_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_415 (.DIODE(\reg_module/_08663_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_416 (.DIODE(\reg_module/_08663_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_417 (.DIODE(\reg_module/_08663_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_418 (.DIODE(\reg_module/_08663_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_419 (.DIODE(\reg_module/_08663_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_420 (.DIODE(\reg_module/_08663_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_421 (.DIODE(\reg_module/_08663_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_422 (.DIODE(\reg_module/_08829_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_423 (.DIODE(\reg_module/_08829_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_424 (.DIODE(\reg_module/_08829_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_425 (.DIODE(\reg_module/_08873_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_426 (.DIODE(\reg_module/_08877_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_427 (.DIODE(\reg_module/_08877_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_428 (.DIODE(\reg_module/_08877_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_429 (.DIODE(\reg_module/_08949_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_430 (.DIODE(\reg_module/_08949_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_431 (.DIODE(\reg_module/_08953_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_432 (.DIODE(\reg_module/_08954_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_433 (.DIODE(\reg_module/_08954_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_434 (.DIODE(\reg_module/_08957_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_435 (.DIODE(\reg_module/_08957_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_436 (.DIODE(\reg_module/_08957_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_437 (.DIODE(\reg_module/_08994_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_438 (.DIODE(\reg_module/_08994_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_439 (.DIODE(\reg_module/_08994_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_440 (.DIODE(\reg_module/_08994_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_441 (.DIODE(\reg_module/_08994_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_442 (.DIODE(\reg_module/_09027_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_443 (.DIODE(\reg_module/_09027_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_444 (.DIODE(\reg_module/_09027_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_445 (.DIODE(\reg_module/_09027_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_446 (.DIODE(\reg_module/_09047_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_447 (.DIODE(\reg_module/_09047_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_448 (.DIODE(\reg_module/_09132_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_449 (.DIODE(\reg_module/_09132_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_450 (.DIODE(\reg_module/_09201_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_451 (.DIODE(\reg_module/_09201_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_452 (.DIODE(\reg_module/_09201_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_453 (.DIODE(\reg_module/_09201_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_454 (.DIODE(\reg_module/_09504_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_455 (.DIODE(\reg_module/_09618_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_456 (.DIODE(\reg_module/_09625_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_457 (.DIODE(\reg_module/_09625_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_458 (.DIODE(\reg_module/_09756_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_459 (.DIODE(\reg_module/_09756_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_460 (.DIODE(\reg_module/_09756_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_461 (.DIODE(\reg_module/_09756_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_462 (.DIODE(\reg_module/_09756_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_463 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_464 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_465 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_466 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_467 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_468 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_469 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_470 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_471 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_472 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_473 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_474 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_475 (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_476 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_477 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_478 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_479 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_480 (.DIODE(net353));
 sky130_fd_sc_hd__diode_2 ANTENNA_481 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_482 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_483 (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_484 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_485 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_486 (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_487 (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_488 (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_489 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_490 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_491 (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_492 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_493 (.DIODE(net387));
 sky130_fd_sc_hd__diode_2 ANTENNA_494 (.DIODE(net390));
 sky130_fd_sc_hd__diode_2 ANTENNA_495 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_496 (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_497 (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_498 (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_499 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_500 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_501 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_502 (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_503 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_504 (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_505 (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 ANTENNA_506 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_507 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_508 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA_509 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA_510 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA_511 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_512 (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_513 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_514 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA_515 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_516 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_517 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_518 (.DIODE(net809));
 sky130_fd_sc_hd__diode_2 ANTENNA_519 (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA_520 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_521 (.DIODE(net881));
 sky130_fd_sc_hd__diode_2 ANTENNA_522 (.DIODE(net970));
 sky130_fd_sc_hd__diode_2 ANTENNA_523 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_524 (.DIODE(net984));
 sky130_fd_sc_hd__diode_2 ANTENNA_525 (.DIODE(net990));
 sky130_fd_sc_hd__diode_2 ANTENNA_526 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_527 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_528 (.DIODE(net993));
 sky130_fd_sc_hd__diode_2 ANTENNA_529 (.DIODE(net1031));
 sky130_fd_sc_hd__diode_2 ANTENNA_530 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_531 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA_532 (.DIODE(net1067));
 sky130_fd_sc_hd__diode_2 ANTENNA_533 (.DIODE(\wAluOut[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_534 (.DIODE(\wAluOut[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_535 (.DIODE(\wAluOut[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_536 (.DIODE(\wAluOut[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_537 (.DIODE(\wRs1Data[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_538 (.DIODE(\wRs1Data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_539 (.DIODE(\wRs2Data[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_540 (.DIODE(\wRs2Data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_541 (.DIODE(\alu/_0203_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_542 (.DIODE(\dec/_112_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_543 (.DIODE(\reg_module/_01124_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_544 (.DIODE(\reg_module/_01156_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_545 (.DIODE(\reg_module/_01408_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_546 (.DIODE(\reg_module/_01455_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_547 (.DIODE(\reg_module/_01458_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_548 (.DIODE(\reg_module/_01458_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_549 (.DIODE(\reg_module/_01545_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_550 (.DIODE(\reg_module/_01545_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_551 (.DIODE(\reg_module/_01545_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_552 (.DIODE(\reg_module/_01702_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_553 (.DIODE(\reg_module/_01702_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_554 (.DIODE(\reg_module/_01702_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_555 (.DIODE(\reg_module/_01856_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_556 (.DIODE(\reg_module/_01856_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_557 (.DIODE(\reg_module/_01868_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_558 (.DIODE(\reg_module/_01932_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_559 (.DIODE(\reg_module/_02010_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_560 (.DIODE(\reg_module/_02010_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_561 (.DIODE(\reg_module/_02086_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_562 (.DIODE(\reg_module/_02192_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_563 (.DIODE(\reg_module/_02192_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_564 (.DIODE(\reg_module/_02210_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_565 (.DIODE(\reg_module/_02368_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_566 (.DIODE(\reg_module/_02368_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_567 (.DIODE(\reg_module/_02523_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_568 (.DIODE(\reg_module/_02523_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_569 (.DIODE(\reg_module/_02553_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_570 (.DIODE(\reg_module/_02604_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_571 (.DIODE(\reg_module/_02604_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_572 (.DIODE(\reg_module/_02604_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_573 (.DIODE(\reg_module/_02604_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_574 (.DIODE(\reg_module/_02604_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_575 (.DIODE(\reg_module/_02614_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_576 (.DIODE(\reg_module/_02614_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_577 (.DIODE(\reg_module/_05022_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_578 (.DIODE(\reg_module/_05094_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_579 (.DIODE(\reg_module/_05100_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_580 (.DIODE(\reg_module/_05100_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_581 (.DIODE(\reg_module/_05287_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_582 (.DIODE(\reg_module/_07525_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_583 (.DIODE(\reg_module/_07525_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_584 (.DIODE(\reg_module/_07573_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_585 (.DIODE(\reg_module/_07641_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_586 (.DIODE(\reg_module/_07641_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_587 (.DIODE(\reg_module/_07645_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_588 (.DIODE(\reg_module/_07648_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_589 (.DIODE(\reg_module/_07648_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_590 (.DIODE(\reg_module/_07768_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_591 (.DIODE(\reg_module/_08020_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_592 (.DIODE(\reg_module/_08023_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_593 (.DIODE(\reg_module/_08023_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_594 (.DIODE(\reg_module/_08364_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_595 (.DIODE(\reg_module/_08364_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_596 (.DIODE(\reg_module/_08367_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_597 (.DIODE(\reg_module/_08573_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_598 (.DIODE(\reg_module/_08837_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_599 (.DIODE(\reg_module/_08873_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_600 (.DIODE(\reg_module/_08873_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_601 (.DIODE(\reg_module/_08877_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_602 (.DIODE(\reg_module/_08877_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_603 (.DIODE(\reg_module/_08949_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_604 (.DIODE(\reg_module/_08949_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_605 (.DIODE(\reg_module/_08953_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_606 (.DIODE(\reg_module/_08953_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_607 (.DIODE(\reg_module/_08953_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_608 (.DIODE(\reg_module/_09078_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_609 (.DIODE(\reg_module/_09078_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_610 (.DIODE(\reg_module/_09078_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_611 (.DIODE(\reg_module/_09132_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_612 (.DIODE(\reg_module/_09703_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_613 (.DIODE(\reg_module/_09703_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_614 (.DIODE(\reg_module/_09741_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_615 (.DIODE(\reg_module/_09741_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_616 (.DIODE(\reg_module/_09741_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_617 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_618 (.DIODE(net356));
 sky130_fd_sc_hd__diode_2 ANTENNA_619 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_620 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_621 (.DIODE(net381));
 sky130_fd_sc_hd__diode_2 ANTENNA_622 (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_623 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_624 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_625 (.DIODE(net753));
 sky130_fd_sc_hd__diode_2 ANTENNA_626 (.DIODE(net1068));
 sky130_fd_sc_hd__diode_2 ANTENNA_627 (.DIODE(\reg_module/_02010_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_628 (.DIODE(\reg_module/_02897_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_629 (.DIODE(\reg_module/_02897_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_630 (.DIODE(\reg_module/_07648_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_631 (.DIODE(\reg_module/_07648_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_632 (.DIODE(\reg_module/_08028_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_633 (.DIODE(\reg_module/_08028_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_634 (.DIODE(\reg_module/_08837_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_635 (.DIODE(\reg_module/_09741_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_636 (.DIODE(net395));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1193 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_980 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_896 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_690 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_959 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1059 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_815 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_927 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1046 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_590 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1102 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1039 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1093 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_880 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1094 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1176 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_968 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_983 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1188 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1215 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_506 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1067 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1219 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1148 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1186 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1215 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1220 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_983 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1143 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_834 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1181 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_984 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1182 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1206 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1242 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1183 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1140 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1172 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1214 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1226 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1197 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1169 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1136 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1086 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1042 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1103 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1222 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1243 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1192 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1233 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_476 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1199 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_954 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1077 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1180 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1192 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1196 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1206 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_962 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1018 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1079 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1218 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1185 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1191 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_816 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_851 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1150 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1202 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_844 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1178 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1183 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_927 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1196 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_902 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1146 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1176 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1222 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1161 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1130 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1187 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_948 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1044 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1056 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1160 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1213 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1199 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1230 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1079 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1199 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_882 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1200 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_255 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1195 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1199 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_985 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1187 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1224 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_644 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_967 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1023 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1194 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1227 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1039 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_843 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1110 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1232 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1212 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1222 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1168 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1152 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1220 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1231 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1000 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1227 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_962 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1186 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1216 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_792 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1171 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_796 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_855 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_924 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1087 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1202 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_844 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1235 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1036 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1151 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1191 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1223 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1068 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1216 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1242 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1063 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1078 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1150 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1228 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_952 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1182 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1198 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1218 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1075 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1207 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1219 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1153 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1223 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_900 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1116 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1197 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1210 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1215 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1236 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1110 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1183 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_924 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1068 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1160 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1176 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1242 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_926 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1152 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1170 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1181 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1200 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1211 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1197 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1071 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1242 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_830 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1040 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1160 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1180 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1187 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1205 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1198 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_960 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1029 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1044 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1180 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1225 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1230 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1132 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1040 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1170 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1180 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1221 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1211 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_955 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1032 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1097 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1095 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1130 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1148 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1182 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1240 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1176 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_471 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1138 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1157 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1122 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1182 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1199 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1099 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1156 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1184 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1207 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_946 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1219 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1227 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1074 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1152 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_880 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_910 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_958 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1195 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1189 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1207 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_560 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1086 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1201 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1215 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1125 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1178 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1234 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1096 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1119 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1197 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1209 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1070 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1172 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1236 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1183 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1206 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_896 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1205 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1217 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1229 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1242 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1107 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1213 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1222 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1076 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1104 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1244 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1099 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1187 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1076 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1200 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1084 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1239 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1105 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1165 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1189 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1209 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1220 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1225 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1050 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1096 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_926 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_988 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1107 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1196 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1216 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1122 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1181 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1191 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1031 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1112 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1128 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1150 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1192 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1210 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1052 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1074 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_930 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1087 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1148 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1218 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_843 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_952 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1069 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_944 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1131 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1245 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1067 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1075 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1178 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_838 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_976 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1113 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_967 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_844 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_986 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1126 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1154 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1245 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1096 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1120 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1144 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1164 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1172 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1180 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1022 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1213 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1152 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_924 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1194 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1198 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1134 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1241 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_939 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_954 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1048 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1056 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1068 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1103 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1133 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1232 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1244 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1252 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_868 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_961 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1069 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1081 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1158 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1197 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1001 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1123 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1156 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1168 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1125 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1162 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1174 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1216 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_875 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1070 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1234 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1241 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1100 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1206 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1102 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1126 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1201 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1049 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1080 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1130 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1142 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1212 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1218 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1247 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1010 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1100 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1163 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1200 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1210 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1234 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1252 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1046 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1092 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1162 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1245 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_972 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1062 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1099 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1181 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1209 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1236 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_814 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_879 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_971 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1226 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1016 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1040 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1050 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1214 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_916 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1120 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1144 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1174 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1186 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1213 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1225 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_870 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1141 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1214 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1220 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1072 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1134 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1185 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1209 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_828 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1192 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1212 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_920 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1204 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_884 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1071 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1161 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1184 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1196 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_452 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_870 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_888 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1073 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1078 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1090 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1185 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1204 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1127 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1171 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1188 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1220 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1238 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_1250 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1039 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1138 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1170 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1196 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1170 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1187 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_946 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_982 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1083 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1207 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1219 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_784 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_903 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1013 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1122 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1142 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1183 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1036 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_886 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1064 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1072 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1097 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1106 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1124 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1216 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1014 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1175 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1204 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1208 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_791 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_947 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1048 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1104 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1113 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1160 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1181 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1234 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1032 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1086 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1098 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1110 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1148 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1160 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1186 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1195 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1207 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1058 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1066 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1155 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1183 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1190 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1209 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1236 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1252 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1068 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1080 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1092 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1143 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1188 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1200 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1212 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_955 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1157 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_990 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1072 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1152 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1184 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1215 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1221 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1017 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1136 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1180 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1187 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_883 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1054 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1064 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1114 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1154 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1190 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1203 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1208 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1223 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1235 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1247 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_980 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1038 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1098 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1143 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1165 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_875 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_944 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1123 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1135 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1191 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_850 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_928 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_985 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1038 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1070 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1094 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1158 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_860 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1014 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1168 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1241 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_874 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_931 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1015 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_1245 ();
endmodule
